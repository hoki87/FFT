��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�#&��#�<����軽���S8��A�>-?�������p��a�sx*|���~O�JC��'��l��Yὥhx�(���������	͠�i�+_C��w�pУFVf@v�r�Q)>�4A��B�x��lcU�w�ƈV1����C��l��͊~SJx���br�,��5�b�XS�	P��d�!��b�-���ز㖛+;L5�
�KP�Q�Fm{;�cNL����#U?ZK�Bb��:�}|���lEܧ�>W��[��=Y�����/i�wd�8M����	Y�h��HJ��-�Vi�iQr���'nCˎ���k�c�h�FG����-ψ'���L�ت[�.�`��@����R^`�O�׻[7¡�t��̿P�4f�b�����(��;�{0XͷH]���Q��5���w����Vfl�e{�X��M�x!�(���:�9y��9��$���)g�X�v/����'�w�I�TP�b����x5�3;:=���.�T�'���\�m2�^􄶟C�p�%A�5dP�cp��T��ۿ�$��`���X �XjΙW�	1�E��,旟4N�s�ō�F��-�q��؛˛v�J��͌3�6k�	�n+���z�
�~G����U�"�o�̠7Fw���D�YT�ޅsFR\.!�Z�m�־�{��+��/�z�Yw�)���aP�S�MnRV�,�UŬ���`8��4k�b�����ݏ�'�&�-�B�w��H$k{�R��e(��\��KK-fR����;�MZYi�����V��,��`C(���)P���9 ��_������ì���ӏ�1A��I�y��
������mi�o0�r���??��l����O<�'/����r����0	P���;X�_�~�f��J�<D H0#�<�ef�&�D}�~f�,�*��F���0|�^�"G����?h����84EG ����sL$��=��a�O�4��1��XO�^���W[�lx�g�R한��#�o^ӽO��D�S�(��N�E��: Rt\7X՗��ܖ�-?�{�f�IH���"���훧6,>e|���ĺ�O⭥�G$� R��<��۔k�]9�f�q	�^G��D&�%�{�V�����.�T���U��<nL����)օ0��VXY!jr�U���L�q\��j	��=��;9m[���Oo�4t���1?,)NZ�U�D ����M�I��ɲ�o���������~CU�$�����J@��_cT���v@�p�
A�O�K���ǁ�\�!"���,��Wp�ne���}e=���w.��a��xљ����Ә�ˮ�p]h#���y�9�Z.����}����s �{%ԑ�2�|M�VZ7t扞lx��·����e��by��6�U�|e�@�y�=9�XD�� T�������o�:ȥ�����\?`�J��u�Xp]�D컘C��g+/x_:�[�̿�_G�|?#L�X@�t��dV�S��n�?.n*������#O����Xm�y�{g�<M���==���#D�T߸ɚ�JE~�����k�4��g@�%&�k�ޢD=���F���Sv֏�������ۄ�v*ԗ��T'����s�A������#yT�7�x(<���Q�y��^`l!�O��:�da�~y*����"�[v�/��������`e��d����?�|�*1?9��Z�Lg0�e�t1�� `�M��FE{�7%OFTɮ�𬆸��6j���X�<�}�$I��1(��"_�
��tc(��O��'�~B�%ڪ����=�/���B
-��Fs��E���k��b�m�LJ���3]�L6).��� �z*��HJ5��E�nغb[|��7�Bi�\KP�'a&7)�\3��cC�4�l�>T�`WN	���Cn��"j��b�ف�X~C,�	��\�t��r�3�S�{��ؿ!���{7�Q�CS�'\�IZ�Λ�V[K�!�~ ��n�]�����⾷vFr�@�_�}|�$M����%�K���.`���L���N��YQ�����Re6ĭ$o�߁P��~���ؽ�?��\�T �-��Ӥ@}}vF�A+7�U�2�����}nT�N���L�"	"��G}�'��9z��TI�ܝ�Ⱦ4��0Q�z�E���^�!\n��0r8��j��H�>����l �3%]�x�,�����_~,X�>�?u��/4Gv��v�U���;*�/�a��:ԙWs�� �;��'�V�"A�߳ �m�Ko7/����Q���H�� y��o2=�Ѓ�0�� X��̤�J�=�BԎ�-�O=��&�n'��S�#�*e�S��%�+�)A~�uXX���~F_o�Eq�@>��e3�^�R��lPl8N�T�^���<ld�H�� ���z���;�.&���8�Xˬh�w�YS;�/	v)6+�ie;Ҹ����z՟Z�KW����Ie�l��}�%�7��q���7�@��Qfg�b�¾"�f	�\���E�?ɮ���7�{At&Ŵs���g�5�2cl|�saɳ�l�TEv��:� W��Ҫ^�o�<?�xE��ݢR���Ҭ�¡k�ƞ�(">�u:���Z��>*�.�B�7h�.է"�eE��<+����;��qQ�h������hw�������T?��Y�*���[vͽU���>+�#��y��m���L���tp6ɉ	[�6gNڌ71,F�'��F^R�����_�ޗBs��F*c�5�����1�h�!�Y���'aÉ�}��D&_��7e|����� }({�Y��YҘ��/��(�n|fI%�k���sjnv��s������q�a��HB�p��uy׍F|i���C���5�谆�`�̑/;��
�7ؚ�tT�+�iⅤ�:p�>��[��Ky�49�<T^_.����՟ǔ;����ި��ܕz��E�*��y�y�����x�Y�Sw�s ��a\�0��KoLoM:���=�����D��P�4��yf8BAeZ��� ��Ձ:�{#�&��e��vTr^~�t�xl�TL��+�����XJ��Ӿ�i�B�ܕ#�F��|�a��r��WL��!�z^�7>��6c��M�|�uff+�2��Yi#�U�-�dF�]������u�_K
��%NS��������	J+ⲧ�EL�wdG�'g(M?�M�����A��t�A� Jc�x�]X�-M����'o����r>;������P �h}��&�	\b�ԯ��]ON�+��)�r� ��u,�����ᴵ�S�y8��{ .��Fh�h�*8���|I=�e_�� [�(�%��G[{e2~��t�B��ߌ����dVY�������N�{�i\�+B��p�^"J����8����M�W#���f:!��}ǧ?x��i&dظ	�u��c�)C�g8kL��x����]`]*�c�Y\ج�XR�$�cW� &�)f��f���Zˢ�;	R3)]q�+��������FTA����[�ru�6&�6O
��|y�^7��-�3Լ��熗�9,6����M�ӽvF022��L��R�H�p�=������r�d��i�`��xIbX���U%���뽲��Ӵ�U�-��z��0w$�;9Պ��x�;�3���ar�k��z�7�)�=��e������:��d�!VBxU�eT���UPj�J�&��g*p}�O#�ڏw�U�F_H��"�LlVD�,s�[�]�bĒ��a+�!�L��"n���{������i5�-�c����|���i���f}��0�B�C�)��97�Z�X[W'���>��(�[���1�+@tw�P�? 1P(`�
�Ⱦae��Bah"}U��Q��]8	�凄M���Se��6F�M=`���vS�|���Z; �S6Y��b��={%Ԣ��lچ�t=Sߌ|���=,����t����)�c�?����\C��������	��t�sq�=G�}v�c�	�ͨ�\�&�i�K~8��ǟ��3/�,J���@��>Q�T�����x�8@"-ք2��Su��z��N͟@cе�Ћ�0 =G%��ڱ!7�)��⧛�z'�����f)�g�p���ʗ��k��@��:��;�ƅZ�\�ʬE*T��GɆ�Ka�Y�T��F.�;��ԝ|�c�,�~~��Iw`�H��� !�J4)�S?�����6�એ���v+&�>����n���i����+��!��VbX�>nI��Q$E�`CT	��C�����,�X6���2�lrl�D��B^��2���C#QSڦ���V��`�a���M���Pư)b�ԏ# �n�K�$C�Vn����>��X_K����t)y}aI�1V�B�.H��9r�ج��`��nZ�`�KFi����U4�%9�I����G�׈��H����r����+$;�Z�p��V�~����#�ݖ�m�e����U���"gg��(ܒҼ�������"1C[њ�[��WƷ�} �A���,�։@��A��<1�e���BЛc���.#r�]ٓp��P07Bh\�N���&�fL�T+;M�i2!���$	Mb��2��y.�33zd�p���=!Ϲm�M7?��I-Ƚ����n��VPM|H��+�<"l1�I�ł�w0�q�ӿ��Oe�tֺ8]����:e�m�۰�o���4sƀ�]�K,~�|�l�5>���>�JJ*K������{9��<��OΤ��B�����8|�,x��>h�j�U������ʛ��I���pugHX��v5��a�$�8߅.�l����v�o�M&H�x;�olf>_���q<�2��!��[��B�Qa`��9�zl��2�0�����`6g���D
'�x��nš=�IQ���� �W�H�t���'�:��>gup߶��s�S���u09�ޑ���tW��{D@�h����l���������udp�EBm�p����OK�[ph�=����WU�RǗ�F�?ؤUH4�h	�L��_��ʫ���6�Ī.�S�~F�'�Zn-i��r0 ��Vӆ��׬0X7y̰�)��A�r���|P��LĢ""�si&�J��d����Ɉ�Z]Z�UA�%5�σd�αj%-�~��x�?�Ӕ?}9�R�ڧ1j�2!}?&��
�b��L�1ڜ��`�Mn�Y�SO=�������f�[I��HW;���F+��f����c銖����RJJ^X�0Y;{�i&��G�To��~�����NF;6j�����x ���TGwo�j�(�2È���!�7��I+�~��� ֳG~�
��t��\����ހ޶8&ɜJI�C�%�=if��B�<;&.�/��|?���A��*5Q�� 7�n�z�5�br�s6#�&�Z��|09��;C���'�Y��f"B��;I)[�����h�^>��(�f�;�kzuR��Q	8����@
5������_�β���J��'HlT.(�����_>��������I�j��)_��1��=�i�V��� �bJ���
��Q�5���.h:>�S���-���O�$m3q��]��3(Qk�
G��2���4�u��$`�ĈD+��@OP���S�I�s�Pr����W�_�@��O��bW\d@�v}*�k�'��2�]����4�W
_��V(uVƘ<�4R4~J�L�8���NE�R��+NUӥ�u��'���[hx���|�0�TΗ�K�]��aq��<����+����ÿ�}ym:f��09�����'#��f���o�rN�ec:l����*;�,���l�g����U}��7\7�yh�ࣽh_�V'�|�I'�xjk�4�����-w�w�!$���� ���.h7��D5�b?��@��x�g*���k�3��\�a��묹C@�M)'&�8��\�^D�=�o��ќH�b/
U�
�/U�Q׃*�֊�>�]�E�Ho"{�T���A��0#d�1D��V`=Z~\�^�>'��i�L�2�;��ar�S�{�r�n�RNǞ��>+���F�m�cA��zy���zLqJ� *�]b��;J�p���_����茊�,�oNU�L�($���m"���g��H-~o������Yw����� �-�>�iP:��Z�DѸ-S{Q��$�=ɦ�4~�Β�T���7�.x8�sY������� 㥄>(.u��<�{�wI��4����݇wP����f]�Z���]4�_���)�x-�
@ #��l5{��`�^8�z�`q�3(#ù���A���e�ǛZ(<6����k���X`�Q0"��@$�6|;Wh���|G";z�� tc����ʗ��7i�bo٨n�����do�� T�a�����ͪ�9�I������sYox�-յ�c�试�M�/%�"��y�c��'�j��E&�� -*�ya��"n��C�U?N#���z�
�g���D/�]BqH<P��Q��q�E����ΥkP�.uL�%p�S�T^���Թ!��JO�� o����`+�p�M�׷?���� �I�Ȧ����:���ն|�5��+֕��}-�M$«1	�~��3ŝr����$�f;�T񩷄ht%�1�e�[��3�o,X'��/= ���	bs�m%�4tO�'c�*�.�rԧ\���/��=,�d�C!�1Ӧν��Q�߫<͆\����h��K�����]ӥ+4��:��36:�!��j�cMni]�Zf���@c°z�_$�����w��`v�@iĒ8��懣/� ���'�|�믉.�Y��
j�$e��Q��S��I4.��2�1}�Gп��-�+k0�xd$��4)��֧�2����@~@�o����%k'�-�1��r��C��\����X�UOA�|��~�m6��NG��$�G�p�����e��	6����K�L��uT��h�Q#�M�g}>�Ǫݩ?�<����d�����{�C�v𯄇���UKU�Z�H�n�l��w=_,�L~^ܵ�}��c]�j潕%�)����?@�bN����U�(���$�'���-�LG�L}�p�Aa��AQ�y���f�-�ަq�`����P4� V��WFBL.�ez_���dB�\[�+�>!2$�L*��4�Z5)�ԗ����|\Iݍ�L�X�G/���\������8���)����P�O��p��~�d�($R���9J�gT�}���p6.�"��*�y�/�m�rō����Gt�0~y��-@)�ju>����B+�!j��'�W�\Q�Y=���Y�C�ٕ��I��86k	�4��]�K0
Y�JGd�+棆�?_�mB��i�-y��Y,Rƙ��QQ>����P,�4CHs2��O4���	�zn���0	;Bʵ�c��R�b�ʶ����q���;�k�� L%vR�:f�8����s8*����7j�e vz=F�2����w���VG�����
�PM�̕��bl}���1="a֝ǃh6kv�>�Xcތ�	�pZe�h��G0����y��b@h��1�2�/����������%�k��˜�H�a|M*�1��Sd���\m���)c;,��-`
�Kak^=�J��n����H��}x����fL�P������.�c���@P��;Q@b�i3	��L�4�V�~����\ܔ�m��9���m֘4�#�iv�?U�#D4P��)�}eg�s[�p�'�U�Z͙!�5/�N���.kD�i�A�vF��%�ՓSrt\U��4��/�îq�Y��_n��F�C����y����f���]���� EM�x�_������o����.q�5>l�<�݊d������ŉ�����θꇋ���.�23ǥ�b�V�e@��s�X��e���Y�����J�E6}��V��'4�D�U���H�?�3<��{�Aݭ�2�8�yp
��"��H��'�c�wަ��/�Sl~Zp����SU�e-�0�k�X'���sD �o��n_������O�C�����ߔFD�� X���*���{�>l�U���ͬ�]C�T{��A둬���� 0/�ޛz�=�����6g��Bp+��j�$>bK{꺉\cw�?��K�cz�4���P�n([��[�Q�@�p�N�28��ǂ0f�	��`\�G�M�����]�E�/���A@Eq縦MOhI5�*7��_P ��ꗫ�,�dv�B����F�`q�,�/�|�c.�RA�����ˑ���TL��<�h�������	�f�驺?b����Ү7�;�wD]K�ۃ����I���{t���6w��&[�gV��9�:�I�
��8�d����|�{��q7�/+�灗[&��p�3��\4�T�<��t2ˑ%���N�o~���黁��m���t���M`Lk�h�\ż��X��e��d"8� ��ȟ�*����o.�,���p=;�=��SU
��`�h�	�UO���_�;s���`�=����$��H�ѵ_T�#�#���Jz��kX��̢�N��+��?�w;����Zf#�9�R�]�#Q��ŒP8��M����%����"X��&G��B�+�k~����n�����ӊ���ֻ��I��� �Z�˦xAJ�p���%�!@=��V7�� V���/{���Β跑�T��_�_f'���֣ѱ�ZBi�s�U[dS+�Dꬺ�P�|�*����Y�7���f�ߩ��?_�X�u�/0k����?��AJc�H��ut���hqc7/�$Գ~��ȖN����^
>��ߪW�:*yI��vRU~k�$jkK:��\���XQ��vX*6���_��m��oW��cw��"�@�"��G���x�w�|#���Bғa,�� �RF����C��[��&��t~&���,�"�PF>ZlD���O4���n��I���Fp���u���>m@p"Ӱ*VK�>6����Q��"�L=*�C���2)1��k�`�l�z�󩌈�aH���?hF�y�F�q�sK�J��>� �dV�J�!���j�Ѽyj�b�Fwk�����Z��v,��g�R'��U��+�h\��g�J��'�������:
�4<������e摬���uX�3�[�~ z9&�
.�ךj��O��mmG���.�bL�ѤS�'�¥C �瞳��Q�r�ʖ��ǧѾ��;&��~��N�!�K�kW�p����s�z/oW��~>�+c�`��:ڒ7T)��/Z_ +D��]~c-��߀63;�"s�S��ΝԆ
�{]8a���w��Ч�؀��3��F��)���ֻ��v͚a]�r ��#~��{Q�R��{[q55L���(���H���V������ɿ	��ٻ�ocΓ�v�F3��Q��ɣ�|�X�!Ub�1�����QU����ZW|<�r�Ȳ���C����	�:��#�c�)#�y��R2�rKqg��!T���wK���b�O6!1Ʒ�۪���o=LL��O�L���N�Z�\@|n�U5#t�ޠ�E��,ʹA�c��$�{��乒'`6?���S]�����ǧ�-��?f�E�� ޏ�&��f<��!�J����gOSMW��{����拫4$fC�ke�ӫ�w�ZQT�+6�tU.JB
L0t�2�	gO;B��_��i`]pO�Njj�޳O $a�XD�ħ�H|������&� �EU�KY��� f��
�"�V�oW�;`C�W9��O�A��e��V0r���\6M�&R�$|�{��@�� ���n�P�ۚ�-+�h��Z�cX{j�W�	���&����>�<��k��L-����ڧ��#i4���g�oEIO(� �q]�G����徭�qey����7%5�W��T�:Hz���<���pI�񣯈OD�Q���G��0�� ����f��v����d�b9���/n��'� �L3��a)�2�������x=��Dg#��%6���d^��,�D����w⫎�A�6�R�1��mj��'i����,���|~��[?�qd���%�У���zI�b]l6)8������UY��=-NbGޓ]c�w�E�-�[�^ss-���պ�����(P�<�5�^���/D��}�W]��'�8@�?�]�FP���2��>��n)S�fa�����=T�
�8�`��t���ղK=��gJ>Z�GA����)�AI�{�O����3q��X������tm�Q�ۮT�p�bm�$W-O�k�%�&(K]���Cp�U�w<����	�3����Ķ$�v֢���qE�3.�g׹ʹRXr�� �	�4c� �����o��\�GA;~?�2���IG��N��4�)�N&v߻�|#��9r~��U��J|D�������k-1c��G��彭}�����+�;v�v��joQ2�����n`���&jM����hH{�����^A��h�u�M똅a�j��8	��!�ħ��8�ԺH�q�7�Ue�f������#�*���{?L���A& �٘Ώ�]�U�<:�b��=�h�@�եM8��G�"�ߗn$����_)T�����6#���iG36��Rԣ8=�����N!M�UN�u��O��.wX�_�lyB�h��C����^!�-L	sge$�d�꒡)T�:q�}U��0,���k���z �F8Qn)����{��~xh�
f*v"6v�y�� e���}-���"m��ȏ��U�9YF����O���ƈ$�/чB�ʴ�i6��<�K��f��݉�._���?Z�9�SI-U*?<p�8��d��8=,"L���f��r)��.w��R]Z|�F�<�x�&����k�3�6�·/���-�P+$+����V���t@�n���v] ��,h�BA��C��fʋ�g���U�#�2�6�d��K	��W�W��L�*��T!a�T��c�݃}(���!��CpVQ����^���n���˞�8;���6o�f݃������=��T��i�zY�5�scB�Zm��m�B�jj�0s��-��� �4��U+��^c�������$|c���$�/=~s�.���������`M�[�u�20c�Pvaj7�E�wr4 	ɯ���U����t3 [�$/���J��Mk{��s�<��0���*
�AT�C��\�������Ԟ?A�`���X�\�u�Tia-�Hu����Ɍ�7����GT���4�?d7I(�}�s}��
W�duo2��h�N��.[r���Q��%�{I���v�Oܭ&��Ρ���:��-��E6ߘ�/u�� �������k�ˠPڨ&Y��-W$����"4�Oh�V��t%����(�� t�WI�h��fi�����s8��-�ffr�oT�]��/fd��G#�;�Ќh_�����k�P�=q�2�*��#c9�]_|`�q�;�a�/�"��.���,*�����i��2�P��=��ک�Auk ��)��Ą��Ne�61(�L7��׽i�
�kd�xv�ـj[��t���8}�]�7~�ŷ9��;�"fjû>	�s�b/�R���0Q���W�Jg�%D��9$�r&�&�V�%���<������(r��"�+7�uj�[X������o+�>��uG%0��ya�"_q
��˖%�,#Ɂ?��x]�7*��̽�v�ѵZǵ�g�׾i��u.t2�c(��5�2�N�,E����Eٞ]�����r���ހ��*J|z��Fn���Ѽ�r��Ȟ,�wo���U��{��8_s�b!���oE�����	��1f��`i*���ZV1��E�P�v��z�<���Y�pulF�r��+�P��>B�'|E��]Wց:���q$n�v����?����-�V3z��`�GO�үX��v=���H�%���IEV����~y+�E:�c�ϥhgř/��Z���e����u�����,�B�NXq��ܰ��׸��J]u�ӷ���s��j���ٲM	f������qfGE}����&�~�	�Kj��m+�����.�K�����{��.1��"���6�IЃ��t3�w�G?�����
B�荘ܕр�9�L7�����Zp�e�	z/��U�BT"��}6�G����+�z�v		��kI9~T�P��O�^S�i��	��9���<K���!�>kT�Mr��I���X��h|)�ŝ�դI�u�",4uu��	���I⦥_}| <7ٷ�o�Ԁ��� !�6~����\�(_\�����i\jf]�韨���)Ѐ�F đ���L�3[�/����
��,8�͋��{_��DOF\�d�Hzl��C /�M=�V�t.'-�&�X��BA{_^qȞصe��-�f�S�>�w������D0O�*�S�=��	�܌W�3|J���>KG�p(�~VJ�,�&�f��h�O�Q�;�ԵNX��5��`h��2?�����7�jkG�JI�;����S�~�@��N+_��_{C�w>���3���HG���:>&��4��4D襁HW��G2>��ݹ�Lc{�����g���\?�1�1�<㴜vs�9������T
d��6��� �P�u���i5g���Kv�`G�	d��d~*J�w� ��=ӗ�tg��l����<!-�	�,y~Ն^�w+��E�Rzj޸�u���b���f�th7�s��Q�2�˱��a~�n����?�
1ܺ���k"Nbg\�8�=�/�k2��K��<AB�s@� 'h�U(Ȓ�X����2���re����	� ���I������c���F�Cq���Р���m s�~�Z8���*MB�G��\�?�q�vf��jB�3=^n\Q�&aK>X�1�a�����,����Y�����N�SV�w�*<�����}�6�ȵ����PF���2�&�Q ���_/����H���7� hu�}�b�F�.O9J�ކq:Y�X��-TV틹s0oGM�V����bO��EK�7� %;v��g�G�ga�dlw.���p��إ�SfS$^��޸�څ���nq����9$���i��i��+�y�cz���#� ΍���{�F����Iq5�h4|�V��vMo��/�`"�
�_�1s��;уv����|���u:Q�+��Gc3�����x�ă;M&��|�M���M�n@�)9�{����Y8|�"�'U�����\$����zq$ݭ=rcS�D'��-⠄0���;s
1����ɂe�#�EQ܆��uK
�<�Л���iـ���Z�������K���Z"��S�����	��dCM_�d���F9%��6��s�X�a��e�8t%D���sA��ɗ
B�w�=�F��F�x�xS���3���c�f|�s$�'�}��!�o�	Q�����t�L(��zжF�*:�����%Lh1�.c���2]�2���Y4B=�M��Ŋp�n�U�g:hP��0�"�\t�m�i\ff��0����d����6'm~�0k�!
Z���X��*3s����*x��_��:�N�\�-��*0ne����2�3�ؑ.?������W�U�n�ͧ8��m�|oU}(��b��BH��>�|�����sA9�f��Dʒ��td��<��#�L��!�u�`_b_�4��Ok�b���({=A�IݺOBͪt�ckOsazH[sNI�JJ��:���� ��C�ڨ�$��?�DvR�����7��T�P�ؘ�K4���WI�k���؜����ll1�.I�A�����\�^`�8�8��did	�=�q�{0ÁѥQ�W&{f��|2FZc4><�Sg��������:���&7���;QS�5:�76R��ͱ#�N�����
�ƻ�$|چ�t��ݵ�?��4�69l	�ch����S�#
oj����%(|F���&6��e���L�v*���kO���W��S3[-�7�}�cl�7���Zak\$Xe�x��a��J���R�t�J�w�]�^9�Ӎ�17��,%S�\�m��tӇ�2L�c&%8�*C�S˄Q��74YY�Hhd�'Ӆ�	��6D�k��Z�z�@���wr�2��f�ь��,w�!_z�ܻ
y��][��?)p�Ag�0�l��d۹ÿC���'0�p��H��B���'t		��"�5�YD����M'9�6q��M��`V��Eke��q�NtΒ�Y��'zA�o�}U����2�B��l�<<!p\d�Rh
��Z��:!2﯋?��&��"A��G�6�>h�?~�e���Wd�N��Azp�O|9ϋ�I-kp̣G7�>��lI]2�Po��d�) r�Qʌh�*�tq�[��%0�	�a�I�0�^��>@,���Z�0˼N�U�IӒ���v�v�I�zւ��㶕��G�e�>8,�`�h~��������^�\P+E�=��w����;|$î� y���N� ���G�2��_�M�򽣛gL���'X����������N�k��ۓ�w�&0�����
�eXd`EZXG��QlJ�іy���&�r�4���D���I��,%�5����!�O���SGmY5�1͏��wy�����5����t��}�n�T��(oq��׈,(Pe���c�?~��ƶ��'���i�&]m�/(�k���k$��wP*%%B�[Đ�b5�]��h��0�{�
��.%߼�d�i�$�P��RĿ�W��Z��J�B�L�n�x�y�������13R{nH���]�`����[�.p�!�e��"��7�x�z-�E�	' ?m�N�������j�oo<�O] ��vb�d�/�EU��?*z4��p�A�$(���ki��^gH@'a
Es�?{ gA��'�Ib��j2Hr~}�y� �r������۾K�Yׂ�X[U.���U�̘�<���ӫv87E9���h�7LYW��W��~�]�r��kyލ�!�/�V]��g�⌎�*ڑ�MM�Ea�d��H��U먙я�KYu5q� 	��W������(	9����=�\��9�!N���[�C	B����A�)V~W�)	oH�� V���b��,J�y7�"����Q���俬ܯ�_cRƊ<����$7�wu�E�H�ق�R 5ja�=b�,�	���@9_&gV�8����ڴUAM�-k�J%t|ӣ�U6bPo~�s�k�W��aNh�=�AQo��0�@�៰J�4��g��l���ļWp�+�J��1�n�,��ʷ���kܾCT\�I���4h�$}��&e�+1�Җ_���̏�K����/&2k��ŃQ>,�s��5�qj���.d~������ܫ�.���h��ʵz�%�7���כ�piռʅv֧Q̖~����8:<w�d5�dѵ��� J�x�8�~�N7I�D��J�"�3�,�\��F*�i�����k�O�$-����j9��tg��0�qd0�i}��������h��n��Ģ��Xz<y����~k�/��<&u7!��ʧ��.���x��nr��������Hd�WC�@/p��V�c�d��C��E�����l<���"L�zm9b�¤>���Џ����d|�_��ͤT���������,������4)ƅ�B��E�� ��݌S,�H!.�����R/���3|�s�VE� $�i�:�L�Ώ��V����y�����V�
���k�-�vXɅ)����yu�B5�<9����(��KG^�����t@]���u <�����[-��X IO�+^��H��*"��og�/��*�4�[]��5�;��F����:�|��3�'iEp����ޭ����r:Z�o�c�\�z�+rA*$��(�{�ۅ���C�ML2���:"b�W��z&���[)�
 �p<>��zA��7�fЏ�T*��Ɯ)J�pV���[_��P���ձ�	s;�~7���-9)����/koS�1�&(Ä8��!�[C���<�w���p���:~���8����r��tN,�Ʈ��^�$n&zm��!l�DXM!e�F�Yvy�F�o˙�gO��].8A�W�E�/Ļ�ʷ���N'����`$�%[-E?�������
5�E!�#��ew�(�D�o���Q��r?&��9�I� $��|�o�5C�J�og�Ez��g#�-v��1��oj�w7�:���5��b�f�9ZH��[t�RX�Z�hk3�s�n;����c4۽�}�;��_�(D\�S��
�Ix��G'�}��e�~vf(�Le�s���=�8�ٶ��6- uY��b>�����C�tg�;S��0'�A���
�S�
�/�� <��/_�LԪ"�6�&h�o�_ِ��'��h��G�p�hP�*U�*j�n�l���!�#W��>��VP�H?���ߢ_�0A)>g��6QTi�8���ɵ���U1���*�w����y1F�������]�a�^29|�r$P��F6��}@�J�1����p��c= Ҋ����[ؐ��t�?X��B�����G	��)b��ډ �e��J3-/!�_2���Z«D���B0L�ǝ��iH���>��1]Qf��7�m�����~�cU��Q�:Oȯ)$�� -�)]*��7��Xel�'<<�MO*��P:j�!���b!a2�V#(M0����=a����1�%�ɬ�(Ĥ@��]��3�sg� �%�sU�CWI�k[�'�#	�ۚ�`�$.̘	&肪T��,>t�Eg�Θf6�
����(��A�Ș�łs7)q�,�80��&;-���*e�fN��b����Q�j ����S4m���J�$-��u�_�a0��ՒY�E��\#6UھQ��$N��d����x�-�	��}�����NnX���r���e�)��
�b�Ф��h ���0sלl��ȔҬT�/��u�W�u�N���������?m/�;�]���Yyo$�=����LX���-U����g��pI�Ox�I8PXKCm�d��0���Ί�^�W�k�9c�,�^�\���_V��FO%-��>.���?8�!<;��$���˂��g<{;��띋��J)@�Ŋ���}a3�7q3a$�����8r�{1��_PV�Q@�;:��L�M�k�#��BWڥ�L�iآ��{���4N�$�����
ti%�n�)q��:"�]���02�h�3�o٣PNo�K'��o��;�ο���[rEv��c�J��{k��%T����/ՕQ~�^a^�9�����C�U�⥓�	��B;�4���7Kh�F�	�Y�h��Ǉa��P=�]3d5�r/epZ*~���DF�y���k�k<�=���V��%�:���I����R@2���=M��n����a]4S����Ͳ�ٯ���s��-`�]*��"�dz�/����F���`�ymm�|�������#�kl���B��S�_g�� k���ܕ���|�'��]�t��7�0��Ⱥ�J,�������F����@�; ��='_]^n-c��h�Q/���@���k�&�Hw�����	�/3�?V~�(��Q��7Q���j$�+:�7��H{������`yB���oXE<l6�ȃ�p`���Фf�����9'z�J�_�����:]P��s�nJ�_��ݕ�����t ���b��[��H��A��rӷ�7�r�c�i�O� $����6w �s.ǵKج��C/�Y3��1F�D�9\��1gt�|d5\
�����+�.'�,�;�F8��=�Z[o���k6[P>����|��~ ����ߢB��62�e��-���DU�_2�߸��f�ti�>)_j_e}��,��;�B�Oc!��[Zͭ&"��:/�٬����	�n�pq���>'��#���x1��y��Kl�>�	�2f�oK$�йP�bF�1�K���&�ʫ���@r����[s�ٚ~I�t��_F���ބԪ��������~��-���\�]�L���r�m\(2C�i�5Y�6Fi����MG�B~������ﱪ*ɨ����B� >x�Dj�ɿ��O����QG����=P�}B=|	L'��������Ͱґ�(��\���v��+�l���K4fdR�5FSW�TH��R2�u�MN��&�~��n��$9O�����T�sEx���E7�0�+�âռ�,��S��s��e����i�<�V��BV�'��L��)葸�T������:���5��#F*54�U�N|+#s)�����B��T� �1R�-�����W������Թ!�h
�"5��2�7�\߂�-;�`L#f���; �c"��N=�uV�EBޮby�u"�g'ϕ80A�U����~�d���&F�JF��N$��vn��H)bS>��i4ď�'k�yŜP������Ϟgv��ߍ�0湶�ۦ��JR��0��Bv����Y��U��~�A|���J�S���t���]v���TغWȬp�AP!�zn��kf��+i���ҷ�4���� x�V[r�>t`�b�E��fo]�����B&,*fA��ˀ!|4��	�eP�^-?�m'w��C
�$��Ʃ�n���5�����A�T�g���R�Ci;t]�f�+�gpa(�U�>6>]i�k�v�:��g�QZN�߀N�'�-W��?���*30����0*�����+M?����%�F@��=�>)�E���-TA�(I�����
�5$c�8�_
��Ӂ�x�"��Ǆ@�ZMV�E��W���W��̟H�qAU>(�/~C��8rۦB�AH�ᚺ���h����B��"E�'1��S���%����B�V��SQ�+�#�L�91��߲���Pg���]Ǫ%Ȩ5|�1��̯C�-���yu�F���a��D�5mN��R�N�B�8L��ǐ�V0�LX4'9og�0p�L������V��E�Ā u�*�-燡U��u7*;�ǋ�LB}�|Y�єm��������ȥ1��<3�Z^�����(�`o��K_a{���
敩Kiװϼٻmt4{�O��W��A>��v�BI70/^A4&�a��[=��?m��4���5.J�`Aʂ(�!o�_S�Y�km��v.?�z0$�'�r]�}���������l��(,�R���!(I��UM�Id����eD6bF�W�]�g���}�?'�Z4�T��'�NQ��K�c���s���"ӹ�h�d�u���_|j��'i��с����(��7�]_޽+\of��1�y����������T��:r�����3I�g���B���m\����aR��,�*,W��1�뢋�Ϋ���
n2�2�	����i�;�NⓇa�W��H� X��<��	Ernۉr�T��HA�3��-_T��}8�;�W�'�^WN�̧�W�tV�����Sx�H��7�)�m<y������k��y]�,�w�ʂNQ�����"?\^�͌����p��3h�4v�
l���y"���~������dk�@�=&&+����pC��s�sR��P���E���������ӹ�sE$X��p�xV�J�t��y�"�t�N�47fZ��3����qF
�����Մ�X�ô�X���&�#0�w�Ā�|�.�(5���J䀸��Z�9{���{���U����ن[u��v�z�d����@�oSDr�ns�ܐ����P@����GbeR�;�)I�+>�?ڹ��ǚ<xI�)s�~����D��֯?6쇊F�IQ. t�=�:�N�>��{��߻�s�����@]��$�@	��sOE�Z��8� :�0�Z�C��[��mY�1``7��&] [����5{���7û�=�Ht��BI�9�V��K�����S"w��s���#���rQ�#c7{Ev�Ⓖ�Cg�q�|$'�g%�~l�9��ysHJ��m��WD\3c���,)-!��2�#�8�ό�-��.�S`7XE^_�ly�	�����9�T��X��a#�fǴm��o8���[�~�Gl�0����:J{�1RD��H��GP�%�|�q���;��ÿ�kg�0!����z�o��X�PΎ���Ft��z�B2�9É�5ٯ2(�9Z3>�_�T���k
�-%����+��5(3�������*�+�h¾}j�AG�\)դ+ڗ�Ê
v}{/��r)��M���S�� �HA&~��C*%��v��̯8n�,���B,����S	s��'&��ȍq���c�Eܠc��&%/���!��`���o�3of�TSJ�b�����we��(����)���W. ���ՔD��r�:�-�z}�A�#>����+�hN��?�"��ژ�h��xZ�tTa�|蠀������Xnmՠ��迖��D��V�D	�˵�d���L��r���ؓ��v��� I:y?�ika�KwU�V����>��*Ys��!zK�<}��z�Rx��
CI�Zr*L��-*@�A}�?��02���SSKz{�R�6�yV�g[� qi��@��J?��I�p���!m��i՚+kq�l�E��i�ke��R�Κ�&�.�'{���M�R����-AV�"�6��(�[³8>��\6\���̗���y4$�g@����)��&9�+�H�;O�T�h�V��UcBQ�pm��=���){�ti���'=X���"�!(_�V�hӢ+*F��b��0����� T��^�oz0M��+^S�?|�$�	X�u�Nb02s�ųX.���=H)8��DLr���x�jZ#���++�I�����[A4��T�I���ë�5��Ie]���ٯ���9�sp�[>�3:'AҖ� ��A�,?�3�$����k�r䅬as�S�a^����@��0�r���d�B�As�1�ʱG��ςZ�H5R=:پGPs���l�xgJ�fw,h�T����R��e�����X{tɀ�
?Y?ɫ+0�إ�R%f�!K�T���	f��w�xf>����UM���yo��w;�Z^S�$¨<�J�^�����])��59�cyE���Ē����#f�B�S��"��3�`�u���bH�=ܣ4�m�9yB��N��;�J��q��1���=[&�i��c�XΉ�3,U�p	��3|}�4Ia�W���p����r"?����ң�2o�9���(�7��V��1���I�Fc�#�R�X=�����f:VZrC�q ��|���i�K����@G��d�Q����k��e��Y[� Ϗ�n�V�B�nŏh���<|�������)�5H�J\���XW���:dR�)���T��S�,�*���>�0p$�6�G`�`�n(�0>��p(*�I*�: ��3��Ma�#
��U�i��g�oa�7��1���������Cڦ�"��2i�y�a��ەD�Ƴ�Y��&����hw&ێ�t���h���3�q�Gzk9,!y{Ą�4K�KU1l��UVۢL3gR��A�q$7����˄�*��b�޼�J�]����=X�f'�tfL�֊�˂��;����$��8]��E��U5S�CV��[-��W;{WY$=��?Br�īA5�L��̷���P����ʿ�Vp���n0\� Θ���4��2T�lYV�z��P�;���èl�v��gp3��^��%Hg��gϗ��i�,4b�N.B7~�N�/�_Wue��#���,���� ��Lk�Գ#1$����U"7�UA���6
�����Y���ds]�;�+'����o�y���8|)�p�4v�3��g�	s(p%�n�� �WO*�4�l��,��#���Ai���,�y���A��i�"�����D
�x���tM�����Ԍ���ei�R�kaǉ�B9���y]T�,0�p�e���r��3��ߕ�	���~�v7�wͿz���<=bl�5Yeu�xR{��J��w>y�{N�>�&-��Xٖ�Q�/������ ��S���I����p5�G݇N�!2��5PM�k���{�z)k��*#O��b�oW�خc�4g��ۊi�ɾZ�����Pp�`h���@K<���O�7n:��5?�Z�O��,U��^v�|V��KPM /��s��Ogc����i�ݏ��!w�����ڞ50J��0��tʌm�MO?~�N��3��Oo�:�Un�[��`�ݮ6�ǉא�dr%M֮�����y��e��de�:GIl{�lu���
c��r>f[+F����>�j�1$f �R{��Rϭ�'n"8j�-@��.�
�}��N���2�ׯU�f�j�0��M�;���0�t4��E�pR]C�Lm`y���[#���b���|;t�C֚����ZZG(^O���|�:ErBaU�OXH�*3���ǌ(B�I����N��y��Z�,l1lJ��z*��0��\/�<7F��nAlarD��F=��x�R�zᩝ;�m޹�C�
�}�R����2Kv�Q7�?	�^/� ��h4�x#��3�.��a�S����X�����O��w~ݧ��+<�m�d�ϙ�J�(��2����n	w�ؒ���K���a ��rb$nؑv˞M���F>��͍�W�>�wa�RN��u[ʰ�qd�˨n�b!"�����l�V͜�J�Q��k���x��ü�����ވ�ԶS�c�a�l�����kW:���|��`��q�Eԑ2�_<�
�\�1vJcc�x,��]J��$�Z��CF%+9D�.�"T1����*HR@b凛��
�H?A�r�,����7���V�Bd�V+�0�S\~�(�T�Ch��s����:�m�cW�0�:g�����j� =�"�Ȼ�+P���n���w�)���擹�NU�Q��C�-��8.���N�Rj����H��!J��Ҍ]���������vL����_!??t싁{��J���z�|����zO�����&w M_�!����n��E}��IJ�݁����5[JP�Vnpi[��4Ȧ�0y[{?�ʦ��?�J0��
�wnܻ���k[�2��S�pj���Nd���@��4�����Q��"��^b�>��dh������Qx9-q��˕s�j.Ow��uɠ��]���A��@|���U�t��ޙ%;�P��e.�m����9 �/��O�>V��^�1��&�&�o�1���<7�z2����nRրZ��]�JWL7��e�[_ç�P��H��ZI֝D��01[�,Q,�[ښ@�j�u��|�p��p9]�
�\D��R$����8�����=�UT�I���`U�B��q� �]ۥ7�'�{���c��D���kݫD
�I:X����c��l��v�� d��+>�s�/��aH��UH��w6:�/q�2�~�YG�����'���0�Vt>�U�߀P�����d#��)���	XVFBÏ�*GtXD�HP��1��?B�1�ȟS��oy���g��ʲ�F"в2�?}@����>��t�j.A�����G�5�)dX*7��hr�ʫs5�'�Z���Ї}����	��~+��n�ř6���ކ�\Ħ�=��3���u|mr���(gDc�8�#��$fJ�앂�g�W��9���,�H��a���y�@�X���/��/��=�z ��n?qz�P��T ��i���"�������jB�� X�����S#,>{�,j��N�St�EYb��귮�u�~V#!9~M���&Ou�����}Ra��d,(62�^{�5W�ԥ���ևa�������`{țI?Y�h�1�ް��S�&(�:��r�2��Ƌ���_���RqtTM:A3�#l��ޤ����>��!�ԆT���|t�Q;k����ݫ�]#Yp��
�5�
n�A�K ������H֋J��|��LM���$x��n1�P�4�N���1�Ҳ��@����h�`G�������ъ�����Ty���7!�³q+#��]�?f����������r���
w1�)�� �����o����S��L��#��u�qX6���ٙ��XCB$�������6��sX�$�B��^�r�6]#I�����=���o?�����#�i�}�ߏ�P�[�b�Y����_�+y�o1�9��Ɂq���c�x8�D�����$4+z��?�
)-X��`�G�aቤ��W}��*���HB��,�4�<4j��ab��:fo�^��� ��;�I�5܂�y_��gf4q�������t&@�,.*�����Q�/	�ky%Gc\ɣ��u3t��'%
��ǜ��D��MS��c�!��3G��\L	�Mj1����Co�A��2�<�9��D]��B��oQ������ⵋ|�	f�T�C\_����O{!�=����ݡ��,f<����n��]�{-���y�x1�l��DZ�d���z�o���n�LM:�Y椠 :W�)w<�V��e�`����Н�)��'a�>������9�RJƶ�+�JYN�
�DS'�D��z�Pԃ`]��Kְ�Y".��kA]�f�Ga��	�fKa��f��뽟��������f_�w(i�([�3pQ��Y�1p���(wiȕ��@v���1@�IB���7F�b��D�0\~D��3c��ګ�a ���3��@��!W�:c��6&�m�I�VZ=t�ȟ��H�&��K��%vSU�`C����Q7�:��tض��#�vP�#�:���+&�[-ԏᏆ��ʌ۟��$�?��!Mڔ��\�-����������'%�疸��l~w����'�!$ӫ}	q�'�Q���]������p:.j'�U�f�m\I5j��㆔��Q�&�9�hc�Ǘ���E~﯑�O)O�Pg��U����60�	����GX?�����b��^����#GAT�y�=��¸�pMx�F�Wi������~�o��ܚ$�>�}��š	n�^MunQ:_�B����U�r����q��-ϐ����<��y�6�� D�}����1L�v=���9����v�?�/W �	>yL��h`��@e�W��IEZ':s/���1���&�Ό[n�����<��fr8�����[�5l��ED�Ov��:0�r
""S�6�mG&������ �Q:i�|��e�O�c�mȷ,�F���I��X<(|T�5{����a�H�p�Fs�X	M�-�3�����7x���O2Iʏ�
�ʨ��H��\FfyF]����T���+)7�:m*(*���A��#e� ~���b��SS��ZNo�j?�9k#_r��H��˴�γ�Iwrĩ&�W�[w>���.�m�o¬�I*�4]O�%a.�Х��t��i燒;�� �y�P��ۉ�.k��m�ί�	��tY��o���f�H�`kk����qj��q22���ЃY'�wê���.�p�ٳJ7�։U��e�ݹ����Ԡ��|<�B�G�Oh������A�%ڙ$!ib�RP���<��A�CK����t��и-�`�H�*m�6��ɀ.cK�lv�����]��Ws���2�|Y�@s��W;fD2T�P��.�S8w�;�n����ܛ�E�bt1��EU������E���+��!<P�Ĵ]cf�!/�x`41NO�A�σw'�e,��v�'�a<o2ބ�,de9Qaj�n���P~��
�0���j�p�zW<��t�jC����Ӛ}�UM�،cWp����@���z����t���54��G�1��)o��/S�u���K�|�� u�X�>M�( V�H1sF6�WU6+ISR�~�s��0��3�㥳��K��(���*��aI�e����T'���O8�@"^�Ț��g_��q��w��$b�^
^�2�ZG����#x��њ�؀����%���M�0�ܶ�^��$����]�\�0οW�����5'Q����r����0߅9%F�ҵR�Z�� ��9ϰ�1�ɃU�B1�4;�Wz�;�^��i�(1��L�]H�#�}[:m)�-V�GH�i���3V���_��a�0����|bí�*o�B��Rq�VXh&
.j�s Տj��pŘ��T�3:d}Pl����wk��5�����y�P+�BKta?Y���?H��z��d��<��Weq��\D��(��1�1���Ҡs���'�J�޲��^L�A��O6�WwK�}!�+������ً�>q�����"�eUB:�:mT��f�0�ك*�\��J4���Oj�����\�N&��?t�â�t�?�h�M�i�!���~�2�d�A딖�?{t�O�t"@����i��WKhKBu0�ȶ���s#�|������Z4����M�S�X�-���)N�Y�.�.�B���x��?����P�K�8>+�r4���@�Gq����E���k����ۍU�~/^4�,&3'�:�藸@ai2�쬥�%�C����LIz�_�ږ[
�*��{̟j�[�l�9}��V�(��S����E�s�B����N$�JLBb���5�s����P����w~��җ�Q'L�Q��CO��;ʇt��.���2�4�fM���A.!����W����g�^ ��R�X�<�T�^A �暖E|�fV��2���r%�^��qL�0\�ߪ��9���gu���!5٬J�v����ia�8d��CKjN�ԉ_Wi�!}�2q�Ծ������<;E	��ؽ�m$�9�F�L��"�7$-��_�'���cT7�F�z�l��~���1ߚ��F�cg%�`�'�7�������N�J�B��h��ꣀ�R�RqϦH��%u���p'�Ͽ������!�ޤ�`}�bQJ�xu��sf�F-Fhd�XB���j�UG!%��c� H�h"�-�F��s���Ȥ|Kj3�Ż��iU�f[�51���7�@Z\՟����6���7yϰ�}����MC\AT�r��b�|yx���cd�bԤ߂�L]�sY��q��a&��ˆeC#*lN\�5�$�W�{����\�@�vT����Sb���ا����^crF���u&�e�x����ʊ�\����z��&�㲝m	ф�)�B�>m�=�%ҧP��	Оh�(u&�o�����J�-�sW��Q���ˀ��}����l�L��C�s'��.�6v�����nD��>��s�F;�w�{����q�z�1�GH�,�����뺫/ՉC��EE���.q��tΦ���;F{)"���gM��0���E��`,��K�:/p�̅P��1��p��#���8� ݡ����C	_E
���"�,�qXp�S���G9�I��-�va}��z�I�7aȰj�
�˽��<����T���6b��h]//�F���,h(�Py��hǡ���`��(*G�7�1� 
�	e�p >�V�����3[�s�� '@,��<#[�R��)ã�	,�z̃��/��;���n��N5��P�R3��2�q��嫓�)ڽ�v��Z
mC*BV�xu^�n������襛��[X�8`<C_2n��C�[������R����{�w�1��|��/]8g��Σ�|���uH�m��S8��^�Su����������{�Da8����ª���$w)���!� f�7�y����;�_�̾fQ��Y���������kj�l�:���ÓC�h��ۓ5�,�ɘO�����G�)�=Ȃ� ��N�ќ�������AQ���7�Lm6?��}�����\�aع�b��D�V���$*3 Tr�ENF��|Ϋ�N^��+>SZ�%QP��J��#b��22!{o|��[95ʆ� ����pKF[�����`����x��N��Ȉ0�3���g���X�`�Gb�S����dq 
��F2ü(��I���kiwo��)z��jR�)WG=�W$,�B�l(�Ģ���I?�����jq��z�>�u���t��o=j�L��}X�qT>�2wnD%-�l�F|�W\��ߏAM��':`��/-�g�qI�ֵ����c�
d�S����pyz��w�u?���|<��ɘ�jds��+0>�O��9����I�ׅ}!:�I�n �o0Ls�j�qm�x@v�~Zۃ�-���]�!p�Z���C	��R�)C	��#�sP�g*W�i���<u�Q/C9���#a�[F�dW酷�l�5^s~/[L��n�}��W(���������ȨIB#/[�A�/!�/I�L㇩������2/��jȨ��W_���s�Z=q��pY���5�)/�]e�w��t�w�lQ���~�/�xJK�a�éM�K�'f�E�n�y�����a�+��U��y0���Ѷ���'{5���:������oeڱη��a�?���f�sG0��r6e�d���2�T�ƊM=�I��A�X��#�CX/�؊M�e�X��`���zVu�(���ݬz�{I��L;�>��ש�@�~�^��`�9H�r\c���� ,�su�������A�i�5~�b;�KJ��VC��x̨2J%t�`d(P���C]�{Xc�6s�//��O��Cyi����H� 3�D�-Ȗ_ ���*���r�����gł'W�1�c0>��(w�٦l���W��IЭ�\���R����Jñ,M��4G�.����T��c�u9��Ꮙ�k�h[� ���w��W��i^?]|��+GG��
&��g��*PaU�ۢ�����IF��&���,� �dB�) ���n�h�J2%8+��e$�"��Z(�
_�~?r<2ȸ������2�L����ٶ��Z����lp��:ر�Z�Μ�6���U@�M�1H��
T"�r��Qe�ٽ15�����}8�.W����Io��MJ����f�Z�/Q�3&����Vz�1�T�l"s@o(FCCc~���rߠ�z���
M׺��Vt����K��G�I�=��Xwbc�&6:�%Hɵ3�o.�a�p�;֕�9�Zhi�����M H0�Y�c�����@M7�B/�d�_�q�|���	�ߧW+�<����BK�^;!.�eq��Dv���ŵw�h�_J,��/X'�̋�I��*|Y:c�Xr�E�:�O�T�1�!�j1LT��"��FVߪ�g�o��~t�6�H[����Y�#��O�ߐ���4o���J+"m��/�^�[C��˩�m�$���h����|���CO?!z1��8e}.��F�v���Ff�*���ԋ(SS�*MϺa�޷`���	�;���c9�D�6�U���G��O��u@L/H�|��mչ�G��e��p���2�WH�f�����b0���nw�P��J��_1ڀ���������C�Ȋ@|z���nI1�Ɵ�옖beAr
�� �lWP��8��tf��;����5�C����V���.��-۪��X�zX�|l��+ ;]���i��!يc�Ԕ��ʺ�ʙ|�b!�h.Ã��+���t�o�TB���r����!aIkMS�O}b*�5� ��a��DIN�!�=5 VXP�+俀D<�1U�N�1F5�ZF��n�������������?�J��"(�5)��M�S�9�^'Qn6�x�AXcAz��~�yb�/�I�}-�I"���g�/Aw�&M0�I5n�y&��Ք41Y��"��`N޼�I��٪:����v ���\wY�A���[��}
د��P���5�]z�Ъ�g�}�#�4�$$5��R�`�	���ӱ��M��_�r���B�0E��N�c?i��仡T���M�u?>Z<}�� q�\,gO��êǺ<'� �O��E����-��E�b,��|z����E�8�m	��?�Fikb�W�1�����Ǩ�����`�އ����4E�V���L�`/����@P���z�`�d|��Y2'�v��Qi�!��C;R}���'Ų�׿��L�P���S��T��l=w+���g� o���5�7����J�L��dh�;�c����p1u�KA�#����/L�`T����K��YJah6�卮i�c_�j��pA?V��)��&�C�mL�&����ͻ�n���]�G�QQ�MP'�V_���*��#�
3��S"��8!O_�YEl${�C��<�+Y���.'�B��0��/���|�E[�:�WkF��c�����!
_��B��eӵxIc��c��v��zm�4zL�پ̢op2��d�)b�ʳ��ò{�e�1��:YS����V�/%^|��,�<�:���sC �R�����x(�H:D/��)�vspy���_7���Cv�9�Ţ7+�J))������vџ�����o�)k�h�#�w�o٠��L:�y�_��y���3�s��������"���P0Qf�<��ŀ�	^���
׌��g	/��6�2I��΁�b��I��8�I�x�2di�8{�ve(��J�~�kｉW3��)h8�4��I_������Q\�Ŷs�X�Cw:��R��Ǌ� m��ܺ��%_m�,�����V�> NUAoL.=�g!?K���V�x=���q��#zf�s��`_г�I���5
`�J
�%'�/� �5Gl�{���"1k�s���/�/o�!�|�D��0	��~_ֵ%���R�vN�3��{V>}G�SPux�B,?4���yj��H��3��	�w���F�9�7y*��_��<[ʧ���g��=Q�����ko���ʐ�CCxx	;ݗ,�W���UlY;J�.+{�6�|4����q�Nn:$��-���z91�	��\��*��ʎn�ɟ����G�:��4���8C��ϧ�
���F��=�jЁA��êԍa�Q��]�0�d.�TL��/�Λ$�!�vΤ���a֞?;�O�⊏Tw4 �!������?���<Z�Q��]���1���]\ڗ�X���lt�@C�e��$�a}Ri�[[�����WI��4���q3�6����+ ���{��k�#ͱV�t�r󍝻�+Յ�>/x�k���;X���{�C�a�Æ���@�G�����6~� E2M��N�<𼁟W$�;J��i�U�L*��E]`������X��D|��Yxuir~�c�YrGs�6lc���
�T�
��8؜F���ڟ�#נ��`OF�y�����v��R<��&�4����K!�5.<$� �\�1�\�5��?�vV�4�9~f�хbt�����l��ȇ�����[�rg��,�bsb�tQ?������
q�q�#�
=��a3Y�y'��@��A��V��v�1�m�wurwcp<����2��UW�*���͇o�}��Ə�xnc�B����ȼM>�F$�0Y��
2g�����?+���Z�������̈�kN'��r����{*d'61%穇wJj��f<@
7�>'< ���`�B� ������[��IĘ�_�!�&�<�qǣ'fN(�WF<SP�Ԯ�l$3`�_J�<F5턀�����Ψ��Ƶ�ɞa�������9��K}�F�	����{y~F2����^�)��W��ڮ��ʎ�@p���s�*w[�O�#�C����	V,�j�wM�2h��3M������wl��f`aw��O�d\Jz��������T�V"�@KZTx}?Qd^+򤹃9�AM���m�|�t�8�F��-���u��[��L-j��A��d��	>�Q����Beҹ� 	>�Io�3���C*r���WE��O��x����0:��p/T�T�b��t�m��ހ�v�j�?>O��W���g�䭱@���:���������h.~�j�s�}<�5h_��/��mg������61��}��F��їN�l�:���lߝO"/����
����(t�\!JC�����YK�=�]i�^sF'�O_���U�~�5��&e��p�vࠇ�i��ī�����9��?�^�z��*9�!(h����e?<��T~NR�����S	�b�� �2�D����V��=2v�+iZ��E��w�N^�����ЍmǛ��'�&aL�۾k�"��)�����R.�޵�絀��qć�[Q�)���n{��-T9���!gU����t�\�7�Z��ñ����ĤH���9��"_\����Ѣ���<� D��0��g� ��✘�Uiy�x�Fą"���*ʤ|ݬ�2^ �$�'j_J���M8#�q�,:LT=�ACJ[�G�_I(}Q�4�s��U�*�[��FP���S�>z���qc���`Y����B]�#�/q3��7�8;���#r�BW��Ѓ����J�|xi|�T�k+�!8�HOX��1��������d�g�W+!��e�l���f��t�����>ul�?Nn���U��W���n�m' �WUػ[����7�s�j��1J�ȉ�wc��(���W=�6�B��ٳ�я2wX=�?g��L�\����PAe��SJ���oD���Wi�7�K
Ѣ:J�4��u�j��s =�y�eQe�\�
����"��MA����c��Ea��^�wj�1*�Z�eã����3����VdZaa�H�s��Kr����*-�Ǩ9c+4�0�<9��VJ��jZ�O����~B�sA�Z a!��Z��\RGE�/��@8..F[��8սf��pW/`q�Z��NI�5��+)\1�o�zi��2Sv�ⵙF��?�1�|���6����;=����CH�"��~��)���K�ByJ����5�k���G��A27����k�gz�[��S� �W�"Mn��$��EF�HS�B��Rb�~o��<3��k���&��6>�a;�d���i��l!��J�)$�jzD>U�\��&׼5�{C��a���Y��Y0�8����8-[�7t��G�$�E%:B�6�9?��Q蠑b�jF����z�x4���1	@a�w?��W��/˪����W����25R�azTRn�!P�.WX�:#�0w��b�4�=}P���Z���xH�nq�^L���\4�7� @�����.r�D��[�jGj��-IW�6j�ߖg�!2?'g&g���2�o��� ]��t����^�	v���ME�ud��;���U�/?�6�0��[��D^��%�'�)V#Ro0x��=@p�������>����u ����"^`�&FYԻ�<��"��Օ�m��@���$��A!b�R௾/�T�$#�RK;�V������	�m	L:B�O����.Y#'
�-D ���P�Ԉu~��Y����d���1�{#�1�Э�q�_������*��Fq,p��0�ް�����y9�M�a�M{q��|��衄E�&,oj�"�m�[�7̶x�94��������.�8i|7���f����O��,5���	��.�����x�R�L/�R�����q���a����Z�AIg;�jx�g/-��,�2&M�F7R���%Ҕ��T��g
�(��W��-�h^ϖ"Lx��lȉH���.�z�T#���e��C��V!���dY�r��D=����Gr{�&����~�
�s��)����%��q��K\8`���J˄��zL	T�dm=�2?�Y�ə����u�t���f9��`bj�}D�t�h�z������]�1�z�g�Zd�I2���;�萴>�����v�f����II��ĹR^Z�n9k�mj���耧�"u���_�ޤ^�ݫи��}�78��>��-��Ƅ�"��)1̓���^���wSiTt������Wj]2�M����iXd�/�J��K7�ٲ> '!Tomր2�{��g�b�G�H���ߪ�ծ�9�4P�po�6��saO{ �ޟ���`�#�����OssE���M��d!�K�5�n�@l�5;xܗ(">0��T�]�����> ��8hɏ�A��&R��+7
��K$�a\�8����B���L��4�u���bz��Р�i��%h�"4�*�|��.s�v����P<��чY�g(H�i?�W��Z=��"7i��
�����P�d�O��Nqs���/hx8 �ԩ�}ބ�����	�(y�As�{ˡ+Ď��#(t��z��V�Zka�'g�������t������R�*�${h��]g�a?�c��f��b��E$X�rS��_�����{F�C��:~79Ơ�A��\~�m������r#�W��B/��Z��h7�k��X͆OE.wF�ٰ���8��w�Jwl;�;<{�{&T8�lps2L87��B�����` �W����G�=ԾzG��gZ?J�P�SxNٵ��y+�P�b`�-2{��������� �yΗ�ΩA���,�OB�@uS����u&���eh2��k����"0c��Dwd����aKo�"}__��p�V��-cKWҏ@�u36P:�nfɧͫ��0�ڇ���L~���y{[c���V{����	r��Ö����{V�K�@�Kww�+U����Y�����s%��7�M���"b�,�����;��~�)�u�XC4�$��!�.7���{�Z�߼l  ����zCv�>H��g��d4_�D��ݺ"�?��mw�@�|)]WS^��L�2����X��wj�����S���n�1�
<��@5O�����4��U�U�`H5kN�(�m�
���kG� �(��~}���G�r���D^��|�s����GY%X�����lDSJ��cz���Z6PS�w2˞8�93�u�8J���
���jK��%�G����	�^�T���|�~�D�S_:HzG�K0�{����TѲ�>�LhBZ9[�m���_����o<��ȩ��cD�����D#D��2q`�(&�k�6nSQժ)J��
����(����>Φ1R��^d�@E�~Eӑ�pz��D���7\Ac�R���<�
q2�0f�t��\j�i<p�,G�yB`��2G�T(���~x�i^xz��8��	a�!}�E�P�{,�o�bǘ	���t8��"�@�����DޢIy9�
��®`?f~�`p&�n���ivO�3e�`fh�'��i��ڜ}��_�%d+H:֡���%2��̤E	��*�$�`��w�2S�TC�*����x���?���ѡ�ro
<R�0Xu�Gx�,Ъn{��*O���+�i���٩����:�<�Q2&a�B0������D�s�R��1�
���{�.��pm~�O�C��� W�-����YFj��7�x��9�	����;P��c����`��Ha��:��2>[QK�x�������[��Mth��߹g�I9����I��-{�q���u�l�Z�;fd���r�|(��(6N�|�İ�T5bRf,�@�P1C�L'a^+v����H��K�qܽQ���Q�If�6�����h���b�$A�	���+���{�`մ���n�_�n��68�k��5mTہ�L���y�!*;������Ҟ�&4�����7)0b�����[��Zl�G�%*���-�)ȵZ6�}0d*:�GK���bId�Qk}K�8��{����]�W�a��I�q���+�^��%����!u�=���]f��) �
�����8����Vz�6���%��J(C��;P� ��C������\�.ۯ�N��1ti�M��C�
k"4����Ś�f�,5I�m�X�����҅�����w(Z�x�|��!\���,�X��3b�T��G��}����O������K<y���!��8�SH_%cC��)^�;��g�0Q������:1�ӁYG��sӻ�ks�{� �`�@��eMֳP"4��9�䳶��3F�Vv�7���m�c*>P��'�'�U����J ���y��6�eq�[WR��W��-���:݌ړ��>(�K��]�r|����$+S�h��58�6`�ˍ�զإ�A1��Ϟ�Ȣ��1�ՙ�}5��)��-���f-�i�1(j�-e���R�~y��,���e���#5�:`�mFEWH���<�)�'�9��Z_CB���� x��:e;Y�/��_������4�)�̞tN���6A���wN̇��$��)|�K;>�}�R���� ,�_W����#m?5�,]��$�ʋs�R����C7��3�
��@��.ES�; ��Fh�_Ɠ�� xc^Z!6U����_�1#P���P8!ziT� ��֍�����a2b�ѣia8Ƣ>[tv��B��|!8�h��R��i27L�F�Z���f\^�,�c��/�ux�Uy�ac}fy��� �9����i�v��Tg�R�C�U(�.��fs\�u�Z
^=Y��V2��g�Shs�����TS	��ra�.�#�1E=��{{^)Dh�Q��1��_^�j6'�8!]�藶
�S�k�ʝ���4�!^x`�h`d�b�-_��~����Q��P	�6�p��mX�U��S4�����S��cGGe,�j��R���D���h��7���Ζ������ ��ԧ<���kc Ӿe� �]H|�&Ot#� �2�K�ʶ��2�榄,~�~�8��8\(�'�9a+L�XZ����+B��U()Y}2Q�$�3�;c�u��PJ�Y��i���yj��\0La��'��H��$*�ߩE�%.��c�'����m��Ma�����|�i��d�`�Ω�Wkc��\�����ƻE���F�HB7⛙dQ��;l�!�2��0���4i���`��&܏��F�^�~��@r��[��oD.�e'���8�b(yVm��]�1uV�\���i��1cG_4�c���,:���U8��'1��4��S* N�,!н{�G��:���H�-�w�ب��`顑�(� ��	DEh��2^� 	�M��]> +���6�נ��Qd4,R����3��$���.���y�o$���(�טsJ�Nu��-Ϟٶ��F��Kb�9����r�"�*��b e.����8F$\ؠy.)�Ly�,f2���,/+�Hۑw������� �kP$��B͟�׹?%a�3J�W;��1K1�Vd����n�/9��Jp,ˉ�c����Y�,�{�b<����F�T���NP@�>č}�����E���֟ C�r�G�0�/{��ڽ�+8��H��jR����<a[ǲi��x��G�\ a�M����G�Q���E����6�,�F%ߙ؟�2�
����B�����-�NzJ�iEc��B��UԨ�ʛ�������uI��u�x��1����}_�(#�g�;MpY�l�<Ơ'�u_�0���f/�ĝ����9M���F�i����l� �dqp�?��	����o�B���� 05Ir(���>t	�(�Xq`:|/r�<i�Z5l���2�)TlH�2�9��+T�u$��UN�0MMNב�����@�;o��EC��&`Y�?`J�I�`�ς��h�sn>l`�?#�R�da���Z� ;|�x�;:�������5�F�g4�">���i�s��H�`��S�^�;E��zDx��SRW���jQGTq)��$Qz�� `���ì]�g���خM\X�-���C��9R�G�@A����u�W�"9���D������anȬ����<�|�]�#�����/ޜN��Gͷ���|"�8[�0�Ё2��l��XUP���{�f!�N-B�n���KE��������џX����ID��_�"�6�	�2�gL�ˇ)$�N|eaxI �Qv���RXmE.5��A�".G��/8Db�����s�:_2ێ�`��ꮤ���NfL͙v!�{�	SC�@������F0��5VA��l5�=���o@tW��g��͔~tXZN��:�l�u�G���B�DsP}�+4�7���D'�����ifr��2����"t �=���J��ܧ��M�B�����/�|�T���;I��J�������%DR�d��7��-L
�2S�sl�H>~(����zE&Dd�A��s��=����'تve�+�]�g�Z��h?�+G��U��C�2�]g�H�^�6���M�3T�8�����<$��+:j��#�Hz���W���h�Y���Ǔ��5�>e���_GL��|Q`)�ꙙ>fC�x)���cE!���*��ι���KC}�\�d�|̘N��p�ܜLE��a(��0��*�d���zk�݉���= z��R�4\�֊>{E��'�b�S\����;r̻�^4t=Cp7�郏?0*��A�=�U�k���.����0���N����q��>���(�٬��l�]�a#�|E��Ţ3Z����>����P���������ԯ�W��\�k:��.L��o�^�G�^jW�^����$�H��)�A_�X��e&��n�ӹyX�K,+�.����2#�h���D�4���!w����V�>\ܙG�9]|ď�YsƖSÂb�zL\�b��0e֒�����G������q�o��@�+]_��9�#<Rk���X�|�g�BP�	b��m�L��o��7��[�\|;��Q�Ɓ��4�T�����X�pt��u�;�w;{�+�<z�@�gvt[��>�0l��8Y��"��(�wF�P��l�2]�c*�Bv/�p�����ઝ�/�ta&2��n-�A�'H��=��CE:��@�bѳ�:��bfz6��E���#
� ��������#d%u�QyF�R,�o�LQ��T��ts�e\`'4�2�Eךv�*�e�7{���L�Z7�o8�B��z���qΩ_bD:��Sy�}�+��_JO�@���]�#����������Ƃ�� ]ZM��V3e�bv'���&��C���	�8;������ަ&�&�Ɓ��z) �X��R����ԋ�u�.A�3:���3�șz?�C�%_�ñ�m�>�N���%�A�&���{-�_����}T��N[���� V�<���ɗw���;�]�.J�<+�WC%�2���N X��`���(qj��UJ
<��(�_�E�͌���{��/��N��>E&�\}�v|j~t��m�����j��*J�k
�:)�Z>����Sx.���3�'7��ǲ�%B�Jė�[�v�pC��*�`6�Y7<���c}��V�3��}|A�#�H���E��	���	]a�|9���_g`�d�ea���[^�a��v���2����?�i����nE�AN���Q�F���Q�@�{���D�<I���{�%����Gr����Cs��^9�g�d����
U, ����
k)4*Ze9�����ۣG*^����--�+��.9D�I���XۦA]+6��dmYk�W�r�p���=�_��l(�����8Ƙ(}zH<���Ej����^�j~]�Y6jp%��_��yg�ĥ��߮v-*��
�u#� �0��p���:0���6�����.&WK�U�'H�|*���ࠝ4N��Ձ�g��[�Fo����Ø&�ҡ��V<4H�L�<�����5T0}>��T��7�([����_t�Z<]sͯ��m�I#L�e���ޯ:P��r4/��e������6�곝����"-K��m�%'�l W����W���U����z�/'��9Ν��§ �v�	D���>y�r�ޣE�`�|
_���P���)�j#���W{.���	�?�E����W�C	* N|��y.�ٚjaA��b�{�����l�?����vH� ��/�Rulw��Sc@eOV��ø�������	�{5��bB�˕�N;y��j�N˓3&��y���lޒQ��qMVv�F%X���Vu��N,}	8L�Qp?��n�Jo`��/;�'-�y.φ#�P��K�W�(Xl�Ԛ7�Ip�ёo�+���T~�%�+IZ�ˈr�*�K��OyX�D�g� ��\�%�̽��ު�"����b�h+\KiHֹy�1iB���"Uh�*��a��p�[z�Z1��%��τHcҸ�Ѭ��=&Il����U�z�?|��1�ZhpdU�5�?+�XYi���O z���ʥ ��&� �w�����m���!.m����ǁ[x.0T>4v?3�6eP/��Ú��������3T���
�]%4�V��ę���"�j��s	��oC=&I�}����qc�Q蜘�g�rܼgz��Rl�F1���b�����o�|�N�l�� GN_�$\b��՜�p$��v��s�.y�2=�x4�Wԥ�l� Q����;#Gڀ�LJ�c�"�����Js�*�J�b��D�Fܩ}�H��>��ୈVŤ�/���\Q���P� �r�<<�k�6�Z��p)�α�bt��+�@Xȩ� D�*�dV�l_x��`����{c�������_06�C��/�5�g��Ԃ���{1$Sm-5ye/����R�c{��O���cu#튆���2�2* �T���m���;Q��֡M�W=��S����I5��������ʪ�%����l/\[�k��@������"a,\D�/�O�wa�ʫ����B��ǮI�QJ1^��^��dO�Bǃ�𤩞{�Ǆu�Ҧ>�Q��е��Nr!z��C�m{���)��� �y<���4��E-h�eqO�9Q�h�
t�%�q����jJZ��t�wQo���rt+E���л����`Y�p��0�սwz"i�����b``�'u���\��lkLq�u�S{\}U��{v)x)?�.����%�
��u��c��&����s'�%���Iy��{�C 8���Hq�f�'����������m|6�:z���Y5&�ntI���K������p �֋�r7�6��86I_���!�����;1^�J�܊�q�m��_�/0OCFG@�C���9ES�Lz�ҥ8�m�M�X�|�"å·�$e��јM;+���fL�NT�I��1j��u�p����~T���bd�����#�r�g̫��J�LJ��"�7���x������I�ͳ:ף�Qȇ�EEJ���~	+#��	�!J��1�����c7|Ǵ��4�V��8������l݅Q���L�{sd����y&Pk˜�s��_.���bkC��+Pd����.���);�>��Q�ᣁ~.IB��)u[�7�����v؅,�i?�x߆�%q�v֥���5Fm��.���B�Z�[H�r7�e��J��wX�_��i�Wƙ�i>!'�����v��[��(H)��ݚw�!d��	�h��8%"D� �X)m�3�y��Gt%���9�6�频�0�
$�*�w�\���")nD�ʭ��!���I�we��!%��o�^��_�,#V�i)_���e��m�z[�Kb�n�A��@��Y7?�.Q�$$��k'8�ҫ60'�1��dʂ��� ^�5u��ivGD��:/Sy-z��_�>��U�Wj���p�m��r� ��%V�-�I��P��{m��2" ��O͌I�e�_���K]�{�Tl���v5��fye.�yP|d|1��6�ۙ�Z��^��-�;F�c�]!-��ދ���t,*Nv���@�{>�P*�B���g���@��y���
ha~(y��h�I��X�vc�{S5�IhET=Y�o���ו��H��+G!�jS�^��k\����_��7茦։j����_ѳ�`E"�A�� �Q�)G���c��"6��=�n������iE~G.�	D�巺<�svG\�0O�1b7��^ B�NZO����_�v2e��B�Й��R���,(sJ=�ōa��܆�V���R,�ʗ�9/����TEz"ʀ���eI|�����Q/���8��诃+�i�^ �]�p=����WP�[/1���R�M����� ��L�
C'�ϑ2��<S<������Ba�8OP-��N<�3a�x�W�̃���Ɛ���t�k�0�˞
�� )-('WzƵa������CX�u�EE���,F"Y��ˮ5�ٻ�CyRD��s���C��&tأ�րl�e�5�u{�Ҁ/# y�$ُE�G�Y�hr�TC����A^�H���/��?����'T�"����"}�����$��c#��_�2���Y͋�?���ѷ��b�D��?�Hp-}jV'�N�[�;�::щ�7*9<�Z��ҦH����`h/�_e�K�U
r8��'4c��&<���b������P�iL�+o��U�g�m�ѺU���[��ʌ�H�%�w��g��=�A��=��0��]:�����?�{CȤ���kɿ�Q�3���$��{�Q��1��/$2�p�V�<���+>K�g��-����)��J8��8і���v0XUju�q���q��@~9�۲�J�X��޹��>����
!솘�2ه���A�A�����0\���``�'�ml4�Qӄ�5�X�^;��/ޜ_(��dpA�Jb�2]�U�����A�����U۾Q���dG�`�k;$~qB�݆Ƹ��V�<�>�̙�
9�`�����r�u�n+�D2z`쩇���^�f�_ڥ����-yQ6����h�7s�A/����D�������i�~���nE�� ���;:��B	����CHJZ(Gr4\���{��K�3���U�[DFS�je�4����5��p�x�jY�n����]^G*����4K�T��ڶ#gS�
�����gmwYh7��܂Ր{]��
p ^�ZS�;�sp�88�����w	���|�Z�&��E��c� ޏ*��>��W��� ���`�$��s)������r
�p.���e�CG�O=�>�� ��Φۀ1!<��~օI�����l�q���?8�/��&!�^�C��*w\+��LTd(3p�����X�F�6�~�����T��~����9��� ��]���u��I���V��
�A��"Z6Sl��:S�����,�q���e�h����;�ډ��ۜ
�{������S�[?���hI 4%��Z�}9��?�O��`1D��Cqu�zq�a^ˈ�oĿ)ۮ�~��o��M+��Ro@ԑ	č�~���Q�$�1qW ��u��u����J|0冱�.��o�
�MNM�K+�W�A�lj���Z��P/lި�]���z��({�yz��il��4F:�/�A���D嘱p���z��G�����tY�r���
=�&[��sJ��i��q��������&,�lP���������M
�hW�����b�+m����@���d�n�/�����2{���f _�)�`��s��W��ޡ�)}��}O9S�B�P.�����HB�\vM��[v�N�'c��ce�Ÿ�L�z����D�(�?�{c�����)�!5R���V�Of�mM7Zʖq�Kں�"@֔�d>�Y.n�±������,P`��ē���: C0�f��f"���;|�K�q��mG��Ϫ���.�O��;���}k�$�Ai��z�:�[�P���;�g0�/B�5��:�%��*|��a_,��)?�8����މ�G�6`�\��e\3��A�Q��S�J��VOq��{_/�ս��)җ7]�z��#Ò��Ms���6P�/�۷\����X����mMݧ�a�<��k��ɠ3�2�_'�N���)����2��WHBy���+��TS�c*q
�̾qD	�K\�l�U+��1Sբ7��&0�xZ!.C���U@�������mB�x���ǅb������`<�wDV�+���1vi�k�?mQ³�<�a��r���]`d.^���T�d���o`�Xa.v���H�un/��>]'@��>�Z�d�2�e}t���ew���,Ώz�`� �N$	�⨓�ٛK��?���&���gG���.+*�L���0��5,��t�4�!�Dʅ
���Cˠ��8�ךOOR: ����A�Ỻ:�*��B�������Vu���������Χ�.�S� ��b:>B�Xt ��Zu��6�`�lk	�N���SW�d�I��~I�5fNlٱ5	OD���t_����W��,���yc�,�5��<��Wx$^�u���s��g\+�HH���:�|U��[�3��]�ń��.�(�J���R�!��ԇV6�?��K�z��+��A��@�J1�}@]�{�W2q��ѱn����c��B��9�}�Nߕ&���$���V焑����"�3�iHʚA�`[+����)
"U���	F�m��ћ6؝�+Nb_u��ۭ��#������܄Z�|+�L��O��ĂA�G.���C�욌Hط�KHzU;�_;ҋ�b��X����zeՂ��=��s�{�=0#���0�oȪ,0(o��8���\���!yi�:'�/�r!�MaO�3��i4��'j�N%���� ̍`������&�75�,1Sk��3�],}|��7N�����A"�i�mh���(�B���w��Kf�O��ܼ��I���� ����h�~B�n�ړc:r��7���&�z�\q�׮Q��M�Ʉ�bv�b=E�����?W-L��r���-ن��WB��J(rF"y���]j"HF�z%�0����	m:k�4���=h�� rD`7.{�{䴘�b�o�O�ϋ	���X=M/Z �2�a��o����\$��KY1����O�U��^D��4��$P��y�a�\;��OՂ-��]��+�Bx�1	�4������*x>�s�a�(��+=��(#�m��vv�I3���p3�({~�ɣJXu�����������Sc��Je����;��eN�>��wh���G��&���m(준�C��3�;�N���	y_��x��g1B���y+����üTW܍g����!��EYĦ���C�谔~�껇�<FZ���߈�9�����,e�%(�@���D�Mh U
}*e|�Xj�!��*7Ju�b2����Ѵ����K�k�\��vG!zTi�|��8�u�s�9�B���A$��SP -�x�˩AX��pR 3�������L�nd:=���ŨQ���(b�h��c?�n0>��-K�k�Q��|x߹{y8/�Z�}�	��"��o^��&5 ��{�W���L�i��	�Cd�V).�T�u/���$O�=�l��7�����Rm��S�zyO��p��@�&��07���G��;c��ƺ�
�%�Z�$ܴ��|�E¾Y�7K)��o:�!���up����-�ƽ�5Q��x@F�#�,ߣ��<n#��=z�#��T�	��;VC�:�w�]�ķ�Q��%��d1��!���C{������/U�#ꏧ���NG�q�Z���]�Q;�R�oL���iW��0�O�]�ڦ�U��O�yF$���Gv�ŅU@�	�'
4�%UU�qBa�Le�	�4��U����o`Oaou��[�2E��)c%#W��Y0��q�I��J�B�����2_��x��1�� S�t8��릞�V=���f�OA�5?j�;��q��ף� Ԛ���H_�z���v�:�dv<�6 ��+�9z]��
,�H#
��`��=-��ws�ed�vR�zƳd)0_"�eI{�a�ɽ=�
�� ��!��������s���IM�Կ�*<��I��td��
얒Z���w`B�)�Ͼ��D-��),5���̛���"'�6�Pz��r+�ò0��cc��,;s_~�Ω�!�2G{%��^Xi��-��}~f`�������
7\s�i�
G�D}e*�&Tv�χ^�����I(�o�b�|=i��b�&Hx�x����]�Fj67�X�>�;�p��P#��+��y�#�ӠP]B(�����	#}�z=|)����Y���o�ur�A�!�L�T������t��蕡C�}1�a}E�]��ߟ� ���h.�9dX���8DVPz���YQ-n>��_��Ϭ
����+�s.�+���!��r�p��/���Qf��:�M�����쵄Ԥ9�[X�|���U��~2d��x	1���iA0�ݸUf?�.]����F�=т{T~�kv��A�ac>��g#ؙ��[@��"��-����Y֧ao����V�⤧(g�#�A7��su�����䗛k�Ik���M_1��Fxu��s��gXj�!S�,�Z�"�t��B��b��.h֝���6���L�j�Ha{�j��_�'��_oz�;2����J���Ϲ���L��ɇ��|diʸM��jK%��?h���^;��.1m���*k��ͽ�*��1 XhJ��=4��}��&G\N��0p��%Uel���3�	������8�\����E+�=��N��KW�MP��6g"%H�'��E��~��L�9��T�z˶P$al��'1<7�$
[� ;fV�������h��n��n.zXj'^
L��`�d�jp��$eՋ̽{\Kq�V �/�'�q��C1aY�:yC8�!��{-����D��R������V��h�`��U�����g�͇��rb |]��σAk�S���K����@y�2|&/�KK0F�C���a��e>�>'	R�HVu`|�)�O�3+�����3�"���n��$�	my�0��js��d��T�g\��~ՕT�li����E`63�T�0��E;����ھM����a�yKW%d��mK����i�>�15����[�����AE$�4�6f��FYNLm"�#��i_g��3�s�/'�nX+�g1��?�Y}���F�����#�`�lpBB6�m��R�nɔ�o����S_㝀nO�+��A��FE��l�f�rc�9�9�h]�ՍAT-�� �����\ ���l%V���q@�u;ﱐxߋ��^0}�JIGd��&���&�� #w�����i��(�u-����	J��{�4��ޗ}p���ֱM���^�e�̠���{�+�%7ȴ��b��V�`s�x3	��"�lh�]f�g��:<���c��%�5ѣ�BIIʯݢ�֨��W+b��R��eᰚ�*h-g���6�������"}��m8ܗ��d�l.#��47:��,T6W�g֍#�4��!ɋvi�ӻ����;�I��ʢbI7�Pq�B?�ZcuV:+z�t�������|K�j$+�B�h�j�c�<�6�������H�P{�ض�,03�G�A�1H"�o]�H0�R�=�tH���5��?��#u1��Cq�W��t���7���3b�|�5��
����N���_3�-�!1�����4�2u���L�U_J�?�呫�+��c��|fR��':�W�[�a������s�T�S6m�av�9�b��
F8N"�o�o4bb�
�L�N�l����.�|�W5��i
��u�x���6���<�1��D��K���ӮD�[�-��+Ĺ
�D�0��x��_N5�~�H�x�!�����S����!�$�a	��!�_��6���)���h�3�0KN\�I#�)�?�h�CC�'u��)�fT$��%�D�V1�l~ݔ�!���W��bCnYm��˕O�K;��B �H`�Ό3}�?��K.@̀G�ܥ� ��oy����:��Lr ��{<��s��TdY���5�2�]�x-!ר8 U�� ��ߔ��Z�������d+R�.X`9��ځ��8X�мk�2����̩]�q1�ק�0ɠ��.T���a�{~�f!�4w�fw2w��ʀh�Ҩ�]߾�@,�	�q�T�!�q۪�Ä �>>�UC�+%����=��D,헝Xn�9��eo^.�\���L�9;��szE����;�=1׆�gV�^�k�5-�i.�Y�
`��_3d���1T2���F�<-��/v%�Y�-��g��e�j)Y��2��9ݜ�8���>�=��Gl��b�H&�:��ڞ��H�%��_`7Zmq�?��!4f�|G���/��"�IbN�0-q� �-'�t{P��~�O 8��,m9H$k�?�zF�n���YT� �z�R���=0���a�3k�x�%֤��3�1��,k�!,�� y�n1��"����dj߹�^��S<Ԧv���
g-J=��o�~�|���	=ЧT̄`<�SM�K(����x�5�t�_���Q�&�;����
>���HH�HV��;���Z�":���SlJ��̅�?Tu������}f����0����	r(Z=v�F�/�qpĐEY� ���i�=8���e�>�ౝ��QG��@B4ބd��,ur���&�"Ne�H�Zgөq��L��lI˔6&��+�w"����&���B-,u�^�Yq�ЯQ�Zȣ�e��8ԡ_:�/3���a!+�z�ބ����1X���P� Œ�L���`�YN��=�/�%e�ٻ!���M|�曊�E�-��Եy����b`��;bqٳ?��b��Q�l��F���U���y�Bj1T�+?$z�����GWƱj�5��\��^H��2�l���ڶ�~VY[��(ږ���n~����_�γ��9�:k_Q���	���룐�����ڏ��3�(f%:Ӻ�o��'n��Լr&���ל9���x��X�~{���̲.�!d*Q�+��Z.��Ӹ���8.�=V\�J�y����Ƥ2_c�H]:r�te�!��"�]��K�27l�#��O)��(�x_��A�!k4D2��#�\����m�e�A�\���՝�#�m��q�ZM��9l7�n�>���]��8���i���܈�Z�>���lM��A�wVZ�����1N͈���x�~s��-�	�x�d��H��L���M{��.��v@��q�l5�(W�|��Ԙ�����=�OV����?0��K,$�p'}4��:���D�|���t����-O��ݺ�����'�r�-��a�u�lK�퉶@h�ۏi�7�#�%�8�]�L��۠����[�Wh&��dir� }����2�@K�p�[�{�4Kj�ɝJ:Csu�	�Q�%���;T��^H@���_n�������m�/u>Q>�N� 1�^�ڡ�B�P��~��L�����]o����L�.̭��ҕ �B��<Ņֹ��h,1z��ɺ��v��,>�n�f�+�O"�����Vb�iG�F�^K$�kN���Zک=�]�@���xX�}��c��j���j� �ֵ���
�2�N-�(�n�X���W��&i,Ɏ�1�
��VQ����o(�4=^���w�)Î�_���Q�%9�^~��ӌ�q:�3�`W�I�u�mLgDqQ�!U��ִ�B|oy�������"QQ��t�Br'��l!�'��m��[�)v`�>X����$�!I�?ձWڟ.���]�T���� |�C(ҹ=kT)߮�Ći�n����n��������N�������=ɒ�󽵫��I���A5�"�j�&?�9	Nē8��
V�2h:]`uO��L��>�T��w�aѴ�b��X��|sFtb�!�w������8A�EK�����F�qh��pB|Z�d[�J9�.�-Ӊh3R�j��zs�}ox�zM8��h���G}�k���y���j��Ǩk��������N\v�/�\�����3���uJ���쀗	��ސ��B�X�������	�B[JD��Mf�{�IL��
Ix��2P�:�O�W!EK�#Q��U�$H�ұ��m�{�m��z��j�S_�O(]��g����bᵁ�Z9��ZY��q�;�τ��L�&��,�͢qh�%L��~�I�n� �'���oA���&� >ԵU�P�m�+w`Yw��4o|�c?`qu�P��d����x_��>.E��vB#i1�3�S����Ԏl6���U�O�$A���!�%�[	��G�6�jr���LS 6@v �SO�y3���6�R�n@Ћqsl��c�c����/J���3,��.'F��z�5$���p��l7�,D�R�)(�ˑ�ʱ���k#����H�i����lb,��Һ�?�_��k��J�~�ſ���3zi����v& �g@ꏿk���.U0�#��{ҹ��# B�t��)�g�8��r;�`����"���)�&��F��8��wé��B-#�I�d�Z:�mu�ȿ`���#��!2�t�4�NmICN����zP��W����g�|M��n�j-e�y�~x�]��o��r���Ƥ��j����Z�$ttu �tb���N�c1������*Kk��J�.%��%��XuYQpty�u}��¢��|;�ʎ\�lr۸"v���  �������ӣ) ����7ڀ>@0�՚�P�d�����|�:J!���|o����VC@�.�W�G�W�F�5.���B���,���G�#�9�Z� �.�������_��wcz�&5��%qTi�����)1)ɺ�	4��ع{��⌞1_��.�hR�+��5S��LȍM�����'�C��^$��y|\�^�!(5Ek>)�D��W�`��� ����Feivj��(��LI���TPF��1�7׮�vH��?-�m�ö.�B��}�@�g���%��2&���T�u�Ky��o"�P}�yzt�<�ä��X�)�pIn�V-�6����s���#'�q�6��;�W��*7�X+�@p\�h�8���z5��H��]` (�_SS�m,���zV�;牃5�oH��m+f�s�]����=��X�VMkQ���k)�#��T	�yh�X���e�rS���j��X�W.��	��B�0��֩I�,j#��De�t�`	Ȟ$� ��t�����'2�rƂҡ�VgU�q/OzE�&3�p���@�>�_�;9��Wa��)�Ѳ���k�Y��)O(����j��I%m	?RI��:;)�K�a!h�84���g��w�Ժ��&_�eu��d�{� ��α�F����h3c��F$jx�w�O�0a<�m�E��5%k%�������'�v��pH;��Q�/�J*l�E�%"׼��3�z�j2$�X��x)�,P��Z�]�o��(��J������G�#o�[x?��h�ᯃ�g����3�r��fd�o��E��b�����BȔ�@��&um�4�F��ޕ �  sRM��/��u:hG@�t�D_�.��=��M�s84�1�̾=��F��I�s`餸0Fӿo�6��Q�Q�*{��(�1�"�����1���&��N�J�ΈR�K�Ga5,h(��]5%w1�M��V  �i��0� ĵ�W�j$}��r�ܔ�Ji��nF��lSv?�|��?�5o��9�e��u�5���fd_i��3P���7a%��V3��+`!�e�)��<#T�M^��5�B�X
 8uO�Z�q?� ��C��U��L���	ZܾM������y���|O�5�V0�H�0)]����B��.����◳�L:�u�x�ad���e܃�y�m;���Ŝb���K HJMJKܼr��a6�ia���@G=0�ڗ��s�ms`�N^�pԉ��{��rM:E���x�l�Fs^M8^��2�8A	y�*�������Vm'�� �������@"B�p�x��a�  ��I����Mwx'��9�]�\<`'�Ȑ"5%�r�����	�箉�¯G��+���۰z1������PZrG���s�)�]����o	���wB>uMR�ٹCDd��$��g��\h��֐�,��]g f+������(@��Q7ޛ��]�$��rݖ�Ltڼ�~7\�j��T�)��
o#�B�󦏕�({-Ӯ�2�'�h����z�����O�[%�f
�݃��>��]���ܷgn�Z&3�Sd�X|N�n��L���#V����[��HX�Vc�-H�(�~�؎^���+���/F%.	���'Pl�a/ϵ�rgɫ�� ((N��S�0b�J4�ME"�3DX`_:$��e"�-�t
��rܗ�iw++i��|G�i~ܮJ�:¦Ml^p�}]:v�N�9k�|�`ޝ��Yz��oM��,����!*��Yq���7s�o�a��j��s��TV;
�ON�[��N�)|��`1���ebP�ū�H��5�i�%�^{��Z0  ��@�X��4h��|;a�.��c?���8���_X����{�";�2U�hw�3�/M���������J�[v�p���D�!��P������`8>�D�ķ]%�/?5G��}�@}���2vR��.>�ʺH<����¿s0T�B`� [�l�xa͊	��$ �~3n�^�|��͏�T߁v��k�^8Y��� _=v%�x�Ǭ�Սl_p�V���C����uT5�!S��؉HM�
��gE��#,���l����2�"�	�����ln���KM��M��z^��|�FN�q����Y�Sζ�U������ta�-O����>�i�[�z!�]�Cm�[-��F��g�o�ʭ�����R��qg���!Lت�BX��v~~�RH\�s�!I��d��^��
{���	A�q^����}�(U&ǃi�U����"�8ǉ�n_"V��gVzfM0��A�Vx�s�T�JUJ�j�8nΉ�
 n��#aF�u��R�cΊ��~���I'a�.�� 5ڽ���?v��0�Q���ƙ����Q.�J���Y�]�|��JL��d��5��!MO�ζ��p��[���8�(�Z����~;��= [8��k	4���gCW�[߯����9�r�*�pbm�$���v
!��U诜�S_y�&��-�G�A~		��c �=@����|���q}�\5P����kf�PTb�����5'O����(`�L�$4h���Y�w>�M�6ÈR��]=�
�AJ>��(�5������?wF�J��/�;X�-�V⃌�p�I �<���Ɂ��j�Jq�����c5�����f���d�� ��<�P��E��2Ҕs6L��f/��<�)C=�kj���3,�}�.�4lTJf{��L�L*�_��h�k���8M<�ksn)Ck~�S�q�"+ɴ�ꁜ��T7��3������k�,䨳��5�xFR.�GU�����n��	1"��H#����h��.mi	�B"H7��}�y
7�a���݁(�8���Y�W�\G�tG�GI=���������Yq���z�>���(��G8|K�OplG���I��5~n�G���z�r^�ps�7�M���Cc�z���ٕ���y�WoZ�{���pq�s�L
)��Z1&Q0�G���:��h��[MjHyB����]���)��°ӷ��I�P�p�ct%*��x�N淜2^_Q��I�.s������~k��7c���88`q�tE��W�����]�����7�$C�K�C\�0����٤n�PČ?�N�����ٮ��A��;D��R^�@zQ肸5Y�e�}cl���Kw�֣����a����F)�l`R�$�q�t�����$�ϗ������i=��s�kHj��d=��R��o�b~�L�w��o?렷i������OX�*MO�~������E�1� 0��5(8p�QRM�|n'���$V)t��N�^��eQ��$�"\�3Rv���� 1t�G.{(ľ�<Kq� E�C/����F�}}i�o�\{#>rd�C���<@�8f�C9ph��՞y^�)����#(���G�;�V^)Y��GZ�5�����7ƙ �]�R\y�W�I�(��+�0���T�\�P0����g����-�r� �Ӱ���]�E(���	��2��3���B����3C�
�\���U���Ƞ4��|��
�}��=+Au�.�t&/��!JR��G焇��Z@�&����'c(�v�M��sp�ct�Q�+ܤ�T�xT��^I:;{c��#x�c�[�O#�d*$�Ю���
�BB���㽻f_*(ƍ���J4�q�k��PVDb# [*�/����f�}�B�8�K�t=/�^n���m����Q�0����ot�� �y]�j5�[kJ�m%���*�S��?G�+�<�?�ٕi�����ʨ����y��^�p��$�P���fK�N2^A��*�Q�V�W�>�Ũ`R�i�	�Y%!k�s����}��$�cl�x�W�����K^P��r�y6�xt{�qꡑ2>q��P6�Q�o�ĥNj�w�H ë�A�:�H#Ϟ�.���2ɹ���V�W[����~#�^5&[Z�kU�p �\�#A>K��YF�� ��aw�����&9����w�����m�k���m�	��BOix<cX�17Ϭǉ�	��5���O��x�"�o0Ըb�>ڃ;���=#U~�K�f���
�Q�<?�$�uXx�	-�������1��z�2.~���谫�6�+tu�&-�>eL����+mҤ�-�Ŵ95�mI�<�X�o{������I�P�2&x�g첃X�|^���v��#p3-�mr�h����y�<�w���f�\�s������;��
��aa�*1v��;����#�	��J}�<Rt=�tJ|3T	�(��k�3���5���_���0l��G>H��ւd���4{�g�����.�w_�kv.Y��Tؒ˗B���  )M,hd[�W�E�G�p;��og���4�i?�߬��C����$�bq�¡W���Qø| Y�������Uf%�%���fV���V�S�h5|ҡ�7��u��4� ��G�GS�/^��Hy^�XH����>)�e�)#�]>�8	��7��M�ٟ�t�l�۳H�/��*�,�,���[k���!���ǎF�l��Ds�����Y��&��- �����<dL�&��0j�)�V.�jk;#X|`e JX��Id����v0��@­�G�T�_�L��K���D�3�8��d��]�uW�S�7p!��F����x��Rcŏ�r�P��]y���gA:;����r��Y!MA7�-�h=�?u4�D��~�͂�\�:�I�I��"oQx��nN�d�{>S%��C���yc���#�����H�5/h[39��C	�B]EtY�5�n��ݕ�i1p�����}��]��v�~�2n��?n��4��0P<�Il��'r���w�^�n��`��/�H�/�-}�צqCF(�'G��|�* !u�)'V�q�3��n�b%��z��l�!�R��!_�F���M|��7�
��k��um�SF��U��#�<�C�58�s����6��#\60������`���0�4<������)�Z���odg��NЀj�X0����Vc��H1��a�:'/�X�Ѡz~�k
�^1c�e��e��_��7��)��;�����]�c�VhK��j�w�l�M\��4��]�h�R����q�3xy��5_$,��ɤQ��+�G�8k��(;��q��{O����;mz$-&�o۔��j(��\��MF�o��W������%�I?����.���7�)�;�	o�>�w�����ġ܆�X�|j):5�óxj���߄�8?�X��H�1�-%\�媋��L���0�F��<.r(v�Z���M�ø9�W����v� ��pu#�}���y����F�imfB:���n ����(�e�����cY1o%og�Σ��g+�#T���S:�3�w��vm�
R���-����7�Ӵ�3NIߍ�;���zIѼ&ƶ��^��&Jl��3�6�Ǎ$����B���+=:�*?р�J\BED��A�5�(�4�t�A>�;��띸`�%"�͛m˰��ߤ
����z�~�n���W\�L1A�YV��r�PBy��/�<Պ�^v�5d�3�F�Q�}����=�%ل�AI��|�j�3��PצЎ\T��t��9TVOX<*)���q�;�)�׷��MZf7�h��$�����r\�uEЊ<gD.����>nNÆ�<�)�h��h	����y���2�QW_L�p2U���	���S����Z����#m�ڵ��M����d}lc���Yy�M�J�\r'i��1���0�=9���)M���>��P		�2��$G��;��~
I1�,eC�������#'��[ܙ2�,<l�J[��ϟ_�;�������F���, HgXņ���(a�5��;���hL�� �[_������%��ѪX�A���RTH� $�U�|jJsd
��j��T���_��[���E5��늲�s��lFB�����H|��6^�NU	up���J�C�\獂7*��B�Sΰ���*2�0O���!��i���/:��l�.g�!�9ȵ,�Q)8��������d�������j�"w�����z�_6��a?�]�N�3I�`�W);�0��fhJ�~m�����Ƒ ^R|N'��z�� ��j��ŴN�yP��.��8:szJŵ�wj��£���X,�"�r�����%��Ŝv��H8�.�~�7��_;5p$Q5��S'�f�˨��n-�����gЏڠω>s��������6f�I{�.�LKhE،[ ����
_YyͲE���a���df ���y+�?�Yek}�ՙ_�]�-y�ȏoO��4���>ٷ�U/ݜ�Q��B�����^�S�*��0�i(�JD���ėGAK�ǬE��cr��~Ņ���3�}����C:��Mu�=O��Pu��}�q��6 �\ܫ��U��f��2���g�MO޳JO8h��4N� ���DN�F~�j�[c��~�� �i,b�`%��gd�S�Н/��~�����P/79(���B:m�y��p�Ֆ)� ؖڈ�j�������'+T�)	ڈ)���G��e��a��Y ͪn����L�۞˓}?����HD���C)S�&#N$��.^�'���K˺��I�$�L؎���C�
�N��Oz��v���ю�C�*:Ӳ�I��О7�|&�J��1j:ʟӤ� 
4��^�[d��1�A��X� :	�	]��@۾Wa��C�;�3���:`�8+�5/��Z�ɭ�vW��xW�BRK�D�'���O@%�1��d�V�o��G�[gg�I��&GR�<���>�ޖ3�P)�ݰl�ϛbV;��1z(ء�t*]K�p"A׍��e��hm�:�꧘��֛.HU}(�vmu�L����V��Cq��*��y� s��#f��{��CaY~�+��{����쁼�R��9�ϝn�8�o���A���*�).+: ����_}F,8� ���,,ZśD�\54��5a��s��Җi�8��W�Eϣ6!s�c���r�v,Pc�����O���p�5N��L�J�P�������lX�Ǥ`�%�5��Q.�	�v	RW׻�ř����Wb:��*O��7��~����fv��z��e�����>�ϱ��_[����i��@#�E7u/���,�O��R]8�A\�<!,�h.����y~ARZ�MC���\4��|K[��*a7@����&u�<�I1a�R����c+��ǲ�5�w1������or&۬=��
���U
�âSG7���j�0��Z%����/����-}*����xR�Kos&>[�� ~���=T/H��:�;���/wP1.�c��,�	��vO��ư�ڮg���:mF���J��<;+�0E������Z_pHQ�T�Њg�g喩K���ɖM����q~���2��uXs���Vg��Ҿ4�}j�m�\��������wvn���u����1�!b��h��N�<V.�GM8�P+�C�[�u41y���hq�h�M`�z�.�B��GEr%`T�瞢��2�U<#FF��V����i7B��Ha'?8�tF@��C�<`w�4�ǈ^G�Ȉ���b������b)�x��=q�c��T�����v�3,�)C��x�Fb��h���W����Oi�6\��Ii��MG���y_�^����y�J��lԄ�X��˺_���'�⸝)J�D	�A	�����hZ��w1)8yJ�)�����0_��e.��i�"S�AoL�����3<�_a������&#�T30$�9�}����{���~_ʽRR�U�c��"G�M�"�B�J0�)���\�u��P�5CX�~�웶6`�:m@�2�.1X(s��7�B����z����\lU&��FAٍHih+p;�4j�Hh�����z�D�E#JJ��k���N"���J��ч\^I1�~ڹ�r��N�fh6��I��ޚ��5�ԭ6��2�.f]������Y���g�`�������u(�@蜲������ݵ	� ax����T�gH����L�磌��V���<��8�"w��Y�Rm��!*;w��\,���X���74SY^�pY��yC�7yW>�C2Y�b��+}¢U{b���P4�Ѷ��+�9�����SZ�����09�#�"n#u�����)�A"����?���sEX������G"
¥������rw�O ���,��d��1~Cj��;E"'s�A}�zVn%����<���;����yn}cf��w|H���C�YP��T�����M�*��\�8f ��3�T_�
=RT@JR��Č����EV�!rW��]������Q]1�)u�1�t���g��ƕL!c۩XZ��֯ON���T
<�9ڢY��"p������/Et��/8n$8��S��#_�E�>���d��5�gF���F�b�nQ �5�]��_�ч�尢�TN�q�����z�LONt��n���w#�Ÿ3-�_XI:�ܱN�͊f������t��ϙ���`R̜�qף����	�S��Di����MGv`M'��}<��1p��-���f|�5�c�}��$�����l���#�8s�\����3���d棸��P�恳�Z��V���蠔zM�ĵ�g���
j>;��-\(6(dQ�BO���2�r{���V�������Õn�Ϻl�{���vm �6�æf�ci��юv&]�<��$ܮs�̯��0�	*�h�=ú�v���q2Ȥ,�=4��1X����h}4Bu[���������2���S�-������Luyz�N3��]���I8T�I�������
O�������IW>��-aI�}��B�{�^;b�g�'���5�L����ޱ% ��%2�)$��綋�-Ĺ��|c�`TO?	��f����k�L6��)�d���g&���i:��7�]�w��X���Q:2�
��{M��;y���������ٖT�e:��8��9r� EX\�4�+�����QkzH+q�68�z�:�g�e��U�֡���b�#��H��Sk
�/G_��T�+U�.H��.�2]fIw:rvTl:v�zK}�_�R�=�<Gvx�r���1w��\�iQ������0��<K�w���3�[[Ǻ��|mT1(yU�Eb$E&�Ձ�����)뜋7=�C.S���+�&�ff�O)��A�q;���=&�U-��YP^70P!��:�_~n���&/�,��K�2:��Zm~=T�=��FRs-����`��~p����u�Է8�\'!���[��:m����K_87�
7�0�g��oG tf9�#`;�
l�뻉��Q禙BB�>���9 Rb��(����){�(65'������'��;:U�3
#ZV��ء�tӇ�A�z(v�b� �eb���[�1�N��LG�8m��;���rNO�O�Z�d��2��qdH�e�wE�J�g�� �-+v�dX�`E�bN�QrEͰ�i�"�K[�4YH)���
=�M�QT��{$�����k��a~Qm��/�l�I�s>��B���pG,�fv��2�:g-��^������`�f�ɯ�-��_��0������;���@6-YQ�%��+IřCu���X��u�!x,*���5I�{VX���
�%e���:���ΓG�H���l�;/�i�G��H�R�B];	�ϦU3���Mf_X�je���{#�>�۱EX�7����HC������)}������9�(�@y�����_�?_���i��b��ĕ����x;_��!�K2>����SUس���h߃V�:�������x�[�Vg���b�0��[���h�cz螊O?�������H̹��틅� ��WK̝<��/Ey�Z��>ɲ�A�����j(�6��A���ZQmROu0��<-�E�m����
ÿA��W�w��r�k�L�_Д��n�,���r�1�����p�@���	$I2y�`װ��v8X��}篭�b?.^$fB�Տ[�]7��Ur�a��c
4N�r�&���2&�#X���n6,�0bMn�\s�8�\�^
��*`:c�B[���8��#D�S��Z�|m��d���=��0����>-$��oU�x�l�1������m֢w�wܘV�s;�k5~ٍ�X�N���,q}
�KG�v�����(7~�&)����D���u_�>UP��?YڥG�7M��>&�|IO9�i������6;>��ג3�]9m�؊��7��'�+�t~--#FB��*���C1u�X8�}J���I��v臎s�ug(��w����6�WS��@��Ş� ��Var+�}��T�ϲ�`즊Z�Q��1���8Ԯ�B�K`)�6�/`�����~��w��Zm���FXq@m&����)��̒%
���F������������5�����_�V����F ��c��̸��e�3�M�Yut��I>-����5I�JlBʡ�Eż��EJ𵾒|QmCL���}I~\�!\�|#~�>�y���j`�#���zR2��q#r�a�s����-����9�5��:hНΣ����[!���ފy��P[�F!7���uAÎ�79��\���M�����5���g�p�s}��U��*�ñ�Cy����8^{#��ϫ�i�&sT�$��+xߺQ/++�b�.��;"!Ka~{�O��!�_��b�Aڇ��&�m��xiӭIn����bb*N`Pks���`\��%�U��-*����]�(�c�Eca�=�)	#��or5�\p���(��G�������������G=�j��z13쑝I
�]��Z5�-F��u�����z.��K֖Fz��x�1���I�F�`|��Vpm䥨oz���L��?�W�A���i���ҷ����e�(�$�d��9U���(؆��_,�ˊm���
nǆC�:l`J����(x���Y���2�DT�7�p'�l�::q�7l?��-��Y,�<�"I��R�1A�{�>8�gV���Ou�Rt�Ǻl��@�		���<WI^��L��T�C��$1҈ �����ǭ{��<�Xo ���f>R�����W7�H;O&8=�f4O�9�W�%ďّ���.8�z��}41�칌��������n�L��dU�甓�Ǽ;P�>q��p�t�!^܋��h���Zxs!��������z
'СF�����Gy���0�w�3m�a�L��"~���x.c��eo�R6�S�cu�"��1Y�~��3i�$�������U�>�q���ې*#��\3F������7�#�^��J��	��8�b�d��P"֖/ޕ�>g7l]>���w���UՐ �({tf�k/pW���a:~-1�'��6>�����Z8��R]�UC�������&�xAkFu���$N�=�x#�qy �������T`n���m��
N�x;����< �!�.^q��R-y��s�Hy�d��g�殛Z���4��T6{cH g����9e%'9��{<H5�r������<K�.��|V8�S��^/	?�IIz��C3�,l��"�S;vUx��C������z�Fʛ�l������B��HO@K�����A��x15]�a��x[�ٯ�P�	֏z.
J9Z�}�R�$���7kI��o�>4d����ަG�M��湁���h�~��nMK����j�m�y��k��a�G�	`V�wȰ,*���i�s�1&O�ii*IN'z��ULrq[>�E����p��kC6 �P�z��}��;t�/}�qN�����F�݄���j���8����� yBp�j�yag�r��T�(���^�F|XB~rإ����^���9�멷�-��]�O
D��}��u/m�\���gG*"٪�#�7���F^;]��w{M�F���߷�.,k�p �_dw��B4����'9�h�����)�����h�D�/a�g�A���"`��x�9K����"�o��������{�ߎ0^�?=�B�� T<5�b��E��֍ H�k[�%�M��A8�}��4�_��PS3���4I��,~�h�v;퉍"TR��Y�����h�4�_�F)1&s��� �mH-��~�� o�9e�Mc8X���T'�Tw�ڤ��$z�7
(��B����7��	�@�K�a/�J>�	|2����-O�������	|�i���R�H
��b��8Tl���@��X[`�y�B:�V�y���Sj'mю�$�2_}C�@��t����,�jt�C��㽻���t��;뤄<S���	u�z��'�	�V��J��[z���;�p��l"�5��������~�[��b��c<�a'�\�2
����-=�9aH	U��{��_��L��T�SK��F���W�#k.aɞ�m�/�	�k�dy��@�S�d̍�BK|'z��`�?%�`L�r����Es�+�	&���}@xN���V�Lp0ۍ��A*���I�mO�v���j_kz�d�s;+�Rq��4Zw�3���%��De&��Lg�/9,a\VG�|N�����n�R� �k��T��*����f��Jc�<eIM�T�%3\Y�x(Bd����ɸ㌪�n*�޷�d.��;�NU��hH�&#�%Z�2?Np1K=q�L\&�ۂ�t�zG�Cd���x�5%��'��Ԫ04n'��}yG@�S�W�9��B]����!@2!����"t����9��C26�u�63(�ɳ�H0���H�#�m9��CI��x�A���J �ޞ���!��I%p�E�"6�Z�~6�Y�m�)9����Ġ�a�s84	4�=h?i�j���x�`���{I� ��r���)ci,8��@bF��L5,�����K%���`���/�&�õ=D�+4�//���9��`�-)Y�W��9��&V�П�g���P�~�a=�H*�
ҍ�7�i�=^H���EϢ�j�yK��Nqv�XZk�6CϚ���e�����P\��+��s����NNW�s�%�Aܞ��m��]�W-��In�$`�����OT�!��c
+�]�@-RP��Z�j�:B�6#����m��!)U=�k5�_Q��yt#���YKi0�`��M{�z�c�(�O����"�P�L��<���sZ{�n��k��S�Z	$�
+t�q�d��j�	�R!�������a+H	����_hm�-�� �I�>�)�Jq�aG�8M��e4�pP�2v��3�=���E]pҵ�)�����W������|G�D��9�����n�C'��Y�;�5�%(~Q]}t�Z�&kD��X%y-�1�!�G���[���o�5պ��@�|`�|aҋo?����AE��z�:�f��Ԡ:��m�j�b"(qnRu��9�^͐�r���W�tä,�Em�S��6��!�ͱi�y3����Y���'��Zk�3GG��׸�.��z���]���G4]Jwv�MR��Vmh��|��zd��Ӄ��%��̪U<��͐o�����@�M�M�C~�u�������o!|�Xl��r��w��sJ_%�鼌`e�M��9�G�9���?��@��Ǐn�[��轄��?j�k�
TO$����q�翅X�CA­v)[~������m���� ���J�v�pnLp������9���>�>0�n�E�FA#�F}ѥ�=�r��ز<�hz�+�q ���R�U3b�/��T�B�����^�#�kJ��%q�
���$M����w=���>v�\t��=���]���hl��5����Od�6hІ�{1�sE���?�k����e�ڊ<���\):��p>�eo�$�DЈZv����-�� P�j�Qwi�S=]�q6�td^рK�:�w�s4��9N�Qr�����Lt��a�,A4&��ʲ���mx�#Կ�i������B�X�ŕ�AO� !��cu��]��Z�K�H��^�){G�����+�S�l&�g5=�b�X@����,':R+~���:��E^.Ԥ�!Ǜ�Mr}BR� ����K�ֳ),)ݖ�]~%�v���C�q:pK�ÞW�{q�Ȭ����X����3�vn�D��(q����#	tJ�LnƂ��rέ�zw����	lLX`�4��c3�ESW�Rfyf���؉$��1	�e(ד6/%�\����.���?��N�W9����YO]��\�I��H�Ly�8DRfO���G����Ȣe�����ϒ.��1���y,��I�ࡺ�3ɼ-�'���� v���~:=5K����Q�����Π"�V��Ac&�}ެސ�	��3N�cqN� Bw�e���f|���!�P�
e��0�h,^����d��K~�G�n���-݁i�V+���A��mV�>���裯T��&v�B̅u����F��Q����y�朗\#WPL����/e�N�ό�;qsy�x)�̼iݣ��Vcý�
n�*w�}z^��Ĕ���lϰ!I��+'�g�B�����	�[
R��Ao��2_�������'�"�m����x1Y��8��_�*b��K�>���/j��̯K�Eu�(���a~)�7��1{�=���y�a+Eݠڳ�P,�xf�����F��1���:P]���ݖ�=�iȂ�U޵�ֺtQ�<��t �9�����^7M�}�*o֐������
pŇב:�\Fd�'d��Og���w˧����Db˺<·GŌ�33s�ﷱ̊>Ûj7�R	�L��"�~֧y�䢴o@ ~l[����Q��ʝY�A������ք��6�<��
nt�܎�X&�N2}f�Q���p�9��8:��bX8"�6p�
�1+|q/aCQ9%\}��!���m�;�|̨E��1�,�U��]�ʈ@`^��y�Ҭ-<��F��Cqb�8$|c_��3����vܻD��0Nz�Ru����u�?^F�A�15Zh��c}LcY9Kx��$ț4HN��t����  ���|�+#�J��-]����Jl��U��� 7����%�\�K\!G��0V�xl2����r(�2�;���;0K�<��x�5����btƂ��H�HIy��ٯ���Y��]���b�2ư�{uU|`JO��+�/���T��$���� �*�oEf���||9*P�L�g�[y��C��Ok*��Ϩ3�?$�z��@�X�R!���RJ�I�^�Q�Ӝڹ�E�E3�R�Um\�'��1���>՞&��J���u;J�ON�
�����t̞*�?�3-c�F��w�ª�g�4sh�o#U��h�F�=N67�Ρ��^��D�����M�Y쌑ym���Fs��b�&m�Kr�;D�L�+�dj��ީ<�Y�S����L�����'��Pl'`��~`��9�Q��_"�|��
[�7g�y�N��Gv.���o{bȺ��׃e�zD~:�����O��p� w�s�G���Q4n���8���0@�Z}��59D��(~�T K���[�e�0���G
�C�_�t�LL,�:q?�o�frA,v�9F�-)7@�w]{�s�"�I��X��i2Se��aV����i��@�˫	?Hr�J,+h3\����\\����-�S&�9��K�c�ow�(�o����/�A�gN�a��<P��p{VլB3��U��Ll8�n���)�e�%HQ^��]a.���	�oYn	n�8�\Ԯv
��	PN[�{E���E2��W1L��_22�2/2�x��a�aR;l	�ПxW۪�}R��w�i�������t0��K��q�n��zN�ᭇ=R�y��O�ŕ�Y��g �pSՂ��^�i��E͆װ"�r��'����``�3U��8�#�R���=���r{#hu��5�{D�t|r��3K��o���C�x���mcW�$v�QM]0���,#�b�%J�*?W()mg��sq`1�-RE�F���"��Yh�6W�I�)jk��������	Ю�U�kN�0�'y��BM�͍-�Lx|��[��<��BQ��=(+�+?�ft��.�3�G���|�{p���5��(ژ��¬���]q|���J\��k�>�����ͫ����(\��c�׾bv����Yd���⏒>.� ��,�]���G[�;~�k�=�9YS�7/�7�C� ����Cٗ�Y�a���+HW>�����E"\��	�
�A�~�Bz���N̭��0h*�2�3�RK\Ӆ���ڸ�'��J]�T'/�-y})�ܰ'2M;�ˋ>���Jj����J���L`n���<ܱ��S0�ç�PJp�E��)�`=1��Wݢf$�<��^�:�5���������e�
~7,%�k���B�ճ�f'ч�䭈1C����f �N�<��"w�T��s�yb�|��H�����[P��H�|��Iw#�@���ja�k^T�z��^4�)Wf�Ɗ�o���=��q�F�+����I׬�ҁ���>�N�`��苓������M�H�)2�]X�-�'��F(Z� �W�K�S���ImI=I�����Ln���PyZ��z�	�<MLS�D&�o�O��-7lb���M.q�m�x@���X��~N'+,��1�	��QK^c$�1�J!� ��@0�8����EV5&8X�,4��Ԝr���oE5�{�-;��"m[�^w���v�D�+���>�B�N7��ͥ>�,h�����M�p%�&�P6��7)��-ڙ;���t~;z��C�6�ʱ-�nd������;�]�D�ޤs�ق���"hi`�t#�S�A��
e�-C�\`!���6f�f�ӋXO�����@��1��f�zZl2��^Ns�<bm�=
" c��&���W�wCo��W���>��}԰�Z��x��-��D�g�8t#y��w�C�&��n�@���Em����G�T�wʌ�������l%�G�ש��]F�g����{lf��a�>2.�ª���d���MZ��/.p�悒[W��-d%�}����-d����1s"z�i�a��s��B8���%�@���ǖ�n�5;4e��ɉ��a���9�v|�%����j92ӥ���F_mFRK}�g%t�yb���g$�h��q��HF�t�;aI�(
��5@�� ��z;��-���⁷'@�x�Ѓ߽�&�?9�?0^������$���v����F�}o%A�̬t0����d
�N�����o �4�R�n�P��>�-ۨ�;L�Μ����~�f[E���#au�؜���X�(��Ԝ��Y�ћ��|�'*�D�� �g��LD��΀�v���%Y�g����~��C���/��m��h.��hbI������]�����`H������w��͂>���n[3�v�����.��u,li?O��9S/T}"c~�L<��pH�4�=�+�]��Tv5[�89�z����+ԃ�hk����/@��Z�T �>84����3"=�+���7����2���SC 
���6D8~
���|"��cY?��� +���7lꕠ�M�UZoO`���}�x�˃�?d���4_4��<K�D7���&\"*q?hR���mR���UQ�1��X��`��>U���;бZ^���f��b��6j�rl �I���W���m�O��z�GR\*�ҏ�a�e�XO'A��[�`@-�����d_\��cW:�8��m�|L
��޺����zz^	��:���� d��X���!_�9��Ɠb�����+���o�d���5�غ�̰���޴(����Ht*K֖��ri��]ok�� ��L�F���9Mi~��(�}�;1�[~�r�M�*��%h[��s����"��R6!��WGu���5Ƅ�K:hiWRwB��x\_ꊰkD�+x�E�Q�P·�ZW@�`}-I7F��}����0{�P�D�O�\16����c��ۆ��gĶ�Q�Mިm�g����#ރȬ+�uJ�]���
���u���`Y�U�����e6M�}�g����5�j��T^"·�b/�bOAS��路#u���������^bj���~�ݴ�Nu�o�W�A����:���y��jߨ�\�R���-M�9�z�{)�!������îi
@0̳\��DR5C���� d�q�'3�sb"�{/��<�Tj�'0�tF#ʝ!�Y�w�f#|��yPA�e���#_f����a����(jʯ�I��mZ�5�e֑�m��r>g���dQ����mb`�4�ޚ��1e"֥�>���ݨ��_�F�p�Q��T����C�uCV��2[s�!�Mt�V��;�iK���e����`$A#�^J�<���p!d�ZwjWy��G�� �I�F�}�{��cT�!�h�{�cV���H9R���A� U�o�+��T�KY��̃���C����� i�YBEe�� g7~�ŤSp{�J�}ƨ�rv�M��d��|��CE���(ԴJ~�/�K�'�I�z�p��Z�b�Ł�;l`���S����!��W����!�$��ݪ�Й�
1������<g��z;��}�6qKB��p}y6�E}'iW�M:xʩL�e��S2��-ۙ;�wG
�ؓ��u,���xgJ�-�^�Gv<��\�(�H�G�����C �hP�<� ؓ��&�e�3�bҺ�e�ۆ�n'&v�:�4�b�<�� ���.��x2F�tW�߃��u�nα�þ�T����q�������[��3��jY�Y�N��G�B,MGA�]S0��5]v�Ue'��c2t�L�};R �M�ODg����,JE�]1ek%�]�슋}b0{-!�>ˡ�R;b��@����}+,�+�# 9���� �9�����;mf'���.�kmcq=Q��Ǽ���z;Oof�gWpr�ۗW��
������Ү���A�#�n[��qK�b�=�����+��w�(�b����ȉZ�S;#�2�����Ao��i�@
~w���3W7x��������2$e�')���ʂ|��B�+�['��6喚B8���u`ѱR%�3���_ X��u�ѷЅvY~6�X�V�c�)��Q/�{�����cB�{����FW2��|�R�ޞSENp^��Gҕ�i<� ��j��/�H��i@�&1F5�(���
���	13�Q.G�I����Es�K]�I��V��3���A�~5�����h��G.�����V3]3%��;*�z�;k�0�{!����I�fW�΢"_6�.����%�Ԑ^Q��;��ZbDY�X�j��������� �pF������6+�<��lG�7������&ǡ�����q��ix޽�rDˬ���F��/a���/(�H��u7Z�^�@�usx�Pwu��s���A�� ����ҧ1�`Q�g-���F��">�W3N^�&0<w
1<����N�-V���r����!1�r�M�� �ν[��Rh��4@/FF�54���E�:f�7��r9�Z�K"YF� ���]������h{vǸ���q`k��\s���٣���cy�|N"R�ن��.8�hFJ�����Q�u:�mM܋=Nh�+D��t�{W��d@��I����ɟ�Ms����ػ6�f+~���5����2s.���ce�� �LY���m��N�B�2��R��4��|�����X_@{����� ����I
�72�ۥm��S�_�ܚlQ"�(<���,�Ox�n��}<���T�G��1J:q���hf�TI�_'�N�5>$��;qT�5�uȋ��A���Aq�XGЀ�FQ��x���_���Qd��rW��g�m�BFiYw�KG���n��\a{��O�i����!� 
ĳ��s�8p�����dq> h�C7�s"��|^�_�s)�a�Na��}l���S��<N6�p ��⒐\14�z��&����|�hph��p[=y���P	�Ŷ�� �ъ�V�^�A��&�Y�&�#����Q< X�7Y�	�qN�ȗ�g������wUr��Km���i�J�H�
����8�ndk�^����<%������i�^)ń�u�k�Q�mx~؃MG՘�W�8�J�V(��^q��xЪ����gd��G<Q���/_�����-2t�e ;�V���	�	�cbl���#�R��U�5}�Rqj���
&����(E�/�ĩ�d�_+їj���:d�tU$Pq[3|�����U�T���K��uc��,?y��u���BY��bҞ��Bv�X�Q�D쾌�����iS�e�÷-�=�f��{MY���ח�k�����f���K&��f����	�sMXq���R��sι'$�tl�dRU�R��R2��N�SgB�:��G%(�uw;�렋Q��B���ˢ/TQpJ/��g{~��p���E��e碣4���Ks5#�]I��_�N3�'3C��>~藺��v�_����h����^��R��",������zt�U�!&� e����P*d�;y�v����*[�����ʗ��ݸ�kfїs]�T�������K�Ǒi�\�Rg�j���a���@Ĳg��6�48�M[��8�Y ~1���vR��+m�$m�΃�S�(���!��|��ZC1���=kX�Ev��ֳ��SN�#�lu�f���Q���:����ѳ����|��P�$�'.�g�X�� ���eoR&}�ӎ���F�6;�}ȏ�~i�p���hPؔ��蝒Hi�mx��F���Q9�yUdN+@b&�+K�Ju�S���D/�^�D3&���y�3{9�T��D��d��K>PC,��^GI�h��6ԑ� ��Ҙ����m.tn�ﵸ�V��*�A���3a���B���c)��	���9%��\`b\��N��Za��\&�"^ƻܜw�_z6�[�b{NBmZe;�	���aө�O{��:,{��p�}�++����?.�G�����9Iy���zQSXOVw�םM��(H�YYGjj���j��X�"_�[�r�^1��k7���0O'�������B�e��~�5�ϔ)��5=�y�+7��۵�`�c��pl��;_���o.��E��� �*([; �9�~lfͯ���µLB�����|���$iv9��?u��K��׎����lK�g���N4��=t�GCt3��1m	u��j�2D�-�(�r�B?�|�]��*걮�4�N�C�J1�O��&�vJ=�^�(�`��Z `��D�$x�f�E,B�y3�p�A����S{]o�ԑ�p��X-K�)�.��4���)s�}��@~��[����������=G�^ӄQ~��@�+0����s���m��x��_���X��h`7��|�>�o!r*������lq���O��M�fw��T[^��G%��L.f����UD���Ѧ�#`�m��"�gI���e�vA��� =R/�
���Ψñ.���s��J�9KX+���x������т��%/TP������I��*���5C͞�(dxt���A�)��7��"�,������g��$E�ey7[��є��GE�X,�yk�CyqԾ�̢c�֚�Sv�L��oF�N!\Df��D歭��+b��j<�w�W!W�a�a��=}��h�%u�?'��Eу>Zj�uw��o�aH���2NnS�Y�7�9pfk�	&x��^`�� ۝Cӷ��Э��L,��>������~X��y�d*Z@i#���@W���<�齣��e̔�G�6-���%�~w��i#]Ԕ?�Yv.*N(?Dn�M]��v��r�4<�@��/LI����W#�=������$X�� ��F�f��i��]	V��y�8�D��U�o�v[�xP���JI�I�qkӀ�_�HΏ)�	���������B�{�Dwև;��q�G'gN'�4kP���S�����S�.��X�Lm+��c�i����݅B�,�m46K�݃��}��X0��0������=���5��,ocSM�}�I��Ų� R�s�0)qp�?�՛C���h�-R�4ߜ�6G	�}�	�5˃U
f��V�l�$g�����:%���A�>Pձϳ����ve�y�D�q��:��37��t�N#6�hj��`'>��t��l���P߻�7�!mάD��m�����;���)s�Z�,���e��%0�`���S���E#{Y���N����\g�A�|�A���nְNF�z	I"�qq���G#R.Sxm�r��A����9�aI�F�Y_9pO��d���d�%�e@���ss�~;��,�p�Y��@�R���S�����.ky�x9Y�2h��31Bف��}����_7&\e!��6�IP�n�'��4�& �gjM�o��C>�߹d���P��`����;-@ӷ׸04�1��I@q�c3������w�`??�X�?��e3��@�nWD��$�uT+�;I{���q�!��������������+v�֔���m0?N$|�Wo"p�0�	�'g8:���Ƃ�[G�p��L���A�S8��F8�[��v�Q�{�L�u���c,�Rm��R%��c��]KH�.��D�>���if�;!���?��M���x�´yg�z�h%/���U�+��9_1WH���&h��`� ��,�:�����ʗ���N$Ҽp���"$��.c��wf@Onz&�[��}��֒XU Y����@[�	Q���@���)%U��2��q�4�@��� -s��#\�����NMY�VN�~�5��� m^>�F���(�:uI�L� ���g1IeUd}����N�U�t�٦!ܳ���S�L��]�p��B���R��?|��Oj�e@��(��a��*(��y��*t���H�3Ii�e>����p��:��[mI-�f�g��n��������t��g�ʠV�����l�`�esx�Yq�s�{��wt�y��{o�WK<�nU<�e@�ڲeȶ��.!�웖։j*H-���6+[^&U�}y����uu& ���[�S�4:�Z:UE�۵l@��Ma�#N�n�a}�%�j�/��]�$V�z9�ݶ��iS�Ɖ�^�~ɋ^`�d�ύڇ�������� D$���,y��ԏ��2�A���JQ��.4���d������F�H,Bj�u�?qs�p�oG�G��p(nE�g����-�,�+���P�{ٕ�f�K���z�����	��KK܀�x����cFE��0M>H{�&xÀ���؆�� �g�K��9�Vn�o2A�N"6��q�5��տ�a��g��S�ﾸě7F`a{�j�u|Td^e!���|J���Ki`�YC����y��Y|�� �K��JYqX�W� �d���̓m��G
	I�A�Γ�+u
.��._����̩H�Q$KH;m�� ��RK��l�E���5$�r�w�V� Dh��b?=�0I���T����`0Ԙ�����R(��3�����K���a�h8̠)V� M	�Z�5��f��� #yE��m�h�]��H��&�}cr�M�[����L 3�9#�[��z]t�Bl-Q\h-Nbr��*��]Z�O���֝>���Yj�]z� �/gɯ��B��������|����1��3���Z!��`m��0\���RKk�W�����n�飺��<�d�]Z����)F�ol�cS�4ρf��T���>��~����VpO�G~��/V˚���]Acg��(r��~��}�������S�@n�6+U���Zk���\�;�ӕ����Q�T�������M\�/��\�
[�=��rs1�T>-?���v��ǅ����G���O�G�K�q��z|p����u�H"�ڈfB�,�ΟofR�(x[�1Ώm�"������?�	N��*!g���E�j��7�Qk��1?����N�q�%�eu�Y����As�RDi���"Jƣ;Y�;��9W��Z���X��ހ��킝x ��R���g���ܬ�餸ߔ����/	�6����j�ݔ��m�:��3�h=s�����ff��\�m��Ѓn6��/�l��p~D�%t���y�M��b -��kU���7¸4�Q����X�M�04{2¤�3��ļ]޵s;��3W��<��?�"$��X�uCe��B0�������zC�^��5c�r�0�f	�l���n��q�^�M4q�1$��ﮜ��!�&��׭˦l�8���𐊅K���A��)��ϓ{��xm�'#�6K��i�Ł���kN}�+�ʞ٬s�'��xܬ��`��]�=FO9������������2�Pb��P�S�=����>.�����F��3`�=�(���6ڌ��QZ%k�ģ�zF���?-[���&��I^��j�Ђ�y7d>�ZrZʖ�Q5">�Z�֫@\�~���HT5(Z5G~����2]}��>Qn��eV>�M�F��X�&T{da!�3Mp��%�.�G=>n��O�|��d\*X�Hޘ��O~�}���c���IEM�
�ۚ�M?k���$�������'ӍҶ�a�\Z�����G�~,%cM��FT���@,�+v�q��b�5�whxΘLR�%Z�]�Mh*ʀ9���Z3�i�-�
+R�t�g���s ���������w���o=��*$@C3@�e�S��Q�����>�#\�J!���Q_$ޜ'<�F� ��/ro&L� A��V�3���ȱ�Vv��Q9uq
yl�Vf�P�����i�F�K<,�v�`s�{q�dc��'v�����{����	K�W��Q��b�?�逬V.	_�d�:ܹ�O׶�N�r�(�Pw8@%!A�-��5����f�K�+��ZJ"H�����5��v�t8���W��G]r�G�ş�����j�9��Z}�Q�>�ƈJ�f�E��'=L0\޿t{�'a��}$t7m@���=���.0{�XB/a�������S'j���}�W�߫�9"�M����c$�U �wH���(�E["YȳbP��@È¤�C�%��G��Kl��_����J��rL�BL�.�	�N��i�o�P�$�	��Y�s�ڥ���ɑq��W�mF򆒝9{/����(���kƀ�]PV�B�[��TA�>�}_��H��$Ld�r�&�	 D����\�Q��~�NH���C�!'�������ОP�`5j.�	��f�wڱ_���!/�7�ZB��b��'a��h�f�_T���N`?��i�Uڴͫ�����5��z2'�[��I���#�V��J[0�ćȿu�}z�\�y�v7C��)�S ��a����4Xء�fxl���+3��rzh����dq-7���8y�J��i�/��ȋY(�X�w���j���sd�Cm�B!K�o5�Jy[r �c+���� #.��?kBg��jJa����7󚺧�U)�5�%G?�?hf�<+��?�K��ܛ46%��eA͑b.J���B�1v��}���q�}�t�4D�ҭ��6��ǋ.]�{�Y�~�e�;n���<f���V5�t���e�U�w83�Թ3ɹ��s�C����eю�Hj�ٕ�?r����Coo���zJ���������Y�ن��=�sQ�9�N�q�ީ�A!N�B6�yo)�"t@Y{r�}S�8� �t^L����!㊚�_&���H�`�5�q_p�T,x
�H�(��:7-�`ˑ��pR��180��a`Υ	�X��bq@M0޴�K��%�Ҧ��q&��Bx`]���X����A$��K�t���/���/��ٗIQ�q�3�x��o�=�E6��w��0oo| ���0��fn)��Q.������vRs:;P��j��EА6��2�aeS�3�T\�[*���(������
*�֮2ݬ�Q��󺂏��j>����qXZJԠF�G��\Ի�Џl��N��3>�F�����r��)cb��	�%e��/�s;x@�T$���:,DRLmu���,�%��}`�J䶶>_�����������(/#��p��kWE�e<��k������N$�P�C���3���r�hr��i/<�w�i�i�W�DȐ+.Ƌ��[	xėᒪ��8eU�?�J���@X�v0f�n^ �w�>�Klg7`��R�7g7{���M�^y7�@�?p�H\��ј=w��o�h��Hu�tH�*<�bY�fc�H�]]|M�e�ݢwr4I�+h��l��!���w����c�;����a��?�19-���ؿ�� 	��	a�`�!L�av�Ǌ���)ġQsz"��&Ikb�L���7�S�s���,ߚ�onJ���K U=��/���JS�"���G+���"h�m���M���2|�Xy�֌k� (���´��G�<Y	8V}�YK3I�?��{��ӭ�����3���Q!S����k�.˸pz^�u𤘦�3:�)fl�yth��K~����Y=c�cb�H�`��E�ݑ}��Mg�[9�sv˛�2��*���]�"�}ycˠѐ��n�_HW�������D@��[�R���H�E��$ѥ	�R�p��jtkM������3n��x7�F�Ֆ?���I
&���^
��ڨZ��".�
���:��&u��l��(Py�\y�Œ�9�8�	x)Vhv�J�><Ok~vi�Boسˀ�)��.mu���$2u�[A�R�f��	�Ln�iSM-P s�Jz�H�F�F/�nɟ�X�83(�{AE���N7hY�IJ���C<RL4�d���ޕb6����M��MU�(c���A���+�y������q�����W��߆t��Ѽ/�n�R�>5���N��v�7�n# ��t��[�G'k�1
u��ĵ��I�7���<�&%k��!��������dՌ)��1����n�u�����ݯ�˸��b%	m�m�R���܍����`EQ��=/&&�S��e�Ɣ�d_�Yi��ʁC��͛�#0��S?j�/�w]���ڦ��D����
E�!_����vF��E�>���-���wI���aP�������M�׽�U(�*�毴���^ZېĕP��(�<M�n#�."���.Vf$�X�V���Р�6��/���S��9���r-R����D�G��$��?��w�B�V+��iF��kUU��gP�r�3�`�s\��K�����oG��,�k�̬�W։B�-�+D�t^�zk�<[ܭ��� z���c
���g	C~Jp�c��X���zJSO�����q��;��n>ڜNA�HG�Y�Z���c�e1b�m���W&���%:�U�A*����3��߹��f����*݉z��7󧒺�T�x���0��ԼZ�?���H����Z�Fp�^A=J�7ᨑbخR_7:��+�/?`3Tͨ��[u4T��0�ow�����X�a[_k���ΰ�Ō��e/,�,G�O�-�A"�8o	���
9�E�dsE���6�Bt(l���%7�������p9�.

+X���W��lr  k� �⯏[E+h��9��� 3�8Ș:m��MYV6�&9���L��%��X7��loO��Ea�T���>�����p�^�Q{@�v��������A�����Ì/ϏB�*� ��t"D%�v�w|);uY�L�$	���^�ѡ>1��;�����H�L�n��[�����H\��E*D�����^S7;ғZ�wjcAX�������ٷ���>}�5|�b7W�A��k_3�:��Eqde��í�1�7���51-<�ے4��-fCO"�.��֛���Xo�t�%|��1� 9�Ҏ��e�Y  �/nC��A�m�X���~t��~A�4ܸ��T?i܇�-�ɅE<�QIf$a�P{�o9r��a	��	6�9+Z�H���G�W��7w��n� bG������w�8O`"�i�H���I{t�5�Oo��a����l�D����\9�5e�#�=]i�K�t��VYh@�(O(hRw�xo�3��6���XW('ҵ@qU��Da�I	�j'E����x�
��'p��e{y�S�A��^�i���ݾ�b���8������ʕM�I�������-�0֦��η';��b�sDǧg}�s����=��{M@S��V��_b[��S1\3
���:86��h��I�S�8���|�e�t�o(m4�·����vV���}Ȩm�G ����yۄ4u�(����7���;�� E:>�!0�Čz��+�"��H߂EG%7+�GY6�� 1�r6K���Ƨ��.|�(ʀA�^�9ѝ
	����L-b�����NP7<��������F �{�&��o~bY��s�l�N��4x8KOGȼ���k�+��2�G��JM�F��LD]����W�Kl���/���5 Fw�X�812�+Ï���oL��h�F�%@�(�摢;Ux���*�W��F�sw��5�#&@T�V̬'����R����J�����.8�ZOᲂ	Bk)�ԡW��R	�F���9�.F�?�� W<Q�b�bǲ��]֫���j�ZsN�������S[j+��ǳ	��R��!F��/�cs��/h��'�ɺ�JS��JZ���w�*�X���Dl�M�lu�� ��㽌���
�I}Yˁ;���b��d<�|�CXB1�R�Î�@���z5����9&��O-�a$�<_� �����=�\U��*����8d��˾Sz�˽*)uӦ3o�):�?���q�
���n@�~������)v5tw�N��8F�-��6B NΗ:�­��TG)�>��?w�k4�^�P��m�&�T1 z����|�f`s��W��殧� U
N��-e�(�h������ɮ#�Bq��	�5习K���tV��jϽZ��Ӂp�Y1�@&�
��������6�ύ`����+����t}jޚ�R�$fMŰ���]���>|L��:���[LЯC�~���og�b�� �05F�<kb+���������5��sx�TM��O�~#5:]CU�I���8噼����Ή��`-xS���3f��S�<[�
Œص�Rc�h� t����b��A�^�z��i;z&m�� �0_mI��Z�@o�>C���:lS�4}G�z����d'��*i��_����Z �V���ջU���z���N,�s|2�ӌ�F����Q�y�q_O�����`�� ,����w#5܀��HXK���f��[o�3��^0a��FE<�]��Pj#�'1x���m�y���ޱI�o�kW���lLp���_!��F��{�_����#�o�D� �R
�#�������i� �����$�D�ե����[����yRS;Y�C����{"dLE94`���0���L�XkB4��� -Nތ��&j=&���<�"�7��(�W�~˹q��{�7BW;x�����m2����3�Mi���X��PXK|�GL�Di�K�U�SZ���J�,ǋ��y�@H�L�g�0�?�h�	��s{�/�m�4,�ywW}A�Tz$a_A�rN����6h�`0��{क़��0$���k���.M��f��O�IO��������0�bv��}�W���i)�?o�5QJ|m[By����{������3�\g}8w��\���Q�����s(��I�qtCA��:��5�-��c�D ��Muٽ�~�b%ʾLF����(����h������x��X�+E1wft*��ow/c���`*o>�l��E�y��!aWݷ09�7�H�f(����.-�4G���*v��;���|TQ({��^Q���{Q�ڀ���3��_�<��we�Ѷ,�\�����R1Ʀ�Y�c��w�n������k�D)϶�\���jՀ(`��86=_�	�k2F����$-��s)n-���܆lw�0�7�Jf*'��K"<u|���t!�e|,-�|jʻ懀`�K�v��$`�缍���&Z3�a�Ӷ��P�Y��$>���[�������6u��S��W��\�K���D��V,r۽�}���B^S�l��!��mlR�h
ej�����0�`JMvE[pEV�����A�P�'J�ެ��/����>�AF}�W�U�8�j��J"�:�"�#�e��h� %��5`��< �vϰ��V��i�>[�Y\i�1$Ch����j`������o7#�
�@a�\�O�0B>�JRK:â
P� [LP�2Id_+o�fD�`�+��<���a�:�v�����(8�N�F~	�1}<*��l�1�Ɠ���Gڒ=�����Wt���.)]��J�jՖt���\�RŞz��
��\�Vߛߡ�'uQ��#������A�W@U_�*�.!�-H�l�d��w?7��w`����U;��]p/��*�^f�Ԁ�N_�p��L{�y�R���y�@�s~B� ��<�3Á��07u#���r�R�C`h�a����{~��Uȇ�������WҦ���[\��s��������5�^
��$��ȡ�i��ї� W��Z٦�W3��5g�dr!��.j�hӪ[���} �U�[�2�ȸ-?f�E_�@��� �W��K.�&�Z���CX�^
@�:����'��M�3�F�U�;��|�ѽ��L�A�nѡ�����!w�t��)?�4:r8n�g�nϹ"fV�B��עIѰ�a
L.�
�\T!4�8ۗ���[J�B@}�� �B7�ޑ������֖�#����}C-��ĥ��������n�81 �w$�/�v2bؑ�^���0���}�,��J��Lo.�4�C��R!] ���#��{��ƫ��� @H�	�7%���Q� H���lM.�ˇ�tW���NwI����LX�Kn�ٜ�x��Y�/S��pZ1�=mB|e!X�*2���k(
�]�Z��2�ۤc	�E��nP��g��Vp��J�0"2 ��Jٲ���ٵd����t�����(�����OM^C��`ݾ��;=���yV�H�F�n�d�=�PLfB|�ɍh���*:uY�'+ȱ�~�p�����(>����BB2�#=�]:}�~�Qs�u�	���<�	����%d�\H�7���n7e�R� �F��W�u��P*�y�O��Af�rؙ����ԥ�RN!z�+���7�ZMᤠwC�^Ц�I�'�b�x����%W̧=�-��<� .�Q��λ=��-����o.�@:�OƩK��7d�=��\r���#�Lҽu���~#�\i��V�}ͽB��V�?��v;����4��$�}b؁ņ��O]��Z2P��/r(pj�����=F�p��<��ʚg�d��N`T��/P���N�ZR�m�,�k���>7�Y�J<:#��mxq��`�#�e�)]��g�����-�e�/��Ǡ3���z�]�u��i��衠�|M�������p��p�%�` `�*D���N���bE2H�;zh)�,3/YQ�O���Q(}�U��9��Ҽ�
��%:��r��VވPr/�F�,z�����V�Β�=u"��!�p���-䯡�_ϲ^?����a:�º��f�촳�q�]R�HUj7K��]E4�}�{�8J�4=A����8�t\'}�i(Fe;%C�H�Y[UK��uo��B���`���%w����)Aw��T�#I�B�%�Lᖩ��uT��7檬S�@����1�g��|��	�$�A�� B)f��G ��Ɋ����-{H\IM�[�K/'���vȊ$�Eu�4܀�H�r��O:B�MO$�����"r�}� v�Fn��9��^�8�O[�ٌh^�����C\� ufӾj]�(������20��mw���KҲ�Ks�U=4<BeW��x��n�7P�5�Ž��5��e1�z�8�?-p/�&�ʕiq��$a蘬���~I*����X*�>�$a�O�<BN�z���Re��ʰ��N R	�킚-����S�*>�q(`^����sL�~j:�J9ݛ2�����%�>�_ޮ� 0�a˥E��<������t�s�� �C^��R��\fhz`O=���YY�.&�jr���J[�3���>�/u���&q��QN<$��c|�AM��$���2����w]�q���c�o�xI���c�#�ސ�>fH��S�N���t�xJ�M���,��f��#�B�W���z�gz����	S$�����Q�J�н�Ju8�?>�������;�Z��qC�m�IO����*���������ҡ��{(4�s���sW󺈍�~5s���f�ߣ�x���U����7%�����0|�Q
f�k;�#􏤪ۍ�Rr���xu�!�w��ps��
�cV��0�̅Ӓ_��ɴ��Mj��~E�vUI���J�����/�C+��O�u�������Ն��'1���w�2����ڀ�]��j[���'��p���}����>�b,a���w�k�f䙻)�$���UO �gL������of/�Q�Z$�w4A�}�l��yI)�&G�+��E�{���.:����k�"�F��]�����a��\"=���VܰݧQ�6�6	�+���CY!�Ӝ΁���h�t�.���'ئD��+��0c��M�9[�0��(�0���C�l�2E�S��ʿvD���D ��+Tl�Np�Ou�-N��벳�x��Oaȿ�����}u���U��zV��X��b%�vn�-�����r���Н� �52 ����q/�loIj�oWvo|�U}��$�7�@�1���i���l��*��&�Ȳ�d>��uA�o�GD������5+7g����S� �����R��~�3Xo���,k�����VlZ߿E�o	��&Գ9�	�n�b�G���dMb)��pM}f��9�I(L�V�2Tv�S��,<&�L.��aEOs���&��K=Uq�������ۡȊ�t�\�i^���1M�d�O������p"$qV�B3�W ��<N��o]徐��8R�����PK�0�M��&Iّ�*����U}Z��Z�B��@��3�$�|O�*l�]O�&�� ��[9�����|x�u��nW@�=V�ȝ�_�fA.��I4�8�j��K�0Y��������h
v�@[��};(� �����)����w0�K_:@1�.D���Y�B���, ����Av0w�#C>�\#4�g���ϫ��y�N��#a ��"�8��Ã/
���D�� ��:��Le0Z��"���9UEn��68ng�wH$�	����?�#Ճ��0X��*�ud�8�`�_=����]pJ�����R��lG ���5�%O���p��<(�]�K.��7�@���
%dX.�(�mOwF�fi�uB��� �����moٗT���ў���fn:L7~P�T'k=̈f�ɤ���fR���W
nsǪ�o���am����;�hʠ�m�w�H#n0J+��'sd����~��:�[{�����O�c6'��rn�Kh�aA՘�N�)��^y��WV�Z�N��-�S]�h@;��� �V
6_���Wu��2Y|o�d{)*�tWۑ8�S��%�m'^6��/�� ��w�ܴ��x��>��۬+g����ҿ
�^Lݪ������hO|��=�k��U��J�`�����0р����*��/*��� ��N;"�r�d}8�\�m$��-���0�f���� �`JyVN�l<����{�����s�wD�&e��Cq�Q<�9��;\r��$�M
�JRy|t�ա�y���/����lG���[����Ȼ����H��Q��;f�[��(��U�,c��5W�\�{"J�=��X������C���v�GZ~�8��S8y�:㩢�~�$��w�����}��l��7�n�1�� �T�/�A�Gt	�͒�q�����.z�������u;�e�e��!�ֈ�,:�4�m��\w�蛗�N?8<�YZ���R?�[�\�{�V��U��:��٤C���cҹDt�Jvi��B�R�u��Si9
�'0��ļY�������(Zn>��ƴgA�񔼛�("�`�� �rpU6lp���a/�J�J�o�uǖ"�����3���Ɗ�8hWٳM�$�T#NN-�a�.��|�5��L`�0�y��S	�L:��A�n?��^P���z�`[L�7u����>�	��N*&�d�F9h�[6m��f���_�`rwJEK�;�7aD���B~ǚNVt��[Lk����ȧsZ���6g�`f�Ur�'V�����a�
-�%4�#G�'�򻬓��|@$6$�3��DQI�S��Q��'\�e�D����a�Ǳ$�e?����	���݊�}��=@�s9����`�$`޹�]�S=���/�%v:u���@�ؔ[q���S����NN��}C�5���b%�����pԻ@cǯ:�~yŘbtE�|�+-qqrǢ�	�U�eu<�7ۍ��up1ȣq��/:��� ��\'���;��s��!N�K�x�e0�l|��M=��A��,�����'�q���vV��9����A�5� sS�d���Dy�x��Љ�_:���l�:"�&�`j$���9�Y0E?�;���ɓ&Hz����̖���{�7�|<���Ƚnn�d���}�j��X PsI�-�6�1�9��|]�'Z�ԶWɣk���̡��'e��6$.��]���K�����a!���� �_�kR}_!�P����Q��Y�BVǾ�������r�����tWJG��	s�Y����* }ҵ&��-\2o����� c�����x��Of-Q�`���>��:����f��한6� [���e0E��v��J�um�BS�p��
]�էy<�}O���1<B� ,c[T��n_&'�@`��>4�*��̽g�	��?�y��u� j�\�طiҾ�aG���9ӝ^�X�?(  �ez�r���q98��R��-��c�|��}�^�M6�U�5�Y������4+I��{-��֪�8.�e
��#�E�vf�l�ϻ���u)���J����F�j�l�pҖ܊�D��������*]۶43�k*�kVh�B�˭`�j����,F���G��nV�(D�2�S�ԝ&u�X�A08h;/O3�����t˚Z
n3?�����;���ֹ�,����lȖ�P���pE�����!^� (bԵ@U��I���}�����_	>n�M*��`n�6��p�zx����d���Ob��ʵ�Q�D��;K�J���q��
�җ�8��e|5�[�4(�x(.qi�vV�g'�1�?Цc���^ܯ$:�� (�]�C㣠U��k�GZr'�L��v���W7r���_�L�"�23)��xY�^�l�^#�u�Pա�za�[�
Wi���J�?��Ķۡ&�aY�'8�Dj	U�����R!?��r��^��>�tS}�[@��N��9S���ӣ��Mm�Ek�\��>>�l>�	�;���n]��ԣb�e�l-~�Hi��_�x[!��]I�oA�/�/:c�^�����[<ї9�p�ܵ��e����cJ��+�o�� C���
w���58�+G��I���֓�/�6��t��@D�;v!]���4Bc��@�I��I�uPЙk�ŗ@���h�:���p��S9֎�
uM*m��&ԇV�cC�h/z��~��d�;��ᾜ��N	�eU`S�H���xz
�*����F4�h��GP>.��xg^����*��v\~�����m6��
�7�*�aƥ�� d ���d>֐ս��B]�a{l��3^�ײ,�G�k��5�fY� ��lt��&�ΏE�����������q��,r�
~�\��\�T灢�Z������c��Z��w�y��7�R	x+��]!��j�*NZ�}o�nȽ��Q�}�;!�Dt�_;��,�ר�����E�HIn��,G��2`�>m���\žZT�H �/�1D����H��H�d���9)�$)�:����{��*o���1���0�74D�g��t/�B;�>��y5g/���[2��k�;��j��_15{��7��ܒ�Tg���*M�3k+@/!�����_��_(`
��d�O��!F5������Y�i��(:���T����Qx�U�%�!#����>���/m+;��G�dÑ@�/�Xn�'�*�n�{E�6ik�?����(���U�����q����eo���m6C~
��%k��5wCn�x��M̵G�/x ַj������ ��Ӧ���z���/h��Z���J1�T�����T9���/>l����߽�ZG'J�N��p��6��X�
+l2&d��w��K G���A�\��n�8���}���u_���4nZ���� ߵۯ�l��Ҿ xd�I��ҫu$��V}djfy}a��������|��"�iY/�"��38����)����F���y-�Y�*�c�3�l�[q��iR������;kc��E⨸y^���,�d0yL^�e����ZK�V2�^oȩ[��`W�P(��WM#I�$yR��@���u_$2nY�*$�A8�k]-��?�aE��](��)�2yp����J�-�c��Gβ��V�	��r���#�j�QtZ`L�T2��I�ES٩n]�z�^�� �P�io�K�3/Tgշ�Fҽ�E�~J�Ge���c��ݫ��5:��F�X�L[uk8�ֱ7�S�)|����v�ҁʩ_�e6��N6�������4g��3���)'��%�9��Z�Dkf��@��U@Cs�f���RB�� K}E��rvۄ#�:���b�5�<������W~B��45����-��i�=S)�۬����e��P����O�&�e���PJ ��ح椐�z����,ؒ���7Ɓd���/Ag��e�kJY��5��dV%��M��E�~y��,�ҋ�9��ݮc�-�SAX�&G��hA�;��9G���9�%'ɇݐG�R�/�fJ6h�9���X�#�`[^������ ��8�� z�� (�K���q��mg��0��KOJs� �u>�m�ɂ���8@?�F���Ʊ9m�;�1pt�êe#���N`���U��Ed�����i�>��x.B��-5�k:u)'4= ș��~�q�D% f��)��߯��[~��l5	���3ufaE���5�<#�Wy��+�$Q �(X&eޖ�}ƭ�~}�KJ�1����ekN�G�i`Qp��l�����m�d��O��|i�w��uY漄d}.�]��5 �0:����}��������yU�Ň��s�Ԙ�0� �����l��U��QS���Ѹ�eXͱ��g������R��G��.K���b�衻�D[ו�!�9��dH6iﰂ����/����΢m�����* <���V(-yz���X�����y	�l�P+���Lx��b��S�L��$�L���ka�nD�0��	�w�^� �P#|�֑�/���÷�2jۻHYLSG����s}��!ISQ����̓T:ᛚ��!��I��-���F�3�+��5�:53���g�Pq�//P����J���y��"�-�T��Wīy$�U]���+�?E#5�yc�L�\t�:!�q�F����>�Cu��W�0�~�i�@ \F��i�K�Pɔ�G/��R��8����L��+�c�G��o�2��㰷@�}(�H�x����F@�R��>�^Ծ�48,gG����lC���K�:��T,�7*&�"Ƞw���ikO
�G8��>��s1��L���^�"�$�Z�|r��С��M��3�hI1�U�=��\T�Tm����{��8��;�?x�}�q��*}Ku�Oi�\�%��1s#�k���j��_��Yr���<7���A�����o���,�rƈ�:w��f��tz���>uiYq�*��fσ���U>I���s+������0�Р���l��a54GO�<-H��Ht�ͼ2P #(�Rt�
A�j/~!#�R/��d��7(�\�#�B�FK�8t�W� �U��驊�x�/t\�&,bW�DF����],,��	�"���D�n�Y!��!>�<K��>�z/c�L�@'����"�p$f��F�y�e r��{�s���
PO�K �	mR�PN�#bA��NX(�Aۻ���2�U�9q {J�?��1���veׂZ�~P�RM��U������-��r��~����A;b����0�F*�Z���S�Nx�)
�1i��$���=�>_��YZ�Mf��
ڿ]�a�Վ�;ږ�uvY¨��_Nm!���CR'����Q�����L*@��y}�������	���'ީ������
��X�����8Y��`�Y�(�r�����o��!�bɢ���/�
ά�Ƶ�Ve�y�Kl#���I�}ˋ'|$t�b�fc9����A��K-�s��J��,9��H�~� ��n���h�?��J�g.Ӯvf�MV���y�nw|ץ�42)"8�^�,r�=y15n����Mi�)"L��D�!Vi��̠Z��~�>{�%��z"e/j�fb�Ζ�c�J1,G1c�~<��4n<m��ҡ��1���t5%�/�i=Db��)�~��#hZȌt	E����u�j�'��o��{�(�]eA�#ű�EWv�)0�`GB?-a�>�03_;���\����0�c$pr��%�49��6�j~sn���|\�]�]?�i�.�2#n�)���v��dH�6Ѿ���"�zP��\�%�-��`1�tk�S�Ց���_���2��s��LU^
� �Ѵ{7�e�����Yxd�/6QPԳ�v��%���*'�,�4r�KjĤr��n+�,ɻm�:h��NNW��X�2����P��2e���OO��P��+�2���P΍=$��"��V>�8��z3�z��E�d��+I��5��ޮ_Fb�������Bh �:X����V{*��γl���ָ�h���秞5�X��
UY���M�aK���Oц]��.�{��I1��\!#���W��U�R�� �����Q�[rawf���Ɛ!��{�g�i�p��.�!w���ػ���=-�G|���=�o��<,aa�_d�CΥ����Q,�攜jF�q�meP����:��G?�����A�g27$#��J�I3]�Z|�EV��*�'4��$(t��
�BY20��M��]���z�w�yܮ��W��Yt�u5�?��%�u��f�Y?Pr!�k���wA#7��FI�C�`\��Xg�%�+юGT�W�NF��Mz������w$�ˑf|�4�#�i�4�"Y�o>h�ٸ�h�@��z=���L{Ę��L�*eW����$k<z�_I��d�$9�P�������mC��{�arWCS99,��{db����P>���  9�o�|��M����.$/��p�ޕ������ϕ�v"[X4'�!
�n�]���0p�I���H�r*����(��Ћ�ޏ
z�D��c��"Q�q/h�ɫ5�;%U��`X<O�*��6Q�u�&ܜ�@oY�߈��o�2���;�����r�~g����ʎU0%���)���qi�k"~N��Z[�R�aϵ��Fq��ݢ�\z4J�A9��_�!�6#�ʔ~=ʒ�u��J9�9\<L�Mbl_Q�B��`qG���z������*Q�·᠎�&�(F��p>l9�z��l�Z'��I5�t�������`���y��K,��ZP2v
�b���@�PH_�d�𴬘.9`��Ջ��[���g�+L�2��W���c/�q��[�EN�~Yj���3���,�6k���z� x���'�����/:�Z��~v�QaJAN�}^��j�����
Pg3��f�s�c�����N��znV//ސ�m9�o���t�ZP)1ԍ`���{�ꞧpD �#aW¤AԱGt�K��Kܫ���<�*�9��MJG�b5�5��M�Ux���8���rE]]�p�3�:��ջ}�R"b��f4����v.֪7�jP��@�2V�M۞���uC���f�DV%���&_f�EV�ɣsQ��=A�E�S3O;<�5�hieS�T����_������3�h�q��C���-�%��Bߒ��Q$��y����USW)��S�*�2�)7�%������� D�\r[0&p�o0"���^n��4W����ľ7y��(�>��j(�V�TS;0�8$QY� ޚr�`��'�V������=����
;��$�ԧ,�`3��N���g^F��&m��*��s)/�
!gB�?��=`� ��BÓ_0�B�I<s�Y9 �n�1I|_�%a+�p���E��|P?HZ�8���\�T��û!��׽��NR�81gԔB�kxy�[L�[�w�Q	���k��jPƇ'־���$TH�Ǖ�����f���ߦ�����|�3wJ# ,n
�Rm@?�~��+)�ٚS'y2����ʊgP	��g�r�ߥXa-�fQS����y����n׸!-,�Kܪ��a�˒�=�tx"B�(���8����0�tY��U9�J/�`�=j7T���[����zJ���U��O+�vA�S)��h0�'�s�b����O�a��\�#�o��]'��m1��5gH	�m��EJR,������$�h�L���7Bޑ��82���++�0+}�;}߃tu�|�b2ń��^f����)�v�r'?so���5��B�� L�e/M���`��K����/����e�ɶA=���j\��W����%��5X_p�XO�Q򏬞
���'0��p��g��ec�|�'#�]�G��z'S4;��^N;�*\IǷ>��`���<~��Ar���m��3J�p�)�C=A���|b�ӻ��驾�58 ����:G��;���Y�쀘��V� ��!
�siwR-q|V%p�Ƃz9�h���7�*f����ƈ*�z�'&\�<�X��׌�/��BK�d��ǰ�ח�G��~T=�1�V��tU�]P���.|�d��b����kL�Ay�x]���H�L ����pg��m��[,b��6��[��i���'��S�5�Vx,��]p�&�<M�?�%s$wL{����������"����*�rm�H.L�{RKы!Z]N���8_�w��������J�z��~����y��vK$��&uR�u��A`���PT��֟׌
���*��d`	�XԆn;~Vq�EF�1���P*(VJ��I1��t�ĮSD��,9��_y��,�1 �?����>os��O�t�Hk��((��;��y�0ȡ.��?�w��{Ϳ���C���tP�ݣ���:����i���/�����W3"nW�q_I�~ߪ�;����Y�bx����^���e@S���[˄�����D��P��
O7]�u��2��Y`�Q6�!����3�ٿ���V��'^�< eG��I�>	�j�VV���h����ҍ���I!L���1&c����Fp;Y��f��
%��Y�A^���\���H�f�CP���n�lra�{X�.�_ny��1x��5����yh�%�̈́����􃸢��m��=�[��3����;v��3��Ѹ��#���Q�w����ҝp��T��f�Cs��RԆ�*�熲@Y[ª>��s<Hx@�G�Q��W�iC��Le7�����(���*m�1��ө��͘+�	W���TU�Ț'h��"���K�-}e�|�.;����
 _9��v���*zm`PU!���T��[챊���v�:K�ɘ�V�i��*����b�'F�4�ڔ���z��ҋP̋`k��R���g�����������㡢�6	�ֹ'��s%��*��kK�9�"y5�t�vGi.נ<�l�AE��_D̼W���P���&@w��'8�Y��8Ne�
�K��Zk�4u,�P��y��JU8׬�p�V.�U��ҙo�{�Y�Tr���9����*;�]wtsw�>��c��-���# )�Z�}�Ú�ڱ���Z?QJӀ O�d��mH���sZoB�=Z��̆��x��� o\m��%�7w��_��3dA��B��C��8�����ͤ�Ҏ���J�ΞY/�!gt�����}�b�s�Տ�%1cE�^	h%H���ah��X[E>ZE����"3?�[㞚Q��fkڢ+������4�ex���;��p�/Pk� ��x�EN��|�kݚ�!5cw&���È�����+���iq����_=е	E�~6��&K{lN�C��H7�'���E�vq�C���_��Æ�!���_���e�lN�$�K����z�@���UZ��K��)�8o��`5�����\����u��tp�
���9��,L=�%��@CP�WT���fL#.m5�y�(�_��5��,��܀�ڧ�ƥ�4���#�s%��0%Q��H	�^q�%"�g�"��["9J�W�!�Ȓx�D7(WW��}��8�@MB�!OBx�jKqPv꯿�11�%G��mF�����%{o�i��e���L�QЁ��x�d}/���F-j�x-D׍V=���Z78Q����b`	�S��ЦnH�!��n�h�8Io����<Wz��I��,��z��������B�jpہ"��fӎ�/t�0�$:̠��$w<�W9i>pe�{9��Ȳ��*�9��|�}Z�7�޹���0}LB�]r;�:�=�Wո��\�g�y����A�q����,��c����'Zپ����(c�<t�F�������L��̴��o���eƜ����Z�n�K�C����xn��L�n���S�C\��\���R�2vF<��WJJ�O�f�9��i5'��{��$�-X�m��2 �	�l��9�(5��h��k����`�*�n�-A�α~-�� ��[N��D��r���h�?#�'s7������ύ|�U�v$3@n�.��0_/���� ���%�W��#�"jU@9�ʓ#u�`�rV~��d�Ĭ�؝�.���_�Up<ȫAOsZU^�;�d#a�H���/��yj�&#��zf��7xݮt���;�x)�U�̨�U�fY�`��*�x�we�))�����o5�q��W��|�Uji���L�o�-Ł����&)���kDϟ�:ٶ�������6��:�m��~�&�+�	�B�}��L��lJLmT ���ɜ�2w]G��|�0���t���/�(_��O�1*�����F�c`U�սnc���j�q�� 6�'�����ɤ-�Cjoٝ�~�^0^@���؀ z����r|��O6X{��Wp�Õ��){;RI�6�x4R���*�/����	gwdѴ�Np$2����yQ$��$K���p��`S�kh˸�8ܘ��]�������D���2��#-��6y=�������͏pj�N�sV��W~�W�`�[��Ѩ�K�eA�"s�b(Gg�jh..�)κ��[�:䭖��E���^"������LNo�w܅����hB�D*Wb�f�O�޵b,$tZ�}M�Y?��uB� ل��LL.�@V7�MB���2;S��ۆ��>[�Zвp����؜�o���EhZ �&��[�����Va����S���~�4W�y
��nDRqAp;>rM����{ �<�.���]]5&UK�dB�k�b��Y�T��"�]��S��!�bB���(�B���p6�/°u^ڜ����!W�G��������mC�^���,���_�3���Ǚj_�(d�s��M'0@���Z��N��u�O�Wh(�U�FU��vK��A�Y�ty8�J��J���(�7|�	���~���e*�[R\C�~;6�C^��#��Ē�XɁi`3F�~C1E2�����kbˤ�o��;]�OY�G'ڸ�Z�AKz��	~+�c�kE[���EH��_4 �|	�Z�m��Y�2�x-�M���6B�_R�5�C;k�5�#mļ��į�������h�@H0���[�\i�uX��q��ll"���[�y	��~��O�n19�삣~S��%58��d��ʥ��U3��F�
vǭ�9�<��m�-��Sߧ�i7#�9�h	��z�m���u��0���&�Y��h[ivml�S��t*��F�+�@}~��Kf�˦�X��Y�9����1ڎ��/B��Y�O��'3��s}��T�Έ�U��|�}"�w�U�[L��� 
����A45J~Aa��N��Y�7��:(���+�4�+y	��"�[.�#t�\H�\la!;T�y��A�B,Ӳ�\hb)���GM�xi-����)�:�����([�ǋ�X���v�d1sUK�4�����	�f��:d�?t3�My�I��m\!f�b��@�.P�^
@� rť�׶s�r�c�/JE�^�]�Z�8�~0���7�)��v�3��`5-�?�r,�K<&���q�;�>(U@������m��KQ�S��t"��ܧ�qJ�o��z��|%m�݋K�Ԏ8E�/�,(��3���a{��J�b-@ X��܅����(��p:rZ��I�����%�+�Q���/-�*�����^��J/	BC��f<�|X4���F�����]��B\|~~?q,��~��}F�xoO`��	*XT4��/9P;�Mp�y�B�����VN�	��L��?0W��B��!��Ȇ�M2W}u�R9O`��䶴�ű|3�����)��\�o�A_d�u��ﴟw�,\�B��UF����"��(.5�6Wo�O-����;�зx_ǥ�|&lmVe�_z��k}[.k���&f�VaF��Wo�w���U�q���r,~`�r������/����N��eٝ=���R��Q�Ry="�o$֪���nj��'��ql6�RB��Oݛ��% _�ef��b�}s��Q�Z����Xm���#����Ke�5ol#�+b�iRV'C��Z� ��ā�|-_p���(#+�4b��<8v�(���d�D}gú'e�B�N[����W��M�>Z�X F�����o��,-�����$=����q>p�*�Sp��v$&O�ڵ2:����3k*�6g�R;�oO��#>����K4!ƶQ>��o`�h+$����&����na�T���8F���*d��"a� ���oY������ZE��	W�m���q�ɚ�Z`&�������D�%d�Rߛ��ެq���-F����@o[��2�s6�N�����O�62�������m#w�2$̂S�	��Љ���`W�r������5<���*�ki��*�5��_�yT��gǗ�sh=�"�D��_����T.ϭ��'��u��~�S�=��w/��t]\,O�-���E��o/��2莨ǝ%�k9'z���y�&��=��F�ۂ�ly;A��eᴦ�&ry���0u�)�_�,��f��iqU���I�Y���ڭT ������n<E[-�Zy]�3=@3���d3�:E��_ŝ�UO6k�&<�U
[|��F	��p6�8�#)=MS!H�������]���Н乽7g �k�GGH]����.Q9J'� @�j���J����r��]	ml���d�O���)2��%�4_��FKy�#�p�$����2�I�jH���bt����3CF�C�n�� w�'�nB�^O���6~}��%2�H�q�"ٿ��L&kmk8�^��ry�$҅$���=(��(�]��>�?���ؗ(J�S(_�s__j���_=*��e�%�-��b$����}�`;9��?��E��X�K5C���s�� �����	�!����0]�����W))��n����6�T�	g(�3��:5t�0��� QR���'Os���tv�Ib]��V��
����cG1�uB��P���� �H<(�6)q� �T���=�#�5�zDEa�X�����-����=�!�_c�l$'	��au�O����w�قֽ}�wk�zW�����E�gA칽�	�Ĉ.p��6�J��t�/X������j�	��5�K�=b=߽��0ET4���w�PmeK�Ʈt[*h���p8q�*0�`]CDf�cP#���&�3V�и���Z��u&�T��x�(�;�f�o�1h9O	cC��0������u�C��:I�4�Z֒&5��Wؐ������`�V#گ�����B����kPPo�.uk��$Ԁ4�m�h�!b�ӭiԄ=H6g!���1|���+F�shY#R�����l�KW.t�y�M�P� �̺X|39�lz�5����X����`oh������!|��w=<[��$��B ��REqG~wǺ����Gñ��:d��Uat4�ּ�����iy��W�0����|1�Q�	�� 6��N'����;0���v{)A��̺��Q���5�m(�>i�>]���u��WC�)p�ܳ�TB,�o�-�>�X/��n-����Z=�+f��-��0-��C���q�N��*��׸b�>��w1�c*� ��tDjK\w�3�i��	��. 0���k��È�x�Ģ���t�GRXq���&L\	 g������u��ZR?:��Md��p��.dǄh�����r��X�^l�H������)�8�NjGo�l�B2]W���\zl\Y�܇�xd�����8�e)e�6#�T�f��&3���t�}ǈͽ�I��#����o��Fr���sJ����<�[2��(..s6����ji�NW)��Y�<�Z�u�j��LEB�؁��1��c���[n�#��ă�&��H�B�T(�2�>Do���o��'��D��4�Yq��Щ�u�n<��N�rp����7��ͳ8��ׄ�S6tw��-o�Y��k֨~�}~'�9�
���B�d٩l��V���^|���M�S]��./��H�k�'��è^�Xg�=�ʷ	/Hl����]6����<��9)����9&7�*��~��Q#��>� �PgXG|wnb�.!��t�?��hs�UIΕ4��&��P_�I/�F�]= p��D�WnL7�U�&�絳Z�i�	>���<�Z渫�ܤ1;ve`	�Id�J���y3�g��c�n�8���&^�Rk�U"C85�A��^T�Q�>8���z" 	�t5�9��3tEu;M���xC�bʏ&X`�(HUC<�!���ޤ��S�jn/b��K}�_�]�Q��).�hv$z�c.	��^�+㠌�z��i�O�QQ�g�_�@SkY����ʑ\Vb^�1��ggV�o��+'&ip���}�G��[����p�5`�D�ܟF������1�-.<{g�+�?�mx�UՎ��`�>,̮L	�E��B��0���J�f[t7ZN_]�x�YR|;�>�I��F���`=�?�CJ�k���ff�qE�bC�cJ�4�:çdRwm���Vby�Tȋ+�@
T��t�nԺ����v�yA�󜷋e "�F)��aL������	�SX�!�2�`ъ���m�B�3k>D��I��0+($@<F��ov��S�s�v��`�q)�J�}`���/8���{�8�؇B��ye�T��b$��=PuζLy//l}b3� x�G/Iu�[j�/̭��sȷ֟K�Ś��!Q.w�������B$1f�Ig���F�:bY�|
.�ZG'���]S	z�z��`� 5ڶ�cK>K����(eC��zv�Fz���nL~l!ȋ� z�3�y���&�߬`�¾z�D�D<S�˥�g� �w��A��'�X )0��L���SQj���Ѯ�ʤ,�i@�50�&ݥ�ZeR..����f���+]E; A��7:bլ
��������sw�B�L�u(��ir9B=_�����j�y�\z��i�Xt�7NK������Up�9hr~�e�Ƽ���+Nkzc=Q�20X�f���(���L�6�I��H� jLeB6�M�zAu����3}BD���f%�	�d�%N�4��v�3%�-]A��_��KX<��H=4�%�~#��#SV�UT�/�I�'�	��b*2�j�NM��nc���݂�۽9o�Dm�� ���a�?E����n����R#�~��l?4i��pC#�����yaf�MT���P.1=�r�#L��p��1JG�x@{�KU��dB1��y�{܄���R�ļN�Ps��  -��ʚWO���3T[L���v�c@N�b�̕�ͨb&��a ��6����1�r]�@y�ma܍J�C-��J
�;�anv�b��]|ذ����F�������I$�d�RKwa��=��S��D�Gnh�i�����ME�M��g��v5�6�E&@�7��y>�I�Ԡ���?�H�ϔ��CpX�����:�����$4�M����aP�i%B�xˋg�EAQ|2�m���S�h.������so\{����2�	=5vB��TP��m����X$���Z̼���,����7p$��
&T��@�'�@�XD/V�{�^���:�������X` �<�@W[�D˓���
U�N�4+Z [-���	���d�K����k����]Q�mS\��h�m:�ǽ�\x-���3�X����[���
!�J��=�ꙇO(< 7[��� Z���V��$��c�����A��]��_S�`l��^9�<�%i@O�E�tB���䌷1��)vi�÷�+�p�����&4'�Mv1��t��ਖ���y�wL���v�p��%�14[�&���.4�7��7�¼L4��<v�+�"������)xL{��Ȏ����F,�(C��Je��x}�`3WČ)r�l:rۙ�yغ�X�^�,��'I��ޯ�f�����yk��8cX�/���.�1z
"�߭��{C�O:*�FN���ӞÿS�!e��9�"!�&�9�K��e�Y���OĖ��F%AI����h>S���jD��c9�(���>
�_^�����|�oH��EI=��C�֘�/��^�9��b�����O�o��ȓ_g$\B�U�����*�myx��Z�z&6(��wn���G��!��5Ѕ�u_��m}��܎����HG�<< r�Ơ�����wV�*�`��Ӻ����X.�4���Ϡ '6bx�D�XFs�|ǖ+��9-\͓]p���\$y��A�\�Hd8�����nV)��b�E��6��,�ӿ�t�13i�F��&ƽ1��*[����0�n�v�4���e!h�U��s�ݳkv.�ⱊ��?�8�������w�/��b�M#��A�]"�Թ�x�+/��l=�#t@����>"wg+���`�u��I�1�3�\I�Ŧb���-
ݥ���A�M��-d���ge ������9"�H:�U�Ln`ko�Yͣz0ʹL��%۞�L��!4D�����3͢�q�%3��o�	g�s��\?%ہ��lY��+���n$�ʰ�2B.�L#}P�"��&���T��|ҡ5mOr|H��	��@������Z��@I����"ZE&��˱�k���,a�	C��oޗ��ꧡ�r��y�r�,�.��lge�t��k�ފq-��C�:b�	E+�U�<�Hb��S�\��S�}!���MC���	0SZ$YQJ#���A�,��|���i ���A8��B���B���0�ĜvCN����e�n���.��V�V'�h|
+<{d�p��OYbd�w�:�Ơ4��(8��D5��r��\=��~��9Z���TT�c� 7W��b|Aãq�#@*����f}���7�vM9?��ؒ>ț:�SC9	������C.�C?��C᫋E���]yJ��έ<�8���q�f�N�;��|�[x!����~=�áb�!�n�}��ս�g��^B!�$ņ;�]L� C�sRU�6��J�5��6~@�@Am�b�c$��Ɵ���ښE$VM�z���Ȃx\�S��� �����rv�9�%�<ɿ^)�CtZk���8����lh����-�Z���a�j_M��*%�(��
t�B���oo��N!��:��la���l�DS�i�2�{�^T���CF|hh/tw�_�[�f{��@2s�������}����'�6��ձ=�������İ�@?(ȧ\�TT��*Au���wO.����!_r'���}�)Y^|\�yz�v6چ
8��0dJ��}!4�k�fZ$�铝]�R������u��|�S�ұ;%`���g�|�q�$�"o��P��
0D���*]���3B7��lTj%JH�(!JRQ�?Φ��j��V��ϟ��0��y��N 13J�2�vc�~���
��}�˹�_x�������ֿ�,@P�#Gf2�%|�~G;��9��J'���)MZҜ3L���z6`�8����CB5�r�~�@�I��]�� �/o�R���O���G��8\4̽���0jhٍ�.��ղρv�3t�*$�Nv��ٚ�L*���+y�9�>h��W��1�mE0����@8���i�H{�f�/Jnx�~/��K�)[z�&c���1O����g#�A��Ӹ�.5�U9��w�x	���{��X���X�k�k����\ h���$��;(�j����O gL=�W�#r�����Q�e/15:� lo�԰!�4�D��Z44�n��� ��~���J����WcE�q�o���L���NJ�9�vO���XO�7�4M~�z9r����hj���Z��I{��5˷��9�QG���*����Gˢ�%(���r	�5Ɓ�?�δ�q����}��g��L��k38�>���!��N��Ź]i��U��S�p�L�s�1�����'�<�$e��E)�ȗF�<���$�j�oþK�*d���=��i��=�D�ن+�b[x8~]U����יK�5��bg!�Z�sY��:��֚͊UB�0
'/1��t���'*'=]
X��[�DVY�`�69��4/I
t��G�3'�COں�J�����s���q�+�=��*���[!��cwE0�jx΃J{�����@5��v�/ ��uc[<�]�����z3���^�ܪ'�HM_��*�	�ꈑޫ:��`��ʰQ�#����Lj%���x��U[�<4�!r�����a�g�7�-�(���`�D�*��T���`?�ʣ�q����=�ﾻ��ed�3�gФ�B�����,Ph�ʈ��96TP�"�Wf|ت/J>��������mu�K?�C�,�J�]��6�s�j�+����d���8~�z��h6k5$ �&�I�e��V�Fd��y��*��T���}��R?�.��!��V���k�ü5'��$޲��a��)K���F�Q�l����6�g��48��Ō���}jt,cK���O |�\>1a��1C�L�;I�MT���O�n��
�9��o=.\2��	r�����	������.��6}�m1)GC�+���I��%�@��=Y�~5�E��"� 
��#x6y��*�j	�/����{�w��������u��4&�Bk��1a>b<�IF��L���*�W����Ep�M|��O�'�ce��Em/�H|�+Y��c+�8��U�Z�$E������2��J�7�������� 2CB��-�K�UV�r�H\���(_���U��=����}x�Z(��~�ѳAϴ�ߨ��D�K��A�X�]U�l� ʒ��{V(-j��@} ݗ���(��܄h��#[zk��ɐ������̋õ���t����,i�6���!HK~ΧR�ƷO(�Q���//���.fa}S���°�����r�{��M��j�d�aT��bV/� !~�!L[_Yם��E|^K	���K�PF۵���x���=ѣw/�B��`�ڦ\F���kQ8��q˚THʞ�	���b�|�%��!��L���S�[w%����t?;�6��+K9���<�BP��z�'���O)��S�ژ�:���%Qk�d�o�f�ۄ�x_6C6卄��$[�9���z�ܘY��q��	��`m:ߓ�_ސD��VJl+y�f�!���wh�����������!V�tk�4l��1t����,LGB]�M�b�"�PSH�MG�ǂo_�z`��z杜��øj�� �v'FY�:D<��R�xP�����G��M��+�|�R�Q�����>�Y��$WkꋂBf]�SCK����o��H�'���s�{Ia�Xc�F!(����C,�աi9���^���҆�vQC�����Ã��K�߈O�u�6.1�^�v��G/^���o��q~�N���F'�߅�t��.�On�<@4��A1��X��Ps��D R.��ǗE-�mi���!�Aw�6�Cf���_��{L�ȓ��ݒv��o��]���=��zmp�>$�����D�O?�d�R�K���:�k�������H���Ӭe��
j�Ї%nP�@a��i�yfk���"gp��{�����(o�G��R5T���A
�Q�S\_��22���vn��>�JM�p��b!uأ�IJ:�.XMr=�sg��.\/��}���uew�:�\G.�8p�Ox��M�o쒘��R�8tS�ܮs�+�HF0 �Vs�C����(@w0"��C: �.�4�1g ��^�U�5Gz��	`��ԁ���hCs^4�@α��ި��j��kV� ��x8)We��cÂbCG��"��A�"��L<��h�<��"�
�S_�b�)�� �O���E1Ɗ%��KJ�S�&p�ˠ�M�k��U�!g�Z϶�n<�u�b�����k��1v�jIE��Ø¿����1Y��${�|��-�k>�9��D���
��Mϣr�5�X1����"�i��H���ͷi���zZ�׍�9�J��;��h�+D���0�2
�<޺3���>��υ���;Z����h�����WQ,X����X.�)hi�x�w_	<~�)j�q����C���.��ݩ�~>iɿJ�(������w/v�N4�D��X�K�]���-,��A&��x+�=�WD�Z�"H-r��5Vr!*!�5qv��lk�LW5�b������\��/��K<�=�c��2(h�Ae@� �t��彆�Ϋ%��B��,Ӄ�L��B�]D� �0)eG'��)ㅈ�&�V��zf`Cs�[������|�G��P��.��A��|<ߥݿ7��T�8-�ͣ�&�\����Ff�-aՃ�ɭc��Z�n��m�|/�r�o��;>���%�;����'5{�lv�g�q�HCd�_��!�@��x䠟�1�#�$�ƾG�
��ʶ���E��iz
݈TS�,���oп=���h*�6�z����z5Hl�qhՅl��nW�Ki��	�jMt�VN�h��J8B�̗�`[c�JC��PD�'тY.�]Y�'�\�j>�7�k��QeIH�&�{V�o`��CL�P�p%Q7e�W�Y����t�A4G��S��06S<������7��&V\&u塆(-���t�˿����f���zv�z��TȺ�'���tq�+.q:�q��s�dpV&o�tX׍J��K�.C�����87H-�!�ް[�� %A*e+��L��pyv4�qñ��I[�k��,Q�m�$	�����[�����-T��H�m�<zz�����?���a�}��U�p@�uz'.F�Xmt���`��T�y�9�JGs��8Y$c؅��
A�`4�-�Ov=׃�F�;!�a��k�{5�S�Up��i��*�I�����Jm���Eq��!�[_����: H�	��T�SX�7f|
<2R�H1�@�d�&���LPJ3_4��T��-do����^�R���lq���jK9K0j���Ѡ�Z��2)��0�C8CCr9�Y��T�G�8
%�`�H+o�NVJ�Ʈ럗Z�#2��A(��s&�[-�'7���E*S~puJQh�o(��Ĵ��̛�m#M��砷@&pJr������N0 �݂th�0�s�~ek̂�~A-����O}j���� �X��Z�*jJ�/ɞ�xjs#�'��������o�Ac%BT[�|y�_����Z�X!��[��ɺ��m���7���oyZ��m�0����ء�&$gH�LؑMRX �uD!p�H?91rp�^�~&{O����:�7�R'5kEI�eJ���L�?2��9�������H�~�:�E^#K�0Q�B��z<vX�ԯA�8B"��`���M&���̞*�-�˵%�����N�����L�n!f��UQ."������q����4@�K����;ڌ(��t\n���_�_N�A_̗��5� �?6+��U�R�fe_\��pE�c˩����6�R�����߾PGSN����p$G�v��qFW�m2T����?oy��'��~O��6��S��4�<u�"�����!D��qԽ3޽�B*Zt3h ���������[��>��{w]A�揘V��9`\���AT���%���+:!Ҩ~�ם�Q����\�Q�e
��3Prnд���[_	85��!��ґ+x_i��'�j4cuݗ;�2]"v=L�)Q��v���
1�/�Z�|)�"A�h4n�;J6�٩��"��"qj��+
�u��;k����o6aД�a�s}�g�țh	������
#��5��?3R^�¸]�~a���/K��=~47�<F�l��f��Y���t|ι���xI�V��.�t���:S�q79QV�Mz#���D���V�� ���C�y�~��d�EE�dt[�/3\�Y�o���6H�YI�Y���Qc$穕v�p���������2�����7�z�T�}~�P\6�UFE�r�&��"L���#��h�I#
օ���G�����������#��}��N�"�B+I���ۙ���
 "�@��H[>�Ӱ�����,��[�����ҷ,�%.8�&��J�)��u}�g�lRor���BR�[T(/tԮk4y;h4A��#�>�ys�N�*=�q���>�6�5a���i�8�.q���,�vmc���\�um��r�.I���Ī�j�����C$�����}-)լ���)b�1�%.X$g��f�}����Y|Q�;v��բ<�X�z�)�\�c	���N�iv��Me�WP��V#�o;��1�nZ2q�0;-71�|�;֧xN٪�a�m���7)�0�KLl�&6h�m��wD�֮YE���nY��;I��::]��c�V�)W�S��;q|�`���x�V��s�fq�C�e�߻��"�°���#]��1��<f�N5�mM�0��W@��F?���Dst&&0��ux��Ӗ4���Dp����
��
s]ڍ$_��{���.���(��T����p��B���|J Yض7�A���L����<��G��l>������J"���N8��;�Ѯ���"�|���Š��qwJ\rb9���-;]����8�9��[0��r�CT�]l�,�8�x4�"���Z���-N}/W�aY�m���%�RA�Ѐ�A�Ѳ�N4�n�9;`1�S�Df[E�9�73�~i�9���9[�*����R��؄b{�(�V���o1n��u`Y��;c�t��B��E`"0.ϛ���Uh�a�ʎ����-4�Z%�2��K]�L�Zd�A��:"�}�g16M��W�XG|LVUH)S���(��un� 7�9>���o3V��y�vʦX�2J����rݫ4%@�/jG1Q��/�"T���p��A�gIQuV�
&�Ҽy��`��O���澟�R�Du"�1&�r�5��C!i:V �io�Tռ�bX-ΰd�i�������J�:gݟ>&��D܀�r�P_�F�3?�`���H<�`i+��+Wr�=է�a�D(�t�E�	��}!>�$EZR`�m�b�H(���.�K����Y�^d�ęH~>[�k|22ʬj�9Ȋ�A�N���s/��p2�!��&����ZsƑ��~�����7/4�;;(�:�r;@|������Q��Ĭw�/2�fl&l[�w���A�?z>��̷��v���摨�^��Ϗ��T�R�@����X���~s9�
r��Vx	f��s�}(�z��y�yl_��1B��뷔�)E�N�����F�F��Q��R�g ���O�����S� K�>9@����c�V>���lͪ|Jm�v+�Ym� �y͵��{6��� Bw�j0��^,�$0����b�����P�����s��Cˇ4�C�Q�+W��!~�&���S�p�XH����gMN3g�⊯K7n?oDϢ ;UUg���[�F���C�؁'��4���'z׋�T����y6�rf'_-�\�R�C�ejHkޑ������!�Ԧ����!.8��qa��Q5������B��?R���ߎ�h݁����?�������e��D0�{����<%D�/�y$��%�q(��$���u��3�?�Y�ti�fup�I���!߇SS���O[��%�����5���r��(N7PD�l�J�x>|�Les�[k���Z-�����b�^,�O���3���r�e��)��iʋ���h;�u/Ʒ�e{�/.H=��|�F�X��Q�	N�U��6��2׉��:q�l�S�b��p�u��5���i�ţ�g5�Q�U�f-G���#U�/ߛ�<�����e �Y�@)���I�J��3�ֲ��\�	;ˈX���1C� M�=��O���?�Ű\��8��] ݶ!<���G������xk��ո�!�6|C�BJ����V�9��N�@����q]�"��³c�j���(��iU>�2�;����<^Q���n�;@[��vȜ�+�v��a����7�Q䏁�OL�7;k�5y���/	���d}-�?��)�%yn��	i����$�s��ܰ��|��K�0ze1!��Z[X�''��}t<�1��=~�+�lʂ��U� �A��ЎIK���
�U�W&\ͽ�ڈ/�t�S��ʑl�A��!�l7}���(��:y�vVR�soF�9i��mn�))D�Q<Z���jGe�����6;"�OB�n�uS�S�����T�yj��98v�;j��"��G��g�u����8�����o�cඥI�� �{�x�pV�D��/~;�2$�x#G?E��1|���j1-���"�4�U�����P��ӝ:��
R�-E<e�y�I�^��dƋ���fΑ�5�p)u^�8�]�kO�s~�N�+��ɑE�eEG櫂�5�DA�A0yϙG!��c/-{��@��`o�@��X�71�5W�Zy��災eq{J/�>!�q�"�Y065�X�i@f�^ ;
����m��x�-2�$n{��uTԧ��n��8�d�C�p�[��/絜p6��>#1�	��%�+�F���+�6�G�Rj�3�Y )c�������q�7<�^�X�C`��թ�S�M�����-�[Q�mh�}+L����y���}�.�����l�
�5ĵ��m+����\��<{�v�)x1l�xF�b��i ����uM��=W`�(}"c,;4M%���ʂ��8����g�dt��N`8HDܟѻL[fDA�ŨB�<��i���v&�{L�I��T�{
Y�[���.:�	�=���9z2��n�����P=��ǘ����<�p.w��O(n������(h�����{����5��]�i���R�`��ǡv~�~�o��'|#�
����*�CF�f�kL����r]�3�����d�EQ�4��-�_��|���GQ������������.� �ˢ�S1���͚���;Ռ��ف����g��X���~��������8s1q�����fsV�4!t&F�Ub�;��J
���e�D�%��U�ԭ��G �*�ގb��oư��/�1��=u����/Ӑ���r��@�Z
�Y8�$�Ĝ�Gr���RY}���\w_(]X�Zlzl -�ͽ�D��uډ7��qR��P��j������Ϙ���8���1���_�6��9 (v��QF�F0?��[!G�Zw��j�x"!�x֐��1���Kdjd�YCa����R���(]Xc�@
5����*z��^��ܟ�d��ڡYS��{����8�t�GZ�O�*��B� $�.�ħ&�wf+F�7�����.aa��*(�>�e�/ވ�R�_*[�������s�KK�~Y+��Vٶ�K�CL�-�S���;��c�ĵܭ���׸�Æ���kz[4_�>4�H7�:��l٭/��:e�ymjNI-t��R�)=�/���rs�я���S�f;D�F�R���%�xH\� Bʏ�C�l�di�=����GmuϠu�/<_ȔJ����.S#?)�e��0C6�>>F4S�n^>�%I5#���X�K�o�b� 8�2p:_1!{��w>�h��	����Q�b�M���v��Y������>�A�)��	aӍ�_�B�>�f�Pn\�Fp8%r�uR^�4�j�
?Q�!�ǅ�Dg��"�|��T-�p����1��' c�ٲ1�(_�L�v����3+�5TQq���;���� ÏY���Bgc�-%��'H�W�QSQ[�B1�-m6��^����Y���&j$���OT����p�Ö�I4A8w1��_B}��o��b�j�#�o8]"Oo�̍�3VO�:�d��8� [���O	��0����J�g/V����
���Wy��v�WU�B�cd_^�
{�ޱ�Z��H�^�J�6���U�[dN\׎/;}�?�Qۡx4�V��b�̱p�:�V7%H�̅=� 5i���G��O
j