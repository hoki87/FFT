��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#���������l��U�~�׏O����j9�PY���`T���x���s����uí������P��"��b%>�1eτy�<�gܰ�N�Y�	� {��I�ɍL�ݫ�G�R�k��Q�!E	�5E��.��:�͂2��y�m�-�.E��i�����YS�
��@�H�ۼ��nD��Y�l"BU�.TԊ�=�-�����q���Ǹ��j��ԋ����tr�a�ٵ�]�b	��%�ɔe�)rYOjX5;V��R�������M\�	D��ҏ����9c=�Vͼu��Ro�P�Jf�tRvsY��c�"n�XO��	3g���Q���^�Bʹ�7gQ+Г���$�-��t�8�����A���<����l-��*�|dG�7�,x|LV����SG�_ϊ����5�ݰ~���^�����ѸsD}C��g�^S���
�<�6�FV=�X�P��ߛ���A�,��R�W{8
\&3�<Ϸa���E�~X�Hm���)�)(���f�5��rJ�� ۑ�Ft��Yd�]N]��@��n���!,W������x���L
H�뉬��pSkI���ˌ6�:�-����u���mEK؆֥�s����4�?�K��tfc�I���M|���6���ǒ�9�Ũ�0��<<����n�	������V���d����t C���	�=u�]��,^�ޤךy:�{��b���5�g{��p��F�И�w*��䃩�
"�y���%zJ�cv�]F!��R�n�W��e��n�k7%4���	Ѥ}��n��d%�{������,�zU�$�����"ӛYd?����k�<W1����{쑘�m��Ɋ���^��"��c[���6k����4�I!v񪰏 ��t}�I� ��4��:�ǎ�	`�w_⑝�� �"����q������ѮlM�s��&�3l�^i�u�]ᯮ���V{YJ�?P�E�CM�%�~I9�.���ra�+	F���ݧ1��(mi���dQ���Ϥ�`�`wZ!7�2g.��{Â�����~��/��$=�.���.6���7�?�KQVYJO�L!=���f��O�A*�8&�Ǔ�4���o8�}���҅�o:fLG�8�AF���P��8�.cjB�u2�b���»>��ic�栅^v�6��b�=��r �����"׋3�r켡X�D�y�|M�/ө<mSM1����╒`M�x�T9�|l��'��L�BOIܣ�8�A�	jоtcX7ā��N���@��6�k��v 
T�=H�9��d�z%���aB�]u�|4֫6��l���7�u
�ѯΧ�H��+���kѐ]�����D5P2���~���Vh�<�wxW-h��6R -����'�n!��9���!Pɸ��\��|+a`�B��~WZ���L�K�����wM	�+�����iƱ������ 42��������4�U��擺��G��bk�|T��o�
r�<)�i7JH���Pw�#�	^3��8��ط��<�5u�0W���6��Y���_����cd4�YP>��4����x�Ay��|��j\������&��&$)0s;ߩ�����シ ʟn|k�OF8oi��ot�[�q;��=�)�~{\�4Y)�Wx?@Ed/�^��(��)���6l�~�2>^���<CSO��Sl��w@���3���I�!��ڋf��[����Y�J�]��4�.X�AM�}n��&%
�P����*g�[`��a"�8@��CƱ86�3s�eE�<��Q%o��	�"�쥒�x�8���v�P��3�G�yX[kq��CP�ʎ⏖���w����v_��>ulK�t,�S���bu�4�j&2�R��#FP1q�r�Kr��-���P:��o���/V�c��~��4~-�4�xE3�_6���mV������a�)k���<uDŻ����Q�(�٘3�Uj9N�\���t�g�';��}-�0o��.����P�Yl\�L��D�9��cC� �c�9 �h���xȻ��ąP��&��_����c�&���~e��C��AA~�%�ɏz�ꮙ)�~Qb�vMhZ5���!��P+u*��5E�S'��TV�6CLB�6w�S+k��&���l���o!���Św����� мf��ˀ��g��z=	�N�9ܦ�  ��y�rWJU1�NSRc�.�V���/4�?	l"�*KG淺9~PT_�������{拀�l���q���rB))l&���.���d�����
H ��`D��Ζ,AoQ�������_?�;w�W�;��ٚY/c�۹Q!Zl��Яd��\�{�}��z��th��/m�a��Gi�q8sې���%�t����W(|�u����W�e����\t6Ӽ=�;�O��p���b����`FM������T`�܌j���!t�	��%�Ql�
{5�2��`7�#Vx�})-�p\�;�ku�
��8����d �|Ԫ��Ld�.B"���	wcPɸ�;��+�0ebXܰ�j��N����.�Gxv=��4/k�o�0�G�O H�HD��ь�[�[�1�I���.4J<=�9��P{ d��EM��i����̙�XhUQJ	ޭ�k�c����*d����z��<g���4�
�0�* D�wHp�y�,컽7,N(�|g�����<�9������1�/"������7�jPb�u��0�*��`٢V?����߸ }���.SWj���y�jp*��2yn���*�bqq���1����F���ʯ� �s��ۭ9�X�q2��GJ>=���.{e��#���s���%����wiw�Aƪ�7rGJvfDXL}�	qP-����;ɅQ���;�^���$�G�j� ��i��~k����oQjp�l��/�^nt��{�ϼ/	��n��9q�+�&���I������f��<�3�lgȕ��5����!���1�3����{3%�v����>>#�Jψ�	]zV���N�bX�9}�ܕ��g�>�$t�����s��b��4��:���b�����%���mÁ���z���~S�6B�?z�	���ăHw��u�2
G�a=l )��"�C=w	�g�����������*��"?z�xG'd����ܼ�&g�9������P)9 �2]-l����9�D��WI�,����Ck?.��=Gd�������� e�q9���2�hF��St�|J�m�A�޶�I��/
�
>���P�9!�[�]���J��l�q��Pz@ؾ0�i�}�;����_N��c_�ZrX0�;��%/�0(���C��E�E>�51:�
/F���H�������ݎo�"I',�L瞈�u�̲��
L8rV+�R9��%�!%�8n7i��2(�6�
Y�H@�rE+VA�L����y��6q�g����V,��8
O�o*1�������@r�1$��-3{lva��V����v�XP��b)��aQ���#:��J3��ڶ�}4�9	�c/C��So��>$� �L��mɠ����5���x/j���D7��P����S����Ò%Vk�Q��-�W1�o(�n��eOb��#v�۷�r�r �&�}s#���}A㵰�~��~�*�ٛ~��w���v��������5��_��G�=*�s���۠^�R��u�ڢ�q#��,��|O���<F5'rFgA[�[S��ðc�hV6+W�Ī�k�:��$S2,s��j�b(d��.56	�A�:E܂��U�isb��d/�D��������J� �87.!�^�p�h�A�wpz9q77W�$K�ά�#�{>J��3lWxt惇�Y�@� 9�%'/��J�Ħ;�%qv�t���Tvi���b��tz�ޥ!0w�~ ơ����Hi��C�����,�LT1Y��c���j�߂E��ɴݗ�i�#�~�)c ꄡ���N򙪱��y�t@�������+���Z;&�p�Z0@M���ރ����n�ь���)M��� �m�g~eZ��'����G�?ٹ�w7 l��F9�;�I�Y�QN��� �o~eV}Ƶ��?+h��i����l�W���P ����x����yF��[��w��i�n���:%��{!^�`,+�j�� �v�|K���l�8��_��xpq�+�_[��n�*�bk���|,�լ�X5������1�7��T�t�� IU��<���,��|���S<�g�#*\�F��Z������_��5:f���L0u]�\>WN���x��JR�l� :�ݭ��u���!�醩�W;�G��������C�Dr��V��%/V� ä�7F]�.duj	�����ˎ����[U�k� =� �"������~�������A�G]C_e��������}�F�Xn����=�O��PK����eT�z���V}�>�~	$u}�C�Y�� �4�؅'\�.h�X�?Bך�1$�1fNA�}iԏ^й��ت=Zb�}��@66��RZ�,�Щ]pU�����9�w�M� f�[-���+��%���T��b�"8��E6�!���>�J�|�5��s+�)T�p�-&�;s�+�~�H�SǺ�k`�g
�[�j�?�mlj��C�G��HV�r�.��ݎ����ʦۧ*�1k���ML����� �����1�קEJ'�L���k��?N-x��Z]J��NK��q	�'��RK[D�j���K�;��d�G�!|Ϯ�D��U�a!�;W��y�(�N��dh'��G!��c�,��.1k�Ɨ���5��X�׈Z�[l���g�V�sc����x�.��KX����`8̊N]�]�*z��\K@�~�>�X�rč��ߚA^{i�7K[>�r|��l��R���yF*�_��������&%�0��S�n3��B��Owr_�u�Y����H'g��w�/��2*`�
�r}ppP0o���9���R��,	D��?/#�N�hc�mڮ�X}m^'�q]�O8bi6�a�hF �l�S�b��ӇԺ�"�Vu3�I�������Ͷ��^���7�)����+�V@�<:�?�ɘas�0�'x�YRL�ׄ����c���W3������O�o�ȡ��W���m����Yԏº�s��ᒄD�7.4h��w���30oʃ��k����P-w���'	x,�"��ι@����\S7l��� Z���Je�[�c��`��L�OY-��t� lD׬V�-�m��tP@9W�
&���D�d*h�h�>w�,$U�d�@w�����N��s��?D<�7σm��{ٟ/W��q���ۙ_�j�	Щ�{ΘA������>0T��8ߙ;􋑮�׊Mo�'��ַ���CJ�$�<�D2dz��*|�ؘר([P���	��`I�+�~`�jD�Ѳló��A��^q��.,d�׃,L�����%�38\_�dH����:sN�E��%���g�����UƧQ���|����1QV�����ĺ����8=cG�M�-��j���٦I_��)�u�4M\��Qջ�lP��<Z��Xb_=PEV��Z���CQjba�1��o���=����q���AK5����N��lh���4�����*3����1�~�{���Zv����<'�AN��b>܌K[k)�N9��/���,������.��n	6���-�D���[�D/l��L��l�}<C�rtZ2��o�p��K�����X�*��f,�'?�ȮHT-���+'}K���<�e��re����"��d�E�!����k� ���<N4O�B\W�Y-��-�Wi�g���S�WD�W��}ԖͰ����-�Iҙit���O5C"��24![s���A^�g��M�MHM{�i'Xs�2�eAn��T�(�H�E@��蹈�H�.��
>)��i@��t��q��)�!�̴$r�i9M@��9����d2P��3�:e"� dba�y(��B0.��6��fA�$���2<�W#������a�y��gs]��g����ɉ�c
8��#���F�WB[�ʲ�⳦vD��8��o� C��D����.W��_?S����B�zǠ��`����kkGx�"�8�l��4ͼ������U�½�/e��2��+@��Ǯ>�������lM�a���Hwd�4�_��㸏���3��P�jEZk1q�}�"�M����t����S�4q�x��ume�Lv��nR����4�DT�U���͓1", �6(PR~r�5y�<��
�?җ�5������hp��c�X}����IU��z���N��A�����c���R��Wst�#g���Ҧs{Bz|������\{X���OV9�b��HCav��7�U��k9�8��#��x�q�D)ܬ�q���K�ł�Hh�s�c�Z�v��̩�J_�7%cy	��W��Z�|jɅ� ������3lU����/K�O�=�^^��t�?�&F�z�Wuŭ���ͤ�0�o�;���/�m���^GW�#���G0��L�dl{|x_����"B�9ﴜȁ����]�)�
&r�M���bk��w%� E��Ҫy[g��2�X��՛��s�~:J���ų�����G4�&UM����&72~$�n�)C��^�}�wKq0�wHK�߰T�R�P?�4xQz����Ogl`���Bpt�gͣ�ƚ�@ע�~�:b >�3 ����B$F��+�.j�<��JA� [���kH�:�m]�*��'0��Um�Yz[ȿ��KG��f�R�I�ug���%v����Fò�����at�$k��������n!�A)���5�R�"D�ٖ�� ��^@��Uc/{K��
�3M��{k@RP�W�4_=�$Rʜ��I�N�2>��	A���l.������A���s�3:ޜ֥2�}�0��=`���`[�վK�e!5�x��gd�(2�/C\�Jabu�0����Ί����IƹnjU�EF ���,Sp��h�@A���C�V$��LۛDat���2���������m|)�[�3̼�Z0up*M����T�ia���+F<���cp[UV]�_��$�`���M�v�.�� �����F��9v�ɹ7����c	K���P���}G�ޛ7��C�����-�G�)�2���.^׬����C�@-��*��Ox�4��g�ё.��5����m�����e�6��#��v��l�T�
�UĂ��栨B{?�p9�*�{��~"��n�n&k���8���Jq�T��jЩL l��=w���ͦ��"@]��� ~��\�{���/V�䃹����݋����H�
��H�R��?/]�_��H�纊IC,a(Ǆ���x��c�琘[��]��°��4���r>h[ 	qq1]fC]�\V8\Hfi����1#pu��g��x��5��u ���Xi=<6=f30��hB�I=�[��B��b�Z��3u��,�a��y���Ԩl��XmA>�^�y���wG=T�[U��m�QA��x3�]Y���(��l7H����'>\��If�K�Y�[�x�@v~����u8�~��&�I=4�g�e�F��#���*K�9Wu֍u�~�x���ʇg�����n!��O�"�5��ȷ4N�>���,�#� ��g �4S47s6yb�یj�+�a�q�?*HB��P�e��~A|�׈=iL!�%(�_Q9��6B�9�������r$��,I��\�,b&Nn��<�e󧲖��R(<��H��d�LC�� 4��@����2B!P�5j��*Q��&W��l l�n�8��p(@�2$�Hkk�:Qݞ^�z^��j�����b6��YӋ!*m3�8�W�9qoF�ʱ�<$�l���zw9d���hI�����^s��Ԛ�GZj�lx�B��� Z�|3������`��ՠ�����E��D��"Knl?@��!c<X{��ibe����EE!<'������	U/���MD9N���Sz���j�K)(�.�;�
r�q�hvt)ro����0��@l�c0F��n1��Z`g���
��.�*:�P�'�o��a�{���GB�ڧ�����@|US����2af�a҉<M��Y%h`��I�/B�-PV��KZZ��vRݵ�(���˝�w�vCgܿ�S���I����*(d*B%"��6cU��Z�d��\���%1\|snW!�B�AO�v�a�I#��8?��\H��$El �f˲L�O��j+z�����.B[ɹ3���i����,�Oy�U�m�\���{Rk"���(	(M%tPi�S�����iT�U	��:�Bܦ�i�#��M:����Q<�8�\���9Ιn�|`d��y?��U�8�z���ܠg�~k'p�!;B�Q:BJ�<�����b��G�W�("B#�ˡ :��FVY	^�מ�V��l�C�&'�����^�����yW�0g��Ù/'�έ!f9-���{�r3�r/�e����V�p�E�/��W^!PV/�h���A�bG4��m����+�I���SP��E�٭"E�y��t�M,,N{|N�tk��-~BK-!���󊭈���^�~�&GE���ԙѶ��tߥ��U��	�����k箆:�n��[��ͨ0j�5��G�L�PdN�HmQA�Wh��U!h�{��%]/
хti7���(z㡪�4��f:-�����(\6���(�E�e�X��{$!-j�~F�I�ߍ���Lt
!o���)m�k���$o�'��b
#���z�F�=Q,�|�! U�q����e��f�Xva�s�J�%�W�25@Bf���r���<��WΤU^��Or���]舡��m�d��t��W �C�0lDI��-C�peS�|��7ȔT�T��.��q(8��)m���O��&��������S}�ع/�}��Y�կ�e?�_�㣩Wڜ
�z�ǔpcQ��r���22���1��E�����4�v�����'i2�8٢�s��yO%�ľ�d)/|��/l��{��������xQ�����0��>��S�=�q�q�Ԝ ��_3jF�/�!��c�-��0s"?�����~��5o6 e��WT���P!��%X�!��|g4:����o�VƆ�wQ�BCe�i�?R�i[7����#z,6 ����Mz=���0��X~M�����=�ZJ�hx=	y���tLQb��#��G�/ݡ#7;م3�
���a��
9�Ԗ+B����<�NkҠiȧ�K�b��%5��/^U���v��ș�������R�MM�:7�"G�`�aNS��С�p�;q&�x�)6���ߦ��B�?���`Q��Cc��o���HO�_����ˠ0��^���# �x���V���L�U�	89��$3�����l &��L��;J�B0��<�SX;ʄh�#O6�	X�!Jz7��2qji�l�ܭN9=��"/���{7�u�G`��A�OS�M9�pX���IZ߯�i�/O��Э!Z�͋O��B��K���ÿ�y1��0o�e�
gvP��u:��8	�q�7$�K��1�Z@��*%����
�{	�h���9�#�<�����׀m?@��������b�󙙷�l4���prD/�1���!%���W���ܵga��GT�֙e>>WA�e{ame�?V�҄�o��&��Bn���E�s�Ne���8�Ѯ�c��8����cAu��	�O���^�1I�H(ݵmG PWy��ĕ �T�J��zj���Z��Ζ��o���u��u3Wow��4Ј�ٝ��Jj}nMa~_����'߰��߈�\�cP"�����1h�	�3Z ᇃ��?�
rXX`�j��*8��w]`܏"��ݚ�����îN�n�� `OR��4�iro�D�..�(f��Z
�� ���Hb���{7I��{��Ul�r�W~�e&���jڱΕw�0��*v���TQ�8�<�(��X�A[�X��M�5�C�ZG
���t2HbڡNaQy5n��Ҍ%B_hД._S�3 �P��_��U)����?�^U7z���&�HU@��+�Bsil�Sw?`��5Y��&���.�u�	�A���_���V�[6�	�៌����h_�o���m�D�ں�:-���	�c�Ӎ����v4�� wB��,Q���B-!�$��?
�x�!�_:���e��@5ѴI�b���an���jȵ>���mT�I.u�m��omW�I��Ս%y,Y7 �<��?�}�Lf�S�F�s���s�kx��V�S467��IyǸz�⸉`r��S��ӥ�4twQ��6�%�]�X~���������_���̞+SV;�u�
�װ�y����:�̽�>�9*��U�o0�xy��*aR�?ee��NB`�ׁW�фnv���>EE��>���S��������q��W��;�;4�>ɣ0H����$�Tۭ?�}lk�����t�&y�@ʻ� ���,�u�xֆy�uȅ��,	N���2����2�^��#�SjMR볖��Ƞ�˦�p�Eo�A��=0B�[����,�7�A��C��i�Y�^1���O{���"W�ya�cg���Mg��=��,p���D*UbE�y"�aC�{ea)�|�|R��������y� �=*!�G���î��E$������}��23���M:ri����Z�^q�����0T�.)����?"��Q ��!������'-�ٝU~�Td�����&�9,���OL@�ɑ��7}��m��

}�C%l��%�@�C_t�Bw{�r����y�ǳ*�;�>�C%����^���?������_��ĵ�z�i3+�����3�A�G�9����bf��	�"P�:��S��I���~V��r�Q��e�.��� ��Nd�/n\wIyNj���g6`��"v��1��M���_#����3u��{60^�OgDS�8[G�����1�9�)�u��P�~x��=�TL�6 �ng��&iG,�(��[��pf�xј�!�,�4��`G��Lo�v��Wɍ��W��U����k��:5N<PML]��,��Q>�X��{��;�-���)�A��2V$�0�ya�R#�v�H��ݰ��b�׽�cX�'x��ԂPqai �H�vZZ߽5�sw�7�=���I��2�|��L� ^�
�a�Ϲ&9���:{���,��_����7��n�z?�m��h8�HE�me�]���<�������� �,5�j���K ��R��(�Hx�O��D�OWu���hW���ܭ2|j1�_�r2��8�-�IT����i#��Z������!��<Q�O�Q;ZR�U�D` ��w#0��(���]����s=��g�Z�.٬E�16~:=���וjc%��*F�C�z�n��4��]��y@*����7p�j:e"��>�'�<��tx;�/~04Qn�4�B�Tb{�^_������ԏ��d�_w��/��,%�n
S¦
Kz��⟗L�i����[�p���C��W����J cQ�����G@-�W�x��Ƈ�X;CU��#�$��K���*Ǯ�P����@��+�"ȭy���G���HI�#,\�-]b��)RyĚ�ZQ�LL��4�Oz	v�:2~>��!:�N�*ǔ�e�'O���rÄ�TO0X�=� ����*o�2��&��B�:!c�+e�D�	`��z���:�둌�wn.�+�h�(1~hM�H]?�����Uԛq ���)��`~Y�����L3����u,�*E��s��[6i�˴����b��X.u� <��sm7Ҋ_�4H<
�#8T���r��ߤeDq��jC2w��'��ĝn��k���u �k��Tt���x�U1�Q�"|�nWh'E�*�W�%�_�*�x7TV9�hx}x�Cm��/�'0t7�!7�VM�&Fk�p��!���׸�ս&�	�l0��E�L��7�u�B�y�*m��9���p5>FZ��0��Is����Ȋ�y^�<�g�h��T�uԞ�I�a�´�eJ�s�����*ٕ�j�N�3�B|�.D�Q�����B�-�]�s���'vD�)<�k.ZH�5�=ŉ�9cg�L&�K`$�xc�ќ�#@(f��D�D�z	h�{��@�˂f�acVpQ-Yh@cy�SԹb ����U�;��A謿��FГ�z%\D�SEc^J��T���d���:�D�q��D3;��Vk�X(�ʹa	3���������Y��.V�֓~Q�D�4.���/=F�u#%�O?���ƊQ��{ׯxUz۝�;t��a��p*qQE���+D2ۻ+{�R���\nr����ګ!�</?qxhfZͧ��&���˯6���qt�v�c�y����U�f�(��m[<����\���3?��(�@�k�P��%�f'b:�&_��c{^�K��Xf�ꐯ$���w�#W�u�N"Ձ�����}+/xaW~tױl�w�ZJ`r���0��x���-2pJ�=�����l?��d9m�Gns�mr��gqs��ds�oM����lj{��S���P�$�|���nA�V����&�J���l�KE�ÌE�y;�����S�7��`U����{����,�㙫�8��"������{+ɅMDF� ��gfްbBo����;Me�\J�3��H�fKA:*��d+��>՗Z�:��⵭��)��Pi�5~�/1�������I,R���\B=�C�p��;����zoB�����!���
G��n�V�x��̡�������4{��>Up\."��9xn�����c$n�[~���cL=�r=�6�*u�!z\�P��A�aܺ�[��`b ,�����ѡ��)�q�`k졦�@��Z�U��Z�u):/q�����kb琽/BG�p��W����Z�Kt����I/x�A��_��θv�+�ر�$�z<E}"�ڡ�+=&J�=O���T�N7�Ŭ�4�zU��#��z�]x��2ǢǮ?��)>��R�>�K��5������
��b��^c�ȍ'~m1���b�^,9�ܥ	�#��z+��|���gQX�k=���Db���0M.9��(���>�t��	f(�qډ+:�b�ĸJ.I)*aN���1;�-e6&cG�ǖ�/�M�hRxݡ�5���Ďp����j>������I[p���*���[�B��A�S:�4m�lg@_���?#�%�����e>)�Z6�9��7��p7�˱�O3��t�+d�+��k����4f�X`���7���DO�pY�s�����B��{��`O�&~����J��כ���%�����N�ẗ́�N��`I�����k�p@�Q2�P�����jU������D������e2鐔}̬w^��lj67]^��SVlMyK�W=��.@iH3��e�θt�3���E�"U�('Z� �N�-������Lm�]��N�@	=��!ߺ��"�(��1Q٦M�W���(� �Q����8�tP��LJNo{��Cnb�͌"���:G������C�4�դt��=�� H���2���V�7HsE�� ��!��a�W�,w �ݙUWho�����Ť��1a���W+��;��Ix��un��l��
��߻����P4�n5f�Q��b�H۠ۖ �	������S����uӾg�	G��ՠ�O�tg�C������Z����/�����,���/�����t�2��W�{�}���I�V�w�STY��G�BNY�#���=�jee�#y*4�����D��p�/���9W�A0ʺ>�L���v�hy��%�a�� ���/���ı�ŐZ�h���V��/��Cei:�R��:�����K��74eZ�OÿiМN���7�� �$OPcS���g�����˿���Ҹ����ʡ��\t�a����I���Z1���vn��5��L����ފr��/��Gs�w�B�K��� ��X�\Ǧ�-'����Y�tjdb%���D�5�����X�@*��?X�D���X�>���y6.���:��W��q��<��Ҩ��P��%�wm�]�_<�Fw=Qv|H��r����;%�n� L��o�&�x�ԝ�iJ��.҉��%QOh���1���E!�B¦���Q=Y���P����������:����d��9K�lP;P �,?S�� �0��[������=��뗋����|umIm����ˍ�H6%��t;��q�yt�#�G͒�w8��N�(�힒P�=D:�?�bSC8����I79ش�8�kt���[`���ߏ=<���z)�.�����FW~�J�;��P�U�:��I���p9�P���Q�T�WW�����[
���3�p(7�y����Kr�6�b@-�eWV��bw
1�g�Od�}���@㮂�:L&z����%�~���V�+#�u|�t�uv���a�t�!h� �!��C�'~9��"�Nh1m��o�'L���$������
�9�R� Y�:Ͼ�\=�\i����35syo��9�5���*D����x�(9�ա)@o�������ϵ
X��g���P 7T~��"���4��Sa��l������;�&��7�96�;��@j�����)ʊ�Tb#4�| P���@�CQ?�;����=��р�R�B�&��Pp�� �S�<=�s��O[�Z� 2�"ڗa���H�%ŻF������V�nMR�z��)z�qI
l}��|Z:����ZC�n4�����9�2�h�2PF�G+���]�/^3'M���Aw��8:GPY]g`�-u����so�W	�H�o3���(mK3\�7��c׺����ȈxQ��F��Z�nʄ_|��$@�pڌP$Z��YA�xGk����m1��ބ�R�h�A*�נN�TP2���0:MiߒF�D11{��v��;��|��
pw�^����#.`�Q��q1��L ;o�nkg�A»?G��C"ܔnK��L�4q��>ޭo���0P˹���hq�o��J#3�'�M�����TK����T�:L@�4��0��*��w�Jj|���a�pA����L�ĤQ���Aa�S}���bz��̈�_x���4�ͼ�L��u]Q�v4����$T~��G�3���+��/�!��zK.}7-�U:���R�Үw�b�G$\V�����u�>'����Z(�4����C.����:_H���3�a��!�{�a܄\�)�<q��K�0��Gi(C6Z�iݖ���b|	��3Z��:�g�Cc����'�@��@Q�4x�ظ��I����@5Y��?+�6��uE0m:�@@T��*:hҕ�5�~�F�o&��W+'L�����'�����'��m��*���L��E{s���>�s1�i��Jv�0��i��H>?�}�R��ϑ�H���F�nQ
��`>#�����6��F'6K,�h]l����c$�����������tRm��>8wJ��7��GP�]�F@z��"_K5(����uݹBͳ$B��^?9��A�K͸':���C����Js }���3��G��:m���y���	�t�9�;��Ơ,���4�;�Ԉ@Z��!� �!�u*�n�{��Ȕ��f:B'Ý��s��<��y�ZJ��0��di�@����Q�º�	OO#:o����ظ*��Oko�C���[�Ǿ���KKluE��/��B�n��az�U����3ҿ-�}#����$�TƿN�� �x��V�{��?�xG��,M�$m
����.d�L��SįKF%������������gh<�HU�J.~�/ ���Mɓ|7���{����6�Y.�F&
�:&yj`5xo�ʀ_f��b�}��'o�yzN>�R����%����O�cco³H����^XGxx��Gw��m��Z��,��M��;-=ꓳ9���H��e%$���$����|d�u�,�k��]��֛ע#�&O.⁶��p�-\k6�.o_~���o\S0Kv��4��U�]�G��ί�j�C!�w+dر��$�[!2�+��1�~<��z�v�Q�]���,AQDK��4��\�Ŀ-�5,q�ix&KI)f?t�����˞���bL�v�,v����Hw�n�&�(v�Зw�	c�(碩��XJ�c�3X�� ����&��ꢌ[X��íI��47��r��A�&huE7�y�v����R�e�s�dk�@��B�׾|���©�m͌Z�3�ל8�E6��i��?�
6��v�G��މ�:��ł��	���f��3pw]��%�}�L�E�t���3�2!���G+�Z$d������nω��Ė�3���E�7~�q�bڹk���SU��m�뵘z��"K0vy.������79��C�R,�l/�S � �_>�G,���0y(׸�Ov�h�n1! M�X�y�1<�����-�JT�דR�����uvfJ�陉M�7�ѩ���+�͕A1�V"� �A�����Y56	�y�o��Ğ��xde�@1��cJg_,��3$}[�hE�	�o��z�έ�y���ˌ��U��N���Qv;ܺS+tj���躝��s ߀q�ٻ���k�=!J���_#����&qc����6�z.����.8���n��ZX��ic,��k@�o]�gC
�$��r$��L`������5;9�r���:cC��~��K��̉h��S�xXz�0�k'��,
l}0du�1�{�
�V�4�e)�\�"c��G�������: N7t}Ш��Kǣ߼:�0R��i�h]d{���{R�	��1�^�ˈ#�)���np#�l�e!��nr�iA��#<Jf ��	'Y�&�:�tod�,���ޜ�1�ۘi�g�P��1�?S"%_^5mzL�C�_`%�@��4&����+o22A���`� �'V������8�w	$t<�-�ɽ͹Ǟ��Plx?�|3N��`:�=%�.^�����R�kɇ��;��#Eq��d%9i�B�h���jj,RTŌ���lh$)��-�4���<�R�ә�3q�$��DǿY��Q�u��$z_6��N��j�F�Sf��-�C�8|hHр���)h�o�$q�%��/�W�"�� �C0���%�tm��δ|]�}�/ .Q^+�hJA�W��N�oJ���,�5{��7ZFz���jj/S@�Ҕ6B}.�=������ ˢؘ�A�Ad��H�|�-�w��%B��)��%��4�a��>/^��B��=��nRG���9mJ�'�u�_���C?.���L�����UD�.�/+�O��;��e�>�3���Jf=6�	ޡ�-�GN��P�%�ae�J�ǉs�u��r���Y0�
5�3W��mV��;r%1�@�={JT*UHh,2����ݿP�`����0�y�~��I��{%�+�u��m̂��=�����@=�<�&3 g�U4���ϳ�����H�d�-/B��� ��2bo�Ó��8�`�Y��S�.��d.n��>-�q��:�i�Y��_�<�(w��Ʌg* Tp4�w�ư�t~�����yQ�;H�p��I���.�n�wN��g��u�����S9��L��Ϭ�zx�#�i��� �v�gv�l��˖4浰J�����O����j�q�yf�A	�f��s>���8�ɪ�_���6��~����	z+�9�<7x8��P��%7����s���N7�vN���ӵέƷ0\�N�SI@%;�
�r�v�����}�=JJ�2�&/�B/[��=�Dj���Bvg���+&=J]�HH�<�~9���$��6��u>O�Ŕ\<~&�><L�K(Qh���u��z���ػ��?qyRcL�׹UrH���T|N�hv\�f�!���^R&�qb7�	b����˧|�t����cq]5l��ݐb��n�;���,�
�fj)������:X�Hv�v�j�ge%�E ��4���R�u&�>��@���<�ń���/��-ބ��U<Q�P�}���H ���å���ULb��`4�B���d,Lq�ғ@���ݳ��NrAВ/기`�O�rݺ�l�K�C��S���'?�×�ѧ����)G�,��$i"���|�k�'���\���>��`�x@W��!P'�l��'͹��A�������3~����bǲ�����g$UMJ�eɁ��Ӓ��<H����Z�K����J�ǸTa��-��� 7��ѯؾ�HR�=��"D,�7��],�`b�ۼ��(�e�0��p6�-���V�ؾ�-����9�6�U�0�|�:@�����$�p$9���
�i��N�b*-떤`�o�+��%�k�~C����l]O�P�2�т��k��~��8�6*I��DV��s��_����N #�V-���B�B�h��{^�7`�R�>� (#,����g�v�o_>��O��Z=�����0"��\����&��\?�)K����KH��M}����[qqu�!���"�HS���_~ɐ��B����+��o���̊1��i>
m�\�ʬ�� ��>ߓE��="Z!�'cF��e�j�_���f����Ke�\�F=?{��l��Zv���6}y=d�_0�R����{��^VRf����uRx�Q�T��`ة�=| �!2<ך^�j�d1�7l<�a��D��eOl_ک��hfh�s_D�����JB�qb{���K�EϰY��=kh�M''�F�
'D	K�ߐ�����}W$=+A��_����h�J^�8𗿿���kx8����=�m7W�#=Ɛ�f��1M�\Z�t�GߡNb��Y���vi)�|^n��w����c��+�-���>zcR��c��B�j�=�R�?�V�P�B���Ӄ>dqǉ]6�rNSە�&���/�p�@=�;�)�S����5bʵ��U������x��Vt�7������Z�#|���=4`	�j���N*����1��#w:ΞH�y��� ��)�*T�m�)�%2�s!�P�6�X�R3\ȟ�+�
����*&�a�	���)M�X?9g�\b�-)��� m�`�j����]�>O>�{ӗ���Kp��|�� w�l��.�/*$���/"^>�|s�t���'��
�k�����T�1�	Kt��E��Xy�0�8*���b#���u�mc�+��1�*�H��ʷ�E�p8��lwc"�7�e���K �s3o�@q *�.G�IGM�h��6�]�r&eͽCb��Tj���7���v8�6�͔z�O&��3�,�L��Gd��Au#Cx�sĎ�8W�>ɢ
,��۳�<�su��˚��Dw?�~�O��j2�ơ1�}�aj-ϋy��j��
yEA�����|�Q����s�p 0bL2��&rZb�G�X�[H���b�K��Y_�4<�.\�Q�k�I�E^�
$ں���FQQ=q �١�3{'��wF�" ��Ͻ���%�Ie�f��]Jd����1�[���<������J��s.�����	ɬ�K�ڬ����:���#�X�(��8�"�7QEY���9'��q��L����Z�k�����R����8��(�[��]ړ|��6�i�Q
�7y��2���g%��I<�����`�v��#s��� �mMŌ�vI_�kΊ���/�``/E(�T������ѥ%�)�^iqI�νh��=b��2�=�P�El���+�L��y�/϶lm� �}tI�,�sC<^-�(�i˳�Ab&�	�8{g�-g�0)�5e~��ˁ;����Б@O�S^$�&Eʓ��ׯF�; �W����rK,�l�ŉ�̢R��%�(�Y50���L٧����[T �.��9�i�q������/Ae>��b��ErO�[��s�R��(��ׁ)5쀢Sd�O�B?��
��À!����Y�V�zpu�d�$|νz�HY^�:���2�s�ϼ��鯍�ל
(���;�dO����a&0:��O>��*�/^��n��+�����"��ܒm*$��S5TƓ�d1�:�]�E��]���,)��م=O��af7Xtɽ^�ᅃReN;2a�2(�����s-�����s�S��V>����r}�:�y���V�:
Z��	,�&�Q��eLN��NYY_�Ӵ�]Q,�}��QC��\P��˛����s؈�b(�<k
'�.���0ݺKق)�q׭�@�
��J���� ��d�����o�-�{��D�fW��qBY�,V���� ����zQ�BT�,ˀ�%�D�
�༜s(1���0�[�9�����C�4�a#�V�z�[x����"6���(aniL��(p�<�& �Ec�	w��%yI�(��&�df�����A�Q����up�ݖKp�R��
4�>t\�.W�@/�p�i� �k��K�n�`����+���1�➱��MF_4D��*�dTR�����S���qsj�qn���H�<��^]]������^d�P�QP��������Ku$>�a�V��|�z�o����՘k`�2+0��^o�*D����2`]�vj�`�c5�h����y����6�q��A�@�~�Mѥ�-��*�y�>d���<���K��2��u~���Y'�K����	���OV?>1�qO�4�9Wb��^j`n	��8`Ed��>?,%�:�L�w�b��'o����z	�O�2��5'k��^[��C����������G�7��L��+l?7���NI���O��̷�������\�����
��L`��7X�Tߖ���m�J�4�Ȫ�l��=)��΂���Dozn"z߈<�-�\�s�(ޥa�3�l�����'���Rw0\����}n8��[�D[n'���F�N��ZY��E��jԣ~�XA9�SE+���7�F%�鼸��;0�d�e{
]��Io&���S��RNf[�j�-}��;A�1So1��ؑpY�h�\2�)f��byX�f�O�#�4C��C̬�!���wÄ����Yc&�vhʢ�)�Y�
Ƈ�u/���6;6B�� ��H|��N$́�V����_@)�/ܫ�{���(::lk� >!K�������s����Ͱ�I�p�g���d�������%p�C=c��E����l'�A���q*�b�1�|F�{C� A|��J_)iC}ߨ��Y,_�3���O��9�rJ�g�v��}�v:R�Ţ��~%�ˬ3���������$��c�8�f�5*��O�h#�4�-m�	A�!�Vo��m��U�h��n^(L�5UXI�#�U�9������	�]���-��m2�fuN�(��C��%al&�Y�XeD<v��ӽ@� Bi������g-89��A�a2�2�;��!a="R����l��mFt�&�s*S����Z,@ 2$��U$�[�G�ton�S����}�RS�
$���ɞ������4p��*�n�h�r����a���߶΂kB��D[_�Y8$9Ne��]�\�s��sx�jzb�����e�:��\Q��H�<]�S0s܋@���iDFpv;��+����)}v⢺W����b��\����ǧ��4Ɂ�έD�Dc#|���U��E��z�Px�LE��������]��hqr�%��	��(�����y�W����ٲ��;0�9be������7*y��"�h���Aܸ9r��5.c�B�@B��<q��[eρ½�q3���LE-n���}W9��ɜ��"���u~�>�J�/UC�b��mܒ���
��*�n��&�<_�����홳�x��Sj�
���?�A���nT++�̓��hL*��|��&j��0�I0o�q�����^�gA��SO��j�
f��|�q�0H�y�)ǈ��p�����"6'gH�M&齦M+��!+BN��DG©%-U�(U�9fzxw��Պk;����154qZ��<�X�t��0�cj�p�W&kM�eMS�����`M���}c��ad�p�+}J��u�z���>�+���^���.�8�-���x� Q��Pc��*!*]B?��`ّmٍ���A���_7�K|��6>�� W9|�E�P2�[������I�1'+�c�˂��I��������� !e�x�8����##j� ��n��q��Ũ�XI�1�c�s�~��V����	���L7Iv{Q�`
�u-�s�>�2�4TpJT��n�u���1"l9y�ho�k̎�Ȏ��f[�d��3f�
ŭ�C��`z�S(��q4��LTƌO˲�Co[-�F��'��mK��VT�-ΊIK���;a5B�
��j�������k ��c:@��M_4�\��\#7/�59V�Ҽ`�����1I�����/�p'��/(��m�=�pQٚ�_����a�=�q��r��U��G���'C��e���ZA�	m��2�f8��J֋�5�H�|*�`����%��NZ���^�ț�j��}�nXC�6��&&�)r��_�p��k�$}֦��m<��&�0� -���}R�9|hE^���Wf|#ϋ6��:2��^�+ȣ�Z%�����,�j��p2L��#�E�S?�P�[� 'q�-����e[,�*a�.{cЈ&�MD��o�N����#z�^W�e��oA�o�*�G|0�{�m"�\
�z:�K���g��=C>��@B�W�s0[o��/�]T����6��|��#�f����70�p�®.�S~f�&�g��9�����i�7�F�ٻ�\Ҝ�n�+��H��)���_�V���x[T�R��8�۩�/��!������(��]�.G�Y����:<@l��y�+"�p�����TC��������K���Y�!��8�(�UmV�*g���1wO�T�}�6�㲍�?3Z���I�3�x��޷y,B�V_���2��N�Eb�Z��D Cտz��"����U����2쿣)�J���pX1Ҥ���q�� 3ƻ^�_W���enZ�=T@��,1,��w���<EG<C T��8¼.'�v�#��`�KeO����,*sd�D���ȩod���Ph��M#�UZ���֨��\�����#�������랍z��5�?�̮9oi%k��Zc����\1��H���uζ�g帺9
�
�M2Px�:��8��yj�h��[4��I���_ �-��0yHyK3X��X���2�?؁&��	�GOO��L=��6������Ө����������7!��h��WJ �1�ŧ�)�z<ǘ�.U}N7T�}�@s�m�	���NP��QV���\����nե��(�V�C�n�钸�z��3���O��2A�U�S�Bu`��D�|�Y`�Y�t��b����ۇ&�Eh8s�8pI�\�p�&v�J�<���Q�Ϧ�h��.lJ�b�"�����&}��M�^�|a�;%��2������Uv��T"̋3,	�0�%|]^�����	�{Fu����s����V2����(���f�V),���Y�n�͢�G>3,�J�T&f�!8k�lrV'��[��D��A���{���Τ�j��˘�O�C$v�S��m��2�`h���Dv�n#z�H�.��8p<��¡rO*�O�6�.��3��|�K����<1T�d�� M��b2%���l'�kd@x$S��8�W���(��#��,*���P��;�}���;���m�/�m�!,(UH4���X�(��,َ�B�X�����v��Q:���$�=b�l�W�cs͗�A�)x�ol���:�}x��aU��i7Jcv�v��L���/5xޠ���?�a���@=9(����.X*O�!����ɝK? )��q�v�o�Jt�I��u(z ��!�'v��&�	����x`����2c��c;��9:�z��3տN�_t���?7��6ك_��.+��2�D�@E��6�~�ۂ��EQ��uA# o�\P$1'-?����H|I���#&��|�w(��.9vM���.*M��>%Qmq���>4�M?Y�1x�S�̕��VMB��k���(����(��A�k9�|In����D{(Us꾥t�� r ]��Ya é&��> ń��1*e��au$b�&����(W�Q�`ɐ;!���j]��T�Ѻ��Z�����n�x⡐rԥ_�ʈBD��|�a��d=��*�W<o�?~��=^�7�0D��+W����b�~�(PAY��:U����oo�u�Dn�K7DpW[O)QH�Z����5�N�\���.�<]�����%����[���<v���HYpR�Ě�v�M<9H�Ԩ��˗(�J�$>�2��{PQ����|4ld6�2;�'����AِA��^�NA^�QD�_,O>��s�o-Ѓfj��`�Nw^�:G�yK(/�#t6LPAEz+��7T:�D�V\��$�	d�ڒ���#�o**�p煿�x-�i�m�fyg��w��k���U9\��6idh��3�/��Ib'���� b���d� ��f�{�I	�E���K��j1I�~����,�n��E�;�����a0'�;lq�;��EЈt��zy͕[����c��x���)��;���=ۯԥ� ���,�[��w�qIʽ�3��\
�KPm�H5m��?CF��_��0K2Q��
�#8��Ta������Z��-: G��5�N��Y��Ic)��7M�y��)�˧��.�n�F��LX�l$�+�[-�F^:z��!�o�7���(iS3�L:ޝ���:��z�l��X��	q���G�#�sHީ\$�A�}�����6G�x�����1A�џz/�lB@��  �d�.��<���Z����w*Hb��w[_q?�K��of<�?�8w�`��n���Υ����K��������
�<�c� #�B4(�ZT�M����u�x��n���h}2��{��M��B���3�]���R��V>����OC��}���ʓ�K6���O�
cH5s�~��-�s)9b����W\&0B'#��w��ύc�Ž��>��$�2�����^�)(f��E�P`a8\�ל����!���L�K��I|Iж�A�˧�Ԫ������ʆ�^�z�p�tv� ��+��vW��;��ö��wg��D~Vh�8���b
�i��)@W�Nl�LK�QK3��WU���,��Ks������R������B�dK�)r���O�8��J����v�s��v� S��ӧ�P]�ϔo�����3eP
0><IbV�%o���p�>k��hC�$��6a_�"t�{��
��G�+��%v�1��� ��ZNG!�(��
�A��	z]X�J�L��^���K�	�+�b��ɲ���{
���ϸ�@6؆��ii¤	!7.l}ˈ{�[��@���uv���'W������XQ�7���2Z��4�v&��A��)�\�W3r�6�=��iю�0ѣ6�:�s"e��A����	;&F�Pd+?�H%5?��"��F)�8��@W�<�~H\h+�2�*�EkUMeS�q����g�<~<�-� �k��A�q6B�@&�$��jCNp� ��+?��JRڐ�Ŕ�2 F�1�/H�"ո�EYC��dPk��p��G=N.O�$L\
\l(	�[h#�P�
�Ou���%�{
j�����J]6�d��~���7s&��]�}�ՠJ����������9@ܩ���H2�V�������O+>����f3@8�Y���������Ѽ��]�tɤ����Qb�Z�V��խzP�Y�c�v����h�Dud]W1+�^�朄�/��lf�7���<H����zT�-��~ ڂy[7��)������'i
.	_���乃�Y0Q'�j%��_�S���8�e�8IoF�d	߁@~�,,\	4�4���G
�%�>�.b$�&b��+k�dD��h��wye0�NotT�@��S�$<e�����
T͎Jl2���k�
�	�u!�=6�K[W��^�w�s��_� *���[õ �f\�)���6[�P˸�׳�QLjs����#E�-q�P����?������)�(�46��b*B�Q��*��9�H6|r1�[�H���n�=�+����ʪʝ�g���5�^�,�b�|-M�|�յkg�KV%Q ]p:�� B̺j׽����i��ƨ����h�.��E�&��j��w����:1�G�LA�X���̬�$h��0F4�Yy��%n8�Hc�����}sԎ&t�,����"qV��L�3��wb�iT� )o���`��R}vZ��@�VY\"�~�|k�;:�X�1����r�R�����G�L$D��U8#�6�co���H�uR�匆Z�uHa���>����5u���c�
�����>�L�x.R訑����\�Q!�)h9_m�7�!e5I���uM?Z��,x�fK\��n�n:[;P�/��i.�{R\���..$�i/ei��V�_���PK�Aڽ���J�o9r�ڼ��U\E9��2�߻P���-� �2 7oI�h�U��2i"�+ :�+:}��o���0�v{�:�҃JV���s�FKӋK2'1g�'���l�N�V�o~��u׶(�o�֘����BH���h�t`#G�˅�N2ȉ"7�q3��v��4[���}>�	�$�Gws/J�r�v^�b���V����A�����Y o�`
�%�5O�D��Z�]���&/��.P�3�CE��A���R�%<�	��������8)˦ �����B��S~L
i,�Rk�$���#ۋ\��"�7�8�M)m+ zG r���9k6�0
!kj�J]ś���.z4�"�� �,
�hk
�-g�3���u��8�E-y�
<�>oǍqg���������s�+}�G�N�a��"���;����Xl9v�������<��	:%�� ��8��jt\v�V�@Z�D4
r��J�#��1���]rn�R �q����lH�/��X��<��+�Os�QD���W��Ny��E(�������Ⱥ��~���Ŷ��GG3ἿU)��xأl֑��F�|��"�\;֦����=���	2�EɈ������U�Mw>V����h��_�s�g�#����� �3��C���[�^(#�q��p�B@Wu9�?֛^=b��x�B�sJ��߰ʼJ5��/j����C0@�I�4�P��I�0yb��~$�AS4�5�;���<wGm쇅sD�&[D�n�Mi���$�z������ڕk���n_[���f��&X�ˡt%C6�	Yi�GCY�ä�����V�$P}�Epg|�a��i3�*�pl��,_N���/Y�g�� ��d$'1L�YI���+i#f�� ��8�`������(?�(���#����/�:�VbfY��+U`�G��qg���EF�<c�x�0b�8w$��7�ȃ8F]B���ޝB�1�k���x�w�I],7`���e@�b�����6�������]�U��r���X�|/��6�h�Fb.�5�w����%g��Z�H���X���+&s��K�;����H^��k���M#��+�O��#aV�;	�B���lT�)�:�����q+|t���b8Fd@�T��W*�b@���Ք [?V������6��Y�2��¾�ث��sw�z��aȆP}�Pa:����X.�;g�E���2�T��Aʉu�Y8�Rv��g��1<�s.��C<��aMX䑰�����T��hYJI���٧j��z*�T�-A6��5�Ͻ��� *�n�ŵ��9�m)����1��V�b����iT}תiR�͟���[EYށl�}{�1��P��v�a��	���jN��ڄ��<|<�>oj�Q�CS�c��ЍI��/��F���ʇ ���^V5�o֡8��f~�}7K�?�� �X.�et����s�o��ݿ�_�O����n #ޑM��׈8�r  �����i�D������5C1W�@[�����L�hIE�ڇ0).���4-��'���/bS�1��NfK����"lH�1 :����%�mMHg_���Sv;�zL��KF9�V�X�jcCQ�(Wu��Vtͦ�A]N�$��E��e�)� ނ���t�E�t�Mƾ�� eB��W�.�!S���98��ū}��!cF�{̅T��þ��秖�_d��31��!�f�!��;���(��Y\!Ƹ�'�%1CC��r�֥VO�B�[~fK�9V$R�DU�5����tQ�G+�ʯ�k���3���r�}VҜ-.���'��B�vD%0 ��O��/r��(�_)a-W�jϫ�5�e(��:ō��<�%ۧ�c�51��G 緩���ا���˦��?�Bgf�B��<��D'�r vG#`[`�7���J���ˏK��;aL�Ђ�������J���H1�9���X6��8��w\�U�S��ߡ䗞��e���Ż �<P�tS�(�ZN�ᴣ\��l�=���e  2��\Bޡ��-�mkR1Qe��C�lg98 \4�mȥ���5�J.�L��v�w�A�-�W�gC='��X��[�y�1�r T�ҷh��$��#I�� j2�t�P`��_I^xX�c5AV?M8�ԡ�`���ź�~v�B���� �{�!���햹�������bm�8�~_|��fG��Q9
�ߘ�Y�+$������I�T���W)Z�p`���z4b����o�8�	X�φ@�5|�g���J�gD�w��d��km���w_�XR|Bx���J*H|DHx����)��՛�4�q΍Md��P� a�Z-���?g���>��S�Sf�>ӊ��WR㬪�
��v�^�[)�#����
��^��'d�b����h�]�������q�y�i�V����Z)"��
��b"��~���Q8�U˿R������Ǡ��\�*/ח(�/�.N�����ߍ`X��&2�g��N��1p�J�k��>�cq��@mRw�f�7�95ٞ��G��a�?������g�%��������~���O�n�2�L���}IaC�!�\W.>G����2��c?
����~��S�:U):|�}Y���U��cO���k�W�Gk?�~*����B[����ZO���dn�X�:hd$�Hr�w�O͛�=��vE���cp���k����O\����`�nh�x��n�Ic;j�t��	)y@O��>�&��_�@�05�6*O&?⧫�X�6{�-�dQ��rJ�ۏ�p����J����.�����܀�p����\�\
G
�N��?}Z�8�^��w�0����A��'̶�h)���%�ND?�+� ���$'Ge�)����I�����$˗M����׍�-
�t?�{���FK�y�!��br}�9x́�G�W��;����p������毢DRK
^���Icq���v�4H���bX�Kޭ��{��O1�aCj<)��p� {�[߮�]�TA�ġ	��n��j�Dm�کefH�$Y��3�ʝ��t�2�*�����T���]w^�s�E'+M;��+g:����w��s���Z�(}{����l �G^�M.'Ԛ�2��ó�d�j4�0��`�f�Л	�!%���.z���	���;�B?�7
�Y� ����<1��T�b�(W4�
�x_���&��rT�aGbL�>�|����)
+p���+����C��`��-� ؼ����H�������In���C���2���<�G�5˺g��%�k���>�1��]�I�nQcc���ב�^����&)%��y� i:�}��6�c+e]�>�R͑¸g�Wq��F��ʜj�䴜.��c�t�b;�0m!l�β�v�N��������M$dO�UBͯ#��5��{�H��F���n���Nw��{�&'ϐEV�y|d��;+��PYB&7�AM�� ����-`o-5�'vI��M�%�|�5i�s;����$��)l3��=R>�r ZӘ3<����*q����@��1�Y�(xe'J5���J�}�oi'����^�[a�AԤ�{�9�77$+��p�!�ʳ>E[N��>Q)���Ϳ������Ug2K��F[��=�%L�Y��²�K)u���=xKD]<f�!��x��ՍN3	պj.9��вawx6Jd��d�հq���W�9�w�����_..y,gg�z�87b�aC�x3���>3 ��+�*e&H��m����ݩ�2	́\6��|���lB��ߣm����� ��	?�|rt�r�r��_�LF�'zx�Ƌ�F`�5�^X����d�r3rL*(@j.�W�4�
���쭋G�S$���1�A!���қpӳJ_�f�q�KN~����kG��q�M8��j��ڜQ��
v��_��,q��O�ox|�K����\�}����d�9��`�T�+@�o��D}Sj]?���
�T�k#LaSiv@��T��X`�0�5+�[n��ٌF����B�m�}��T:���l��Dvp��v6Cb��|[D�9tïQ*σI��As@��q�`	�&k2�N�BR7źmݷ��<��3�$����xݮj���)Y߀3b^(�az���;�~����;) �9��2ϙ�a�<R:-����"�QK�s0�7S��.X��w��xUg/qd�ML�|��VwV�p�>�;t�����r�j��s��tX F8)?c_�/�$�֊y�~�-�H�L���t&Y}�+�M�4��������A����"�	r�����'�r�F�s�#!kڏhd*4I.ƃ�g��nK�J#9���#�v�
� �@P�)g�:��+�(��0d������+��dxݢ�JF���Y)�D���G�AC��|\3/�pZ!�K�KP�G胫�[��q��i���j�Dm=~G*�k�����;���f��9��S[��[X�{����Yx��M�^>՘�9�{�p��-z���mw�	�'�B��T_�/F�Z�J[)����sB�EܹL
J����5;.�������4��n[�=pH�����k�ec�,�(w����z�i�(�^��ۻtp]��X:h�A�]3+r�tx�����_c�d��g4	�|���ՋF�[��q�8���?�f� t\U���4P����qؐ���S �Ǔ��aL<s�{ ���}���cK�%���c�^[�8DiaaR�B� �,���d�g��k���� ,T���<}�#O��E��)�1��,�*8��*�1��SƢ��C�l��Z�6��u��`^�$�-��G�h�S���<�/%��j��b�C�u�*QT_�(b	�y��7c$]��"euO�.2�9�H�d��T��`�Z7�0W��l�Ԩ�J(pe�F4�,uD-��`�z}�����!�\��1^��b����==
.�?}t��7quM6�g4u��Ȏ$�@��e�f�D��''�[@x�������.�b؍�;?O+�NB_L�{6Lv���i��Ꮩa'���JD%�s}�8��iB;5a�P���*E�B���r����s���,0��E�*ǖ�+W)��B����.Rp���
�K?�{�������>*�m���BF�5B�tr	��kn�	�w�ݎ^P�%�\��V��P9k�����Ja]�9M���ZYǪ�v��#��-����0��?�r��Z gn����"{a���E���!l\���ݦ1��7� �i���<0�o<'c��%�/��%��~bZ��|���j��C�~ʸ}�����N���m!�3��^��sm�GE�q�Zy����׻š���gmg��5��zRi"���l������1���8"�Z�$	%��&�u.eL�R�h᧖�m�A�~�2ʹ�YJer_z��|�r��JVyJ�T\4�A�8^�V/F�I�Mz0G]�D��X�����f ŅU�8P�9���f=��.�<�<A��Հ�R�hX�Q�i�0AweO��a����]pʭ4�C���V������TeFޫ�������Q��7͛B����3�s�S#pVN���LQ�-y#K��@Z�Oȫ���˘=7#m��+����'P��� �'�����z��y��F_P���-ΐ�yg���Hi���?��떐n\l�`n}l� �
�qƫ���][�U�G:Mc#��?e��t/^! yQ����<X��P�%���}O�����#���gw�sf F��xrg������-=D�im�": `v+Um����~���u������Ҿ[DR���Ɉ��,�5K��יwl���X���a�Um�fC������0�J�5�yο�c�*�����u�ƂD�z��՞����;�vq��8煚3'��ݩ����jlܲ�q����eXO�BzQ\
��
�d;��tP�N�� �>fxf�s�0�p/�@K���Կj>S ���O9F�4l�u���8t�;��P�T�Ъ��v]�G��_.�,�J�SE5�N0$�
q�G�	p�l��AU�	B
%�J��A�nG�^�YDR��_o�I�pQI�VV�b�Ӷ@/���F;���BЊ�� Ƨ-Q�^'�AzB6�lS!�)qB���	�Be�56V��"0ʃ��ᝠT��4INiJy��a����x���CZ�i�&�s�=f�"A��@�z[��ĢZ.}
�A�@��-w,f�r\z؛t�\�����Ԉ�W!�k-���]P4(3(��� 0���>�����]f���}��CS�.���v��Z���PU�����(�X��і���~m��(F�؝��i���sl�҃�-|^�=WL���g؀s�ȟb-�[˔���/.�f�(�ta�fN3�"�X��~�+o�S�!f��{��K�h�g� ~*!vv���t�xB�r ��O����hH(2W�j�q����1��������� ���������W�ب,m���9�pH�Cl����x���g��|p�p���-N�v��]G�e���UyɅT�Q�7Qbp�T�Pj5���7�%Bq�c9ԧ���¯����Q⑒���?٥Ԥ�	����wED�̃:[����J�CV�yʠ�|�{}O2VM����$���%�� �+����&�F��Fv\C�:w(�J�A5����^��br�1xיG���X=F��$����R�G��*Iy�
]6˯%Y�S�,�9�U��q|�RA��!-m�9~�2��<��H:�*E�dOl�+��0ʅx��ÿ���X��&|�&7�nx6K"�}�vAL �7+�(���1��?U�̇j8�HV/�[�ߑC�.B|V��9U�WT7���ILlO�f����-i*ğW_J��HL����Ƨ�� ��c��n¢5LJ�Q���<����s��k��yӨ��Z�7Ac@�0�
1��s��O�^�W��nU(눅~��^�+0��I��"�Cҿ �w�2i!( ����(�q?���6�(�[�ܹ2����e`Q<����4���U���au�������7Ѝ��c#�s�?`��""`2���F�^T$�Ud��(<lj�J<n�>�Qq� �R�,Mz*U��()�U����"��Md���]In\T�.-94ן��@���.����1SM�:���a�1*=������F�BQ+X�:`¿�1Z V���^5�t��O>,&?Ad�[@%�g��jT��Z'�=ʧ�&��,v
��	�*N/z�I���`\-AV�*�,�E�����h\;����.��O�4�Y��Py+���T��Xm�B���c,tO����9^���!�&�ݻ�V��3l���N�ٌ��^A���Ic>�P�����)��(���B_�;@iO���ٯ*v$\uKV�r��'p��2]a*U���U[}+�����f��umgt���t��ż���������4bV�'�1��B.�8�Q(8�#�Z-"�*MXJ�{E�Ek"Xӊx;��닗�m�s�N��m��	�m��L�.�q	�F����<D����%����*��(��7��*T���	�ױ�o�bUs�� GH��.��ReY ��(�b��v��ˑ�f���H�0�{̐��G��_�e��H��!���]��_�6��N�����/�Y�M~+���RC�Ԝ�hd:3���0X�y���L00���I%���9�(�����N��a�[Ѓ��ڥ�kf�#,2c�K�qvݠ�e�5`�d(�k��s��������Ȥd�����T�9���P��O7����@�{J��WWQq���/c8IfG�𥉉B�V���#�L1O׻��q�s ��Q�u7��%H�#��|��v��׭G�e5���B٤!�)n�s��}]��ӛ-�3B}š�m`c��;�1����~:긛�;�R~����f�;��>W����ҽ ��V0�=�Ơ�������I������_I��Y������}��ud�����Z��d_���!&
��m�� ��X��5�<�u!f�G�N�G%8��������]Wu60[�k9�l~�_��@j����خe)���GW�JO��ON�>3�3d $??�����V�U�aW.Z�F�t�G�/��Yj��!�s�� Ni�+_+��\>����.@P6A��PTq�Z{�X��l��z5j�fA,����0���Xfi�/G����t+��+�-�H������F�mV�h����y�gU��%^�?���G��h�A\pA����.�A���C-�\���COH,B���s�`8�u�:#�GHo$8zS�:H�^B��G��v�8b; d~�K���va�I]��[p�\1�+*]������uz������xU��KL�ڋj{�*U�TFVU��@���8���ng����}�s^�*�6w���)3$?(H&yD=�ª�gm����R�êg^6,sd�TK��n����N!��EtD���Z��KX�s���'&.���F�Q���:Q�-߬��{�	Zs��ٌߴ��C�`X�E��-����j� zy�6
�Z�A?<�TXϫ��D�*Z�d����]�$�B��[)U`-��:��2һK�X(������/]v1%`�;���h��}��'d\�d.v<���mǧ����)�a�p�94�u�3�l�β���2����6$T�6)��ވi4W:#J���S����vEϚ�b����,l�vh��b�}�K4�\�Ƽ뎓W&"�0P�䨘��V ���r,�q���O�Ix1E�7�(��c^Dȷ�����9'@4,1��c��@��1<e	ey�D�_�!<D�LJn�������۸��矷6����& 8���.vEV�`i�^!�C�g��Ǌ��\�x��4�;2WI�߁rJ4�NR}A�T�f�LZ�
�|�r+�A뼔�0B�LJ4��~�i�4�~?7�"(v��F��b���}j֢����f��i�v1���a1���/�F����8����
 ����Z eE���,��9lέ^��]����� #�[��8Lܨ��� j��n^F�$�v�&�4�#�Р��ew�-@���PM�>O%�=��5������Uy�f�'��H�-�іM�b��8�`����I��@���T#��+^�=G�#��HJ�$`�3�O�.^J-��������(�|�I��,�@F~X��E�I|V~���<�`9K<�Z�E�Pʗ8m$�j`�~N}�g�;+h��b���Χ�w	ډa��q~�n�Ǎz�e�U�`zC~��J:�b�=�� \�fu�k�!�%״�u+�m^iʼb��ũtzi(��j�O���m�g%�� 2N��B����&$�ƂMp=��tjHQ�v�_�ܲ�������U$ڤ@4>�r��q��}��E�ÕQWѺ�rC걅_�~����8�I�x���zY�������pe�)rr'a����h^���p����#b�^>*�mZ]ʲ$3��e��R�����6&[���MWf��z�H�ǣ�`���r��J&dʿӽ�T�شk0|��L��m�,#�UqFh� �K���{"��e/kQ�����£���+;`�T�o����\�� "kT� ʪ�@F�����o/��8�����+�� %�e{�n"S���w�FPr��mP]�2!m~��I���1-yyH���/ ��VV�ԕ��e��F)�"Ab��h[�~����?�޲������[~Úrl�OG�t�>oko�����z`dS��@��;�\`�
�W�
�(������J�Հ���=b����.ײ�Yo1�O� Î���i�fC:���I�Pc�LC\�&�G0܇�	��䙡�^�{�r��r�n����f�3X(�1��e�s����u��ApY��_� x/�̛1t�8�F�r�3_˺r�W�U��m$��+�X�|���-�r,5G!�~d�%�"�g��}Un�vG�|'�;Z�Y3�7�ց}��tr�����"�nx�PMl� �X �#�M��V�<�T�7P�s⁆>#�/n�#K�-��3�N�)�x}F��hP�h������]�nz�\S}�H~��7�>&~I���h���۷!{l��l�4�-?��c%���f�<ƛ�k�����F�\�0o(�Ue	Z�%�H>�>�j�eH�cc#��y[�M���&�0��R�R������FR�1��
��k�y��R�N�7xl�:�&���޽v�Y<Ur��,U����o�����&D��n������������*�\��^�(V�P]��F��� ��4�;j�p�5�����ʮ38ksa"U�Z��0��.�_xUsK=�o��d7a:.���-�o�ix��[��i>eZ���gU��a�/�Z�k�p�*�V��M��%����+hy�5&��l2���%Y{Ƴ�b���q8}�%[��8ʗ@�����xBYo�Ԑ�ă�ߴ���OG ������0��:_�	�X5n��1�K�@��v0Ҝ�[��H}��XB���66�@Hl�ȏoX�?�������>H�9��*J�ߝ6�?0��\�3	0r��:oF%}��{�(Q�ϛ��r��JႝX\�
�먮�~!�Oy^d�'�p���>|M�N��}���m�-r1�2L�s�(�բ�Kw�®�T]�@�Ü�)D�oul�j�H�X=x���Z�g���?\�[sؤ6�4ɓ[+΂"(��Z����h �%݅�m8R{y^����5��í���x��	\^�Ď��R���ܛGOx�e������V7��	�O�DƯГ����G�w)��{C��g��ګ��J����bI�.+��wOkd��һ!�pi7#��֑d��W+V��A�c���錼.�GhB�����͖��~��bX7K�i�e~O8Zf
t���ޙ��'���S(��ӡA������	��~%�M��wEՏ��a)��C�B\R/�|�w�8�3j�9%F�O�( dO6Q��տ� ?l�'������k�X�-����u� �Ь��0|R���j��M$��������0��l)�QZx5����-z.��_c��֯5q ٮ��QR�j����aW��zGU*�`(�x]��CB�ϔkO�7�~�u)J�����ԙfq���z�]$ZpFT���Op��F�ɀ(o�ȋ�8r
F�`9d��x㶝�C�.��I7EE��a���c�b��R
»y�T"�YɅ�����Ȳp6u5�����N?���V�A�/4��~uҶ���Y0>�:���k@}�;��������xB$���BA.��&!�lkFɋ)�O�F��;��V���k*CL��0)�i�x3�*�x_#sPY_�su�kJk�����#r���i�kV%��fh���j���	x/��^ >��K��O�#R�7�^��SAu�Z7u�����QDؖ�n��,j��*���lu�߼O��O�+�1�_8����������b\����1�`l`?��f���h����oY�9|�&���M�㓡*��O����_��+/�7?\���E���*
'�Tf�g���鋀��N��w�R�QH��Ʉ���_N��m�kޙ���P#" R���0�S�F�5�L[Rfz�vm49!+�f}�jd�`y��A�%N1�1h
w��c���qd��d�=>���2�a,Ў�=��R5M�ܲ��whnV�\9��Dt?Ӱ�j�s����9��US8P"��G�(����(�V'‽�vCf>~�뭎���>����np��~a���Zp���W�
�~Ff��ך�C�R;��/����Y}]iqdr�ijey��qS���j�@5@�rrFɀi�ˮM���o�۳�W�rE-��������w/�]aB�#�41�J�S��+[��D���:/(��[�(Q>.6�[�|2絴���Xx& I�ҧ^S 9�+f�!�n �7D�����B����u
��v���q�`���_x��2xhŷ*=&�VKa>�W^��>�;��xo[&|bN��W�Së4[!���P���P�ǿ��s��V��d���*��͌�\����(��lL5/�mhu"��y��w����7/�nP����]���m�αǞ��v��P~�ũ O1"�DA�J3��!qTi�%���m�V]K��C,�j�sP�[���P��]|b��t�����~�j�k供>� ~��B�Da�̀o��oҧ�%����|�@�M������#1�C��(�A��f>���aH�s�:@��ҹ��`�� �`��=�K`��Q�� ��7x��K�Ov��o��F/`��>t�c�7lP��@".V�˄0��Ȣ��?֋mdlg��a{d�j'��H%���-��@xP9�JO��UrT�ͺ�^������E�mPE�xMߥ�&�B�� ���4L��/��X����h���V$�,��b�7���E�( ����؃Kd%�?o0T0x��oe�P{�;�?�z'���,�sc�Pq��~7,,K�G�ved��s��y��D��%�}����N�{�gX�����=��ƮEA�qp�|8����n.�a������
N(��Vk)*�/��J�G�Z�ʴ�ԃ��J����`ix�ɒ5t�M�+@�5;Ql�q�����W��r���" ��@e�y(�����ͅ^���d<$���Ο�S���q���\';g���ہ���P-|�&{F��X��iNo����q=թB�#AUY�R� *÷�M���۟��1�$.��\'�2���H�ۍ�թ�8�Ɂ��G1)��'�����U�3�_�1�ސ�}���|ʳ�^��c��f���6�lbm��M"3� ��X+��b�����ӥFR�r@5L���&%X�1�@>v���hb�|��>nդ/Հ�S�-���߉����1��F���\��_�ݶ�,hZ�k�h*�6'[0o�8�UPBL�kǩ����@���/`?��Im�4*CG��i�\�W�5�D��o�Å�!��m��ڶt�t5^c��1>1�3}Ӷa��og�d=��J1r�%�u^���!]�9���j���qC�@���M|!�N�"���%��z�as	����z.7H��Np���*�Yxbv擋�D��F�K+���m����bt�&�t��}�B�~T��wh�+����LU�b�[6s��	.3?(yl*����IU�q�	rè�����wߍ��YL�[T�AϹ9�5wN?V&�gN���!�a(��Лy��y����Ar���%���Kް�?��ʈaHzm��c;�M�*B�MP���rP��wz�ϵ��DP�C���M�ו� +	�#�ۅq�N�M���JiM���ˬ��
�  ��K�->�Ȗ�m���	=���D�7���YN���ix3�I�w���C�L6���~>{���8_�|�Т�!0�g�R �o���;3yX�#30a�o�$B�c� ����
�mqуf�3+Ç|0��b=_�b��]���_���y.H[93�B	��L�]4�mI�-0C ��tH
ojՔ�b�q='��4��U����7qQe$bwT������gG=@�����'z�@#o�=�&!����Jv�.� ?p �*O��5^�
se?�eȉ3P�1�U`/w'�)z2�����4{�����M_�Jc~�\FL�k�6�/��� 9-�aLFF)�/(��_�j��VD�O� 
MM#�d��;1����T7�t�?�*��H��Z�ekTN��n��z?��EܬX�O��W�w Ekn��-��;YZփa��uϻ���@�Mxa��S����f�\�{�Wͼ�|q�f� �@{�{�ˀUw�z�׈�*����Gi~j�?�9�E" '��6Ⱥ��y��nD��b��";rY��|pw��5{��)e{x��P��ְ����%�'�j��Qt�~r�^k�o�� V|��g�>����`��?�%O�0����"�mƨ��N-?����!Toρ�=pt7M�~a���b�o�������[�r��G�݄<���RҔ����n��B4�.�+�gpݮ�f*�A����B �5>�����q! O���S_���L��rf������Ç}��U�CI{�-Ϋ�������o{��眲%`P�9���(�1Ǡ��,6Xz]d��D|�,�O7���9�j�D1�p�r�&1����6==����8�Z[�-���dH��M�C��UQ	�m_¶�W�����P��ּJz/ 6�F��6�Q����d�����ITQP.���?�w��*�������gĥ��+��&露�b�J��%���m���䐥�\�F��K4]~�k����'$�f�(f�9��Ffx_�L�������i��|����õu�=d���+�m�0�,Ĺ��D��6������{�x7���v���c��4ǧ�Z@���B���l1m�0X�LŶw�f�� �db��R��Y"]r�h�)��Թj�pn�V��4g�8�v~��t�N������+D�3�s�ۘ��:�8�խ�Wa�����aέ�,h=da��h"fr�H�\i�|Ν7�~�� �	�2GX,�7I�����l�J#Vor��~�M⺵����/�Q͡C�
�x۹���)l��Y���,3�YH�u�j{�`W��wiA��hN���nD��u�p[�J��'[2X��=��F�Y�ƉS��`d��N�B_#���̗�Q���!U|N�*�G�i=��y�*�M+j�߻f3��˽0���6Pyid(3E��<%�;�p����-�W�&ʹ�jẘ�v ��d���N��}x��L��P����A�1��,�?�,�1��qm�>�ܥ8q̇u�,Xi'c�-����'����ϟ:�|��Y�OSk���ѷ� T	)�@���A|��l:L�ze��Y@6�0gY�"Ia�{�ޮB��׃�R26����Ƙ;O�8F�5h:� �=}���V�/3	Kd ��"������Rw�/_g����W.+��s�N�>��*S�:]\&�1\T)r*��2��'�v]lS&-��9&c������g��.Nh�9#��ٶ8��!�MWLxG�p ��"�>�})�Մ1�jOZ��Vi�ao�n٪6����f�^3����Гd�,@KaVo�.�~�6���ZX�b�����k]-:���h��\!ߍ&��,�^���F��)��޲ɖ`j�1M���u3�
��(�9��`�+Ňa��	�� G��|	��Y��.O�\$�t1�B�j.ڬ�a�6`�}%ם�	wf�!i�x*҄��A�dS5��p��Z`���B�ZH�|G�Qh�'�w�1�K�� [p��"$���Q�ީ��sD���ym���)��G�iH�.�J
�ɫz=!����ӿ꠶���F�>?���t��c��b�0\����ix�X8�o Ќ�������2�Te,Q�K�]`]�=��8 9�U�X��e��>vF�*.����'}���D]_4�:L�<p�T�Ky��/��v䋖��;6h�D��=�U�R �c"I�t�N��w�a�^��%��9C\��*�&��N��Zk�IX^S@>C�b_���҄&��k��Ox̥��$��3#g�:sU�S�:�B��$�m�"Y�s�:�]4	���X�E��C�hC\Wy�~��EӥE����	o�A�[�nK�0MG�� �����wr� *j��E�HS����*�V|0�%���գ��Ժ��m�I���r���f $)���9�$2r�J����J���s���Ծm�6�0�{v�6�0)?Dy�����Ol� �	��
�$�F^��N�����V.���]~\�2lz4��n��&���P!�<��l5���W1/z�ce�g�h��*�t*N<��3��|���5�ة��۟F��u/��(څp�Ѐ8������T�\c��i�垬�h�+�*#��+�\|��^��c1U�V�"�.O��3�H:�)�trҀ|���LzG�z�.�U(;0� ���Z
��N��rIPJ1���Li�^�xM�_�mko���������phe�#^�[�Q���[Hzͨg��+]6��=�`k���+&���aTi� +Q����cI�c�&�	�D�KT�0Z�3�3?Wn7����[xP;���-�b��
�I�N�7�y=_t
L�����e;�3S�u��c�ƥǪX�6�q��!�iaǾ�ѣAސfs��sx�,sӅ�q��a�[T�2W*5�	�"��0.�$)E��70m��T{W��/�X��g��d�^��^������p��"G�cMBe��>Q�<��r$�}BO��Pr�hn�h�����$h߾�%�$=ᶇ�_�͏�@el7Ӆ&�(�n|��AmWݸ��݅B�C��gP8�F�5���0F =��m`�h�=]����t�S}F���0I�~XTtf\?_�M�6�X���ݏ���g���DL:��pg�����-������p.�/`���Jf��X>�g���7�K�3�����&i�~�_���S���RπLm2Rl�`�.�!\�0������5������ȁg ���
bQ��I ��s��<�B�	c�x����ɚؗ�ފR�G6gW��|_�2nK����B[F
Ӓ�ixX�q��r�)�QvC�5�L�o*����g����`x熀|F�ꆇ���8�ᥙ)����O0�[l�<;�6��R�l�	P�KPw͟Uv�}�Т�0	��:���J��3�G�[FG��	τ�kP�ꈭ�E�X1�̔�;2P���C�N�Hڼy�C�g��S�_���3xܕ�`��m`�dv6�����Hј�n�>a��b��G� ��
��m`��N>zut���߮����QN+�/�^{	7I懁�c��{e��2P�s3F��[��!��B��[���Q"������9�}�5�գw�)%􉐸�*��������MsO���&y��D�{t�n��**>�T��!~�t����]�ď+�΁��̎T��N��O�z`k�m̨[\W��o�wR���G)��2�Q��i�N9�^_��2�e��q$���g ���-:J��B�����@�I	��Y��K�;�Z�9�����t�P3�l�K˺s�E�i�:R�ђ����-�f���J{X�@]�*��t]�\4���wY2�ꍢɸ�N����u��.��������~�d�^�Y���	r߮��q"apfx�ǈ�z�tL%4�T����.x*�����ե�<;Rx�~�:$$��2�#t�W�/�#p�6��FT��Lm���lK���N9�O#ǣ��Eku��k����n�j~4��c�1��@��i�D��%�Q�;g�0t��G5���P�Xt+.�d|A^^�a=�S��F����Z6��t���o�[�������zo��_l��v@;�1q�e��vZ�<�� 0�ۓ'�����E�2�c��3 ը��?�?´LC8�k3�S�7L%A`Y�&���Dy_�j���i�BKڿ?�.X!���ȚJ�˙���Է�];t�槕O�ם�*����䔂����YS��?��7r��--��^:�'K%Y��� A��`�Ű�~���w;�@*�I���x��[����)����E�j�w���yI��qr�Ρ+b�oY��h2��>�5O���Rv+c_#�)ê�\6�t���O���g�FU�R
$�땟�_�w"Q.F�^v�`y�f�٫�I��sij���z�f �LY�r�#���]BL�hJ`�>��]� 踬��f m���Ư �bĺ��ԤV^�a�!._J�1�6�aӢF�h���Gt㕟��;'�t��d"w��$�=�b楋ˑ1C�Z�7�ׂd\�Vcg�r���v{�Lpj,�:5����eT���h#7م��xf��6s9�xq[CN��0�KǇj���~�Zli)��ò$�L�W����hUS��n�u;QW��&����z>�t�6�c�N�Dq�k�t \��}Wk9�į�^a,��9��h���TQU0�����D��+:�
\��?�@�wB��\,�Hn��2߅��֝�o����oL1��Z�x@&o0c���BA	����\9?�$z��TQ[�A��j��'��s
���s�4��!��?	%u#�������m�ƫ#��d޴7������j�<��d"�^3�����Z�n��V������^�\���}u(�.#��:�M3���2<VMX��;�~����gT����i�M����X-jLn�j�xhDdEe���FQ���9�_(7�`yˁ�O��%Z����s�w%Ә�h�T�]+n��}"Ů,c?�5<��TH�ƖAD��[M���1�|�ꔖ���F+��Q�\	�,����M����Lg����c@�'�-i�֨}���)�e�Z��I "���(GT��!����+����0d5FGfm�+C9mZ����T���(g q6^�@�Q'ոK�m8�e��Z���覇,=�U�^G~�ȅ܇}��0\���J%��!�	>��Y�ޝd!�9��r�M48�<�:�J��M?�cU�Q	�DV��������T����^��"��ud��{�DU�}Z�N�^�,�����B뼑�� C���ķ�6�j5��V��	H��n����Ɖ	٨���,��zy5��#W����V����A�U�\m��w:9��Ms�Vާ��T�Rr{��`��oy��Y)�n~�,."�z:�I���$��u��������Y�9~�����gP���U���n@T�:����sW�_g��e�s>2�,�·r��؟�݆߫lOd��<�f�5F�8;�����6vX�N��P�,"䤏.�~LlW���u5�J����ȕ�`W<��-+���]�w����K�ު��.FM�+s*YTF��7��x<Ш���7y6����	�t�4$G�?�h'/�oҔ�<�U!���C�uy0�U]��&������g�|%J���C��
;:��چ~��.�7η�?��t�'`]��8�����qh�|��K���T=K��I�A��"'N_ԥ�_U���l��i+e��uz��
T
Ăx�5v�k[Xסn��ݮ&�6j)JL�F��M��+E�#�wh�K�z�ꍷ߭�F�v')�>4L�-e�Fh���̽<��ZK��߉�ʕKܯv�P��XLK���Ft����y)�.!��2�9��d9SiT�i�F���g1��A�#���'7���q��R��Q9��T��t-�q����_����4�ڡ�\�`}�w�U� �Q�{��%�ΣNao��~�&��ByҘ5K0��� ��Q<�tK9��<��}��4À�ݔ7����5,��rWm(�
U��]G��za'�BPc������'�u
yn��~�%	U|Gk=t%�Q˦�z�{�,PL0�ŏ;����$8�s��;@��N�L|Ze#}���,��y|h/V�)��8�p����_"��Hc|���ɱ/�W-����wR\��)%�Գ���;6]o{�����&�/k�|�\`G+�$�mG]��P=������MK���	�����NQ녕��)E?����a��r���EBƥ{w'� ���zuC�eߡ$��R![ק�� 5� ��y�f�������������B�N��S�6�c��4	�om�:�3�V_����14w�I����0kB���B�{p�9,׊U�ϔ���){Vn4/�H�<p��D��������'��0�*���'y��S|�U��K� �ĝ���giU��ί�0��{-����|5Yl���� ��Q'+1>J���z�&�ᔌ�S�l���,�0�r��u�=�6�,Hg5wb�t�������'�y�������Z$�����2d'�t����P��bqDy�Du��;�e��u!���G�s�u̔�a�F%TQ��
�\@����t3$l�f�.�ۦkĢ�4���d���:��RM}l_3�?��8�xQ�ª�ag:O�K �o�1���CdQ�M���3=b�ik���1�f�,�3ς�m��#���L�J(�Do`�^�nr8u�c?��|� �ϙ�k�^�j�]��}N�ڗ'1}6i��S���ai5kq/lQE�±��]4��s~!C���������鋄�ߕ�	�1`?�뤾�|@������a�.c�в\7��?;>�06C!9��!�u��k�i�A'l�ߩP�Bt[z͋�d�y���k��P+�7�c�b(91� �^��F8_{������W��_~� �I.��
�w����U���pgG���B�.uɗ��;.�	o\
Y:
	�A,d��Վ|̇��,`J ]N�u���=�c�#�L��
NV(Q�V|�s�����	�p���lU�<�\t
�VG�[,��>\@��t�f���_�)���Px������P�����G�]tX���ըl�$P0c�B�Tm���8�o3���q�&��N��{�ʵ�&�쬿�V�����@&{D��0��xymц)1F��x����e+@-�8��l�U��"�k_H�&����Hl�Ƅ���ԋe��(7����W'�[�A��_8��P��>��d1z�W��D�׳Wm����?�t83mP�`!*��;L]/v�a%�'��u�U�|:�2�0{ݐ�A��/_�Pٻ��fPg���Z���=k�d�u�9�-qǃڲ�����i[�Ǩ9L��8�J�}�I�нr����n�I�1���O���'�sS�H�v���o��>nq��p�!�7Y4�(Ct�)��_O�.��=��>�!��aW��(�,mzϠi��w��DQ]��-n���� )���ֺ-g��g'Z�ֵ��Ϫ��Qy���:"���@�w�9��
Ĩ�<��ѯѪ=�����y{j4���>%��Zk[��n�V��B:kH����ڱ�72j�_�sW��[�m#�/�u��u�;�z����'[�m�+M(c6KΡ��bMJ�H���d!�����Z�c�u�����z��\��~)�B�
{����,R?LKwuf��>׻��9��V/
��/~ ��cz��?��.�<���1��6�o����+/}V�B��S���D�50��%
K�6�}/����?T�H�O��ѩH�e����~:DRԈ(�z�8�`�����OҎr�K�},��g��y�5����00H���f���m6w��D�y���1����f�8\����y�X�y��s^L"�|��Q��,��~��L�XV�7_�;�9�s�Ei�rh�)��������;�]ة���,��NV���x����>�c�<ڕ��k�y�В9>׫Gґ��/�"���eAM��i��X�ҷM��橕���@���/ţ��>+G���w�8�i���ν��x��4	�U��ˢ�{�0�	�H,��fHc��ʙ�L���0�//b��	6dxK��������/7Kʌ[q�E���i��