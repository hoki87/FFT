��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�#&��#�<�����G��՛��A����_���E��{�o�j�-�wmy�#fnqąMu�=J�(��]�
h�٤����[��wHOWeG�# ��'Y��l�ݱ_@1 N迱L<���I� �9�F3�6'kn��[��cv`�Ǐ�՝kb�v��1�gE4���5(	�����,V6dd*�P����+J�z���!�!�i��b�:)���L��pp1��|>A�&�p��ᕙ�.��{�J}N�3p��ڱM�+�!�s�+��������Z�)���n���K�4�"fU��Õ�����W܃	�-���˟5�T����,貈���$��{݆qh̼gY��h8!!ֳ`L֪gD���_sz�TE6h�v�����f&���+��6�j��)�lA��0'��wb��K�b@�����P�LN��Rڠ��#�bL qlnc��̜�Fܿ�o�}���HC�t�?��ǫ�%��s�蜻���6ak3��%�XөMP���C�l��l@� s��W�96��[7���5d�����h0�+�<����T
䄇J����{~jQ!����W��Dpe�����̧�������t�Bm��V^��F5�xG�zt���M�S�{�Ll�AA���]>��]���gF������M��b�\Q�k��Z_������h��ͣ�a�T6�&g�a1H|W�<��p@E�HMNV4��%Yrg)���N4��r��g����W�6����rw�w��|^&0�ҧ�~b(u�'`A���vj��U�?OH��ӥ����|+[Z�A,{�&�>&Y��q~c���������2P�����)i��������ы�P��j�Q<<p�ӄr��EVde�X�J�S�mh���i�./�&�{@��KRVMn�
Gmc'�ʩ_��,�N�F�MJY�TZa�p'����L��2MRm%��S�x�\��P�]]�X���i��[	�ߖ�N�g�1�H@��!SiP���T���Ơm��	���K֢ٹ�V|C��H�c������1�dg6A?���^���;������wN��#:����F��֣�X�
>��Lq����8�K���ӿ=���mN�c�|�w��rgɲ�%��D/�U��iO5��*	}."�]}*�y��vd��X��p�u��-�����eԋ| ��k�{��l�i�X�-% /s��A/�o)V&r	Nhc%�e�. ���ֱ���>�QU �+�.$k��Fʛq��S���Zq��L�ok��N�|t�&!\���)j �K��M���:Ic���+;(� �Ұlf{��}N'�Ly�)����+ǔ׹R��]�h�#ʘ�x߯���	<VP�	�>�t%Xy�!l�Q���EX�)�o�Ż�y�,$��ѳ?���3;m���bU��0ϰ컩5� q��eaR��܀��b1����O'��Vp'd��C3&�J(�D� �U�j� �J����a�p�a��9k��z�+o� L��5)��L@9��b���]���������@��J% ���C��+��Š룐�1�A��}D�Z)���Q��U$Q,�[Kč&�>&�#�/`y�g_n;����e<�}�za�6Z��,�ص��l�s *}�Wn)���^I�2�0��?Aև��˲�n
 c_�� �r���a�QPH4��V��}�M��o@�;�4���~�mY�f��6ٷ�#�5#�z@T��;"��عw���V5����ߛ��$�)�f���-���Z���V��b:�<F��D,a��r�+�M�II�NUҦ�x���3�,]���Ap��_tNy�,�Աa7T䆃�:�O��p���b�BN/�pX�e#5Ţ�I!F{W��^TC��uΒ�����D[���&�nj��Im���Wo=�02�$R�G
�I9A�Ŀ�p�"փ���l�	s�P:�S̲ي���2�|�i�wƲʋ�o�>��.��ۀ��H��YO�����{Z�-��@�N�������j}�y�,�'Z���=���Ŗ�d��%�Gnm~F�@4"S��tl�]��'�i&���bv�<Iq�H!��X�W'<��I�8�ށ���`ƨ�����y��G}%g��-��y���:�ApQ����Q���"a1���}Al�c»�\Y��O��Ֆ`l��/�T@kI�g��tCF��ɰJ|���򡣏�S�7�#�'�B�K�
n� �v7�r-^?#����-5�u���_C�j����ߛ�oPܢ��������Cy�(=���J�`z���C��.1���=�GS��B���!V��?n�~�L:��cZǟdm����m��o:���qw�}2��mM@�k9��n�} ]�oW�yl��_�Z9|��P�K�jo�s�@�-/�9�:^��Y+��k뎠r��83�B�"��GIVKO�a�x�	d���)v�ܝ.���U���^�e�����u���$�V>
�W����U}=�ol-����=k�X�����o�C�͎��ڡG����fTxr���\��L�h�F��kB�OG'���a2��/�㽊��x�S�#�R�u]�1�G�a[���W�HQ:��Jے�3P��H�$f��w���p���B����R�_5wY���O�V��s<���&�}�����	Ǔ�l%�jMw.�_*�`�ʞ�[�hV�#�(樰1����F&V��A�Xk9�fςhS����O�粛���T���٫�%#mm<BЫit�t��0n�:��xkq�*��F�԰(�j>w����~g����M�.���8W��qȌ:�?�eP�-|-�c�Ð(�ց	�@j�&�v�,���f��#��d�Y��^| ���;���ʽ:;U��H`��`И(�5����7ʚ������C��Sx���=��F�t�>V�/A5���D�G��ۣ����;"�[w^@���ouI����m�������I���_�[ds9<(���h��(�:��0}ɿ�mve��b;m�t��G=�p�yŐÓ^8�,լ�d��W@٭���\�i1p!���B��b����j
i�N�mK�P����k [2� ;�8��ۦv�k۰3����E��KXqG �I��݆veƇ�o� ��,��7Zl#���B�/ �u��G��[֧���V�k���c�*���(d%o�_�Iގ�A4Z)\�����ԏ��*�/�d��G�p�`�yZI'y���xǣ�y�!)�'7��k^hP�:�;�oz�d�l0\N��4���ϕ��^[��k4�����%���=���E�:HFe~���0�!������<; 8�޵�M�\�ɰ������*UO�k���k���V]��F^_����)�WtOb�`��{�fۢ�pg��9;6��_A�*��AUhHy��\�ʰ���L���@*�ME!�+QI'޹+��,H�
��MW��vA/@�1��Y�\-A&���wc��$���`F(# �m�#�/#�׷]��&���(�SF�N�J��w��E��KR�i0���:��2H���j܅%J�ƕ_(6/�Y��kR�8�(5/�STYCֵ�k�	h5憶%�5�����G��A��)�&.�]���YI�H#�:C]`=3Ȥ���1���W���	��"�I�4� ��Zn��R�Y6���ovw��q�̣<�ܳ�8�:eU�������uG����-�Jg:��(���#���J�!A�f���u&O�;j2�z���m	e����\�_
6���Y^H���֙��S7�|��L���@�'�r��l���		�[
�$^�A��� w�Z��nń�@�>:ׯ� ��is"L�'�:������DbV�hMf�Nx�e�v�E�b->e}?�a�Q*!C�\)!������JR��j�zZ3\�En�0��)���q��P��7(���{n_�z���RI��R,��%��7��J�ٯ��c1L&]���@`S��X=�K��.L�0�[e=I^+- �N��m�� Z��x�K�f� ��*'����/:z&�1�ִ�TA�"�ᑩ��զ�c��=+~�i������s��� ~�pz�F8�W�W%�ti�����^D�E%�L=�Yig*꩷Q����X��{�)[������'�:�����)��I� D��|���5(���.�U&�����'���g��m`���!)� �@�Y��LҼg��1�檰���̵�Rg�²���R���o�-
U�I�|e{��c�������f�6[�����@��C/���2��F�V�GX/��Jn
��ffe���!D��s�,C�/;14��e�%�Δ�uZj��e�t
��v���a��.[ws��f���P�ɂ$O��sm�!'��7;`�af�s�)��4�ɣ+S���˃�O��7E �`��?��tl��t�b*��!�褘�:����l(%�xR�lp(��������x6%n��95��e�_��W�$Tő�&:�s�]*'[�k�2� F_}�	�`�ꎛ�g\�f��Y#�>��zU����������vy���3[��v��}�;r�#䋢<^˙�i!���<�*�G��'y��Km�q~yc�zS�-����d��ԂC�ק��!McpV\������5|;E���#_}k0�!���6��z[�C5+4��)w:����q'���G_�r��'x�Kb}��%V/��ʡQa��b�Q?h ��܂��2*�y���F��Ar��qK��ȿkŗ�>붥V�}�l�G�̕�@[TƵ�l&܊��@Ot�y������ӷ�Rض�G���E���5	J�(��i"����'j|�E�jjD�~0~^ȯ�%i��/���g������lM��&��b�RۖSp��9bߜ������*�|�}��+�\k�yˍ����`2aO��j�����2��4w�����j��OY��A�Z�E�)I�`�X%�k9���;�m�v]����8b�5�(oP�ۀY�r�:VSq�5�U�7��R�5=_�������K=K�dv�a�شe51�af,l!O[�3p���������2���I1V����7�"�O~��F��j�Z.w��gs�3���z� Q1j=�Z Qh�k�G�ҙ�`�p�^�;j�cwHp�����k��JD�m14��C�o��ii�iг�W�H^������u\��W�Ru�[�w��k��J��s�|n�ye�֍���XhJR�W�C���Ǩ�,���X���-_x6��7h.��8z!�o����.����f�G�
��S'i!���ߎx]�~�c�X�\,���̶�" s0j^�����E�Մ�9�[[_���I_],�x�
�Q���v+��	yj�rp�/�8����,w�縘�6�d>u�śY���������%�a294��<��?� "��~� ��U$K���3U�20˒�&'�q��Ӏ�؟&J�]��Ei��n.�E���N2 ��1�/�Y���i���Z.Nę�*'0p���uÙ���X.C]��jk~��uku<�67b��!���W�n��X��FM��l䷃#��_��Аg�?��!>;M;?���QN�k%i{ �K����iz�j���z�4�&e�dA7�X����mT�|]`D	�� �3c������Rh�q�~ x��=�pM�]��'yM�4%m+� ���^��!�W�n�\G;hG�Id�YP�c�5�nXDv��Ik��b����:�����V�KU�7f!�l\�}lѵ�7c��6?��p�OD�l�O��RdG}��a՞�ZZ�:�җ���i-���o~��V�w�|����P-��$t�j��$|6�^Ǎ��Y�=U�J���qO!zy=�pu�]��\#i�������	�M��8��!�n8�>����XI�POJa!,��~���W-���a7����VL �:Y�*p2ຠwd8��Z��C6�V?�l���A.��Z�!r��;_W,��-5�щ��!�NB��-.�0�Y
&��v*���?�<*�^zx�}�����%�$���l�(A�_̄�)l�y�%�VN��xr�I�󦡔Hs� ��5v����,�rRX��#8��\��R_g*`x��>��u�p����t<�avKw����>����X@Ro0R,#֜*-���Y�u{�Z�{�T��Na�+��+�1���Y�B����.��}+}:ɼ��f6Q��{j�Q�=�5�$̫B巀͝GH��$�i�ófv�'u348yMT�Oj
e�^ŉ9T�-�J4r�� �M�b/�r;L��>�6ɐj��ϣS2�W��Un.Orm��Q�u�P/#v�'`��z�P|y�r{�ˬ�����R
Α"N"��.���
FL��\)<�wS@�%N�M񵅣���_�8!<�����in��˧��i��yR����W/b��Whr�C�����2�|�s�0f��Ml]ƶ������Au �i�Vp_{��yA��{z�&e/8��ŎRNx������*�TH��}�'u_��I���8f���d�R��|<�W&��d�r�t.0۽"�+wxC��
���]��U)(��aw ǀ���_E�}2gSP��P��� b��-��fh�w���@�g�H���-�I����u��BP�!�
���W��&_�d���	��R7�I����������y��
(��[�Ý2�7��|�^so��ݯ[��
L�|�#��y�VL쁍��y�#�sY�:��O��k�X��������-�ݽ��t��OO]���}��JQ�I�i˟)���=���^Ƈ+z������h��[^�&���5���+L�ӆ#M$�$�QL:!Ϻ7=\t���_�XO���N��
Aܭ�D,��ex�������6Potvy��HDG�^wK8�����o�gR���P~�\�5+��0CLm�? !8{��Ū4�<hg�R_�Ѝ�W|D�F���V?�.��2�9���ت�H���D���|d�A�Gu�&�3'H�{Ŗ|D"h�[;9t�-ne�2�\/�b��)�=�AZ�{��~�����pJ�U]Tvu���ъ�������J�e�|�Ou�຿m��eX�{f
���ٔ�?�)�Oj�����^�4�,�����;�H����p��Xxq=
��s����)�j[lX���,�;�Làwqt���&�7}e5�I?(Wv�|�n���w-h�kbm��l��sq�h��f�/��*W�������t�"&5l����A�'�H����xTQ�!�"��QX8U<GР��]=��,�lmQ�;��E�D��ھ��CG%՗3�.K9w��i�[ι��gݠ/����;�lc�<��-Ԅ^ᳯ���Z|��4D����W]�.��ㆋ��1�\i�R���!�G�J9BZ���r�
E�2A�Pha/�N���R��\c	��#-�����v8�ʖ��oG@=��p&�r��$�C�W�~q�r-.��0����'�u|w.K(��a�t&_��l�'��0N�����H>�8\Ç*8��[��;��=�����d�<���S�94�>J�aj� �Ղґ�wf�z��g�� �S�(Iqb5�e�VH��<5��8!�c!����!��-D?����_<ᥢo��lx
�6���O����ِK�,��_Q�ByfH�l6Fay�.��lr@��S@Y��-�q#�������p��t��DiY]*dH����i��0L�YUp���]Xd�<����Ծ}���"��8������i�kQ�RU���,�w��4����Zû�5�e�Bu-#�=�����~��θ�b:{HB���B���'2�v{��6��T��]��{ű�j`��+�Y�ɑ�?r��6y�--'T�y���-嵞�D�<\b��Aom�����]�]�S'�Z�4�m�5�@g��σB�S7)�Ĕ�`��Ӝ�B�UH�7�,����a�ug�q��%n�U�
DK+�k���>��$��X�*$�'�N]�"�����5M����^w���'��G�������u�N��(�A���i�IT��p`7������ rZ�h�y���c\lI|��T�0�[Μ�$o����䑩]�qQ�v, ��2��� �חY�#�X�o׆���	f�P&��Wj�sQc֣����\�W�V���O�&������")�pQ^7yA�욝�?V��¶�ك���v���|�~���]ŗzے=�;�Q�.~�	gB�Z�;h�"�,���O"��):�/B�E!� bѫ��!��t�2M��j��ˇD	�<�pl;]�,7�G>/��t�����<�n~������kdꨙ|������M�,���l����[	�tTe��� N,�i�@!r��?Dep�)ʞh:O���b��,A|��l��w#(���Z��^<\
׃Ul�i*B� ?��i���%[���6��\rl�{qPU�D-���'x�Ϛ�Z�[���NlC��m�����[��9�e�U<�L�0��`�l2��82o>�e��a�L(}�A�=�?�"��R���R)gS����3X���b���ϑ��2l��ZHi��gH�q��"�q�T}c�����S�?�Z\#�͗j�x�%�Q����X;,�2\`q�����7`����R�Jd*��gvǴ��<� ���P/f8���3�����a�O���'s�o�s��ڵ��VL,������� �-���0-ud7 �m �[N��^��e�<����f�K hVO!O��70�>��j�J�#�D�AEo����߅��g�n�HߙTnQ�~��ล2�]��O�Y*G�4枪)�[A�\6�1ǯI3�.%�f�10v�y2��+ʌ����}�@�b��G����Qⳮ-�R�y�	B�]�V�5W-QHi�h)����9OJ^#�a͛ ���l\��t:����w#�7�_yB�0 �o�vk��b6[�v)��h��ǩ�}Kᢇ��i���wȘ��������mf����Ƶ^.�5��
���R*�V���~��G�2O��䇾e]��4OedF1�s(�,�n��nu�ʽ��+�	a�R�����W�.,�0�LA~:6�|7|�	��=1����pJ)���A�H���Q�B���x�c81Rw&�%RD/������Z�?��4�����1��Gu�13�EH��"5�R��.�M��;�u�n�%k�`򢭧C��+�ב�4��^���pz���Ct�+֏NK������b��)�ԛK,�7�i��絉۞	��ٮn�ԑ���^|�U�*'�����3�S���йz&>?� �H��YM��*笘Т�?���c�-�_�;m�e�9����n,!C�B�-ٙ4�ώi��^�ˀ^ړ�}U!���l0�mi�a��@��r������cP�����[���m
����I�_K�1E�l�A�t�xY��Q��ֱ,2)މj��=�P+����jh��Y,\3�v��Hw�8X/�]�֒	JvE��h�=/���ru{�In��/�k�س;�:�Whөu��:�[�;��dB�P�[��?a8qk��E�������R
2���}����R	VQm�����d*�?InH�s�l�3l�#��4o	��i�ۿQ�ʶܒU�jJT�u2�ޛ��|K�X�\}���~Qz��^\F*��r�>����0'����!��Uq��)e,�~�`˄^�^[Z��S�Y���	Ofa�ޙ�x�5�v�Md�صE�v����!ߛ���ݠB>�5�F.^�aa곉"Ū2o&[_�u�;d#�6�9��l����f۔׍����꺪mfN��J;�Z�ʂ,pļ�U�q5S��p*����-փ���]���}�UBV�)�]�@w+g�/��zvJw���
�1�����ܨ��p�[ȎSd��ֹ���!,{�B���1��ܙ*�zs�X�Sk�����c�k=�$ƿ��k��!��;�_�1�.�x�s��`�/D;ð5�Z�*	�/J
F�l*ÄΥofw	���~�8��ӝ6~Y&��z��֕�j�tl7Ap����lFV��dH��}�@�Ä ��������4g�-�	��L2IG��e���ڬ�j�-"��`}�,f�����N]��.�S�ќnd�����~��5��wy؁�5�>�� ��bΉ�(yd��XN`t&�q���V�O�,S!D���f���LK�|�J@�8h�z�leM�M�O�����G[_�����`����0�pH��͇I�6�x�C��  Qϱҳ@ S��9��}��!ɛ�+O��� �ֿy	�jԆ������0ߋ�����)������{qnP�#9��ƀh��x�Y'܁�9��(!��t���B�e�BI���|��x�QoJ��)D�ȳ�iz� }js�nT�'C&�u�˿�o��4	�5�q���
�R =~e�7m�w�E������[���������[q́J|�h��<q�|jm��m����o����BҚ�3��{TeO	F69`0[��n3<i
�w�Ix�5�@����D���H���o��v�M�M��510j��#d���z�,V���k}��L����M
����a�͐sHޟ���<�	�k���i�<�v�1Y�޽R��}��wT�5n�T��b~����TU/*V"��39T1y�'��W�T>�L�u7�-u���3m��@���v���=l���<�m-#z���p;�݇�h�ۊ��pS���&��Qm�,@�;��H�t��V@��#r#	k�o��Ņ��<֟PJu�Y:��� 3I����I�{���G}0�5���|Gf�xt�߬}��z����*�]�U��(���6"�륭}k�<YS<�� �h�F��v8#���O�6{�.��	�l�l ��2J�<�ŵI�U1��B�K���Þͺ�O�/�����ͽ��j��i�*3�&��:���8i�=�#�����ť��Z+��3&cW�Ex�q�r���'*מ�!益��'l�M��^5$]���_���Z�E�=���6kt��q*�CF����s�*�� J��U���	��V��OL��C�YNv�-lP�����O*������i�ȏ�'��݌��zb'Հ?�+��k��)�!g'W׹/nB�TF�!�<�\��J�""QK'�E6d�N�/�ZP$�/,�~����?(%I@=��d��N��#H)��u����'� k�"�Q�ΤL��qF���Xp�V��<͗VĄ�r�U F�_%�ѻ�y=��X�qa8uTa/f�P��"��N��}�>_>%�����Z]芰���<t�RэK�iq+�2N\��s{��������"��ݑ��ٿA�H7�̎A	=�L�.1����?Oϐ��[�-��[(C��1FbP��PPrM�7�A[ ���Ow�Vl���)�&m�@j}D����6y���ڪ���g��nNӁTP���Q�DY��&�jXq�c6�:MI�>�'tx�8>g�u�R�P�ݸ�҉D��k@7�C�s�-�:p]p���5���FOlH����7��O\E����(�r=��~����}{M(��V�}:;t@:�Y��S�U]_�ҝ$�a0��c��m�p�O{�|-gu��ݲ/f+��>L�3K�jW'� �.�~N���	��|9XR޵�(_�����曪Ca㉔��ͭ^�F�VK+$]9�b,��u���w�f}�_�f]N����t?B������e�js���^ V��kt��\�V�B� C�������ۿPt���w�� K�����@�dW艳!��:2�oI�]�`��'I��J�p<KHY3�V)ɘC��i:�	gw�� 4�N���&�����CY����n�B� �x/֐�PA ��0�Y��lƹӡ��і�����sޒeW��Ŗ���UG�<h~a9ui�r3�Ƀ�*bPۺy��=ꍞ��q.���r�nF��@��"1��L���m>����>dR��<m�B�H챫[�M��Ã��ʎ�qciD4�r�/W�:�y�\��S|��|@��r0���*Mz��h�]<���SG�L���;:G�WSP6��e�N�^A��hE��S�^���}���a2e�B����.�0��O�����T�x2�S���@����Y����/<#y�)t�����V�yj��?�!�Q��.Ba�i��s%�
��a��`8?�?�{��p`���}<c���yh��"�������������"nҚd=�23���N^!K�o	U�<ߎ�*GI���2��\5�y��	�1��׳�����r4��02��
j�����
P�ن,6m-�nh��s����s�D�,���F7��7�=���Lޢ���YK�'
�ש(�0����#-�|��߳A��ƚӠ��6<^��JC��cbN'K]i? ��mGҔe����ZU��b#Pc��o��s����U��N����؞)4�6�����mʋ��d�ة!]!���+�6��LߑA�A�2��҉�6�ς>3�bb�s��V����ǑGŔ�9�s�{/Տ�=\��$>g|O-�@�c�cm�>DSq
�'@����ᦵ H��m�'��/
�5y9dmf����B]c�G��qs��K�3���f��l��cr�R����ir킙c,3���))���\�Q#���N B�h��#H;8�!銧�l
 'yQ�UFZ� �W'/tE�UJ�t��T���r֩T|3�fx�V �/N��6} ��R�dvt��,�
�+�S&����UUs��>$8��=q��_P��_�>,��;'���zGJ��G��g���S0�4�?)�VK��"01mE�l��q�������x�H��Cb&�7lVjs;4a�렖��	j�	�h��VK����xZ�߿����c�@��ނ�-
u�e(�eC�mڳ۹(�P�w�Jv+��"Y�8��6=��:@��7��j=`�ZD��<��v�^�ri=����w���\���@�1:�t!�u`�����6@�M޼�B?����'�#�ׅ����{^MEl4o�s��)�ۆ��Ԅb�G'���_��y¿\a�eT�{gA��7ҙ�R�R-�\���=�V`R��@�%���Gi����vw��GW�h���ӣ��D����~�r�c����=W�ɴ}��~nx��	�e�݆��	4ʹ�_��|�,j��JT"5<���&�x�{~wc���7m�-Y��V8IS�@�����Mc�c���
Y�-�-���:.�Y�,V+�@��'��R��/7xEK5�wd�d�/�7�w��s���T;s����C�KZh�l��kf�[I�ֿI���B��85� ��1��<g�{��(�T�AJ�ow�[EV���@P3(�g��a!mT�uy��ѧ��Cڦ/���@S��n�K����/T�f�����i��7L \���8�M�Ԟ|�~Ъ�ӌ���.��*�k��Vi�Z�?�-T{,�P�����1V�&����=W��ȝ�����~Ź�N�ǆ�,���/}2A�lWn�Hkn��նz)�c��q�~�v�u�td�k�:W�:�ʽ�<�[~��IB�ނ7���(�^���zZ�H�|PLA}�q(a�p���b�m)�����Ꞔ���9���Y�A�z?y���5c07��G��8a-*�G픜�eǨ��ು� ڴD$�zl��$�Q,�x������6���sS�2��oQrkL�9�o��]�J=^��a�¹��bہ���'�K��5�N9|�&��o�?�vu��`p	U�1���^r�F[��eܱHO��s��Mv��֌�iع�����)��Bw�_Oh�y���V	��kvR,^��5���ƾ��ءs��ε��} ��g�bZ���Z�N�����:9���tW�d~�6�;-���6��G9hM�����S�	��}�-� ެt(7s�Ӻ�/�1����*X��X��h�;{&����]��ѽ&���`�u�������b�����{�jPi,����� ���"���y�F������`�"�����;���b+��J�LÝd<�?*�R��QM���*ۃ���|��~LL,u�)�$�p��P�h`	g걌]�A}(r"T@�j@���F"�K�j�Ƭ�pu�)F����V�{���.�s �%@^Rj���$�\<):%��=~f ހ�6�d��f���m1 B�Y{�$�����k@9�#�ti���6g�R�u���Rb`ʃSMn��Z�����k�$�)G�d�4?�)7Ҝ죵�H ��
	������:�z-�+���2g�$�`����W�ˆ�L�0�Gغ�2�I��P^�*��/�4�w#��s0@��#8�'�SH*� ����cIb� ���X�C����	�I��v��p�Iap��z�"ix[I��6���^�%��h�w���נ�������Dhڧ��v�&�h��Ao��.�2�Z�s�h��U�i���������Nj�����xʀ2e׌K~$¼D�YY؄%�+G�J��m�ڀ�L
Y�y�9�p*�G�d
2袹�f~m�^j��k-?o��_�r��r����Hd�wqŲ��w�jP��H���#ml˯y�U�� ���
Gzg*r`�˜��j-���wo�Ȓ�%D�ţMb��Z���z�d�/g���n�������d�s��ۦI��X&\���PT��0!��_��d���E�d�W��� 0��3a�H|�`�L��yj�g��"�w#A&ͪ���1���Օ���5�(�՛k��~N��������m���d�*����g�|�y���!�W%���Mќ�F��	�ԑ֑-���d�W�{�#�����bb�����"^d
�/!��b!�Q_qi1���O�,�Ǩ�A�,��d�\߾��! ���l�b
�B�y�$����$ 7����B���6*g��^�D��&IBi�M�;�8D#�]���M,K/j�yt�Oza����.�v�F�րNJ�@a��>��%8���G)nݨg��6mi�	�z�0k��ë�o���;$�����\O�������+��ҏ�U�Sx"b�dj��u�~�f{t��ˀ5��4�d$@��]T��OOg��ݱ���/�.R��J&Y1GȈ(4�]�q�n��B$�(�=ǴjP���C����q�7yO�'�~r��!ץ#���ǹ�6������֖s�΋�k�z�ek��?�̓���&����`�cǽ��"�G�J	v�R�uTZͬ�?�;����u�,���٣p����M��ן�sF�I�'eR��5H���J�zN���J��}��ُ��*����ڙa�8�rH0�o�	y�$�4S3�����͢�Wy{r�֚���oTA�l�i4f�O��S:��4Am�+� �"2Fg`d�K�$G.Vc�]{&��X_&����Ί���7�yn�.�N���KLb���f�u���"��r����K��S�M�4��#�.��Rip>b�'�і2M,�|�����xuk<<�Gpاk����@(�p�L6���t�<h�����o;ꎣ�o�Df�5��q����N�E!1���:�o�x�\�m+��oeua�ɝ�W?㻿�z*����=��ڧ��'���՜)4���������S�R����5	uI�ڳ�$;�g/��>3�}�d되�yXC���y�v[�ӏ�C(6G3�V?���*����Iof���GݰM���<�C�Ԭ���WL������H����(��T�;1�+"E_1j��DT�:�X$���ĉ"�6yk�/�^֕}=�F�M�4�Ϻ%�rz8*Q{����ei���D�a��'���E 岣�F45��]�/�}��Zf@{@�-}^�� � �M��`�酱�_�8���i٨r��v��>-����������Pe��i��]V�e�P�а��[Ħ��B���'{\@4߷|S�Z;!o}V�	�	�5��ިt�)�*M���P*��Z�Sݛ�/3ը#�3݊�~4���.�t��g*^�%��p�Ӊ`2`<�ƛLP�����^����;n�c�ph>�gg"w;�pQ}���d������i��Ɨ�K�!�lf�����P6�\>3�3o�<c�C/�	p�Q�2���Ԑ���uD�����'��~Df+�6o�ZÑ�Q4K�U��>ht띏1MnG�f�^ �iu[��X_k�VI��'���"�JP��* LE�J�qxx��Q��5����p�u����P����iE�j,�I�<�s��?�G���,D$t���e�"�����-XtcrB5o��J��<9֎���6��8�:�C@�����yd�%�=6�^W8��>��8�8,�@xx[��.]3�J��g�vFt��G�|b��j��2��U-�����2��G:$.IN��Կ�)��Ni*����<���N�p�}r����ړ�^P顕 8�L����b��זpn����?�X?�>���.|�^�a� ��<2c��ń��IWj���pP�m��?��7�����L)������u�w +����&\�p�m��5�3�M�&�;ڱ/�f��"y�㑣�c�Um�b�'_7���l ���S���:����j!$��R_�{�d�cT����{���g�w%�:r�Y�En�*��j���k�j;��9���
�#lA��2F/���KH~�툀6� q�#�ykQ�a�Cyn}���c9���R�#��e��f]����N��4�� 7��Q�V��%�����cֿãu��cT�V�t��wr�k'v���8���h���OZT	My��xj�(/�R)RY��zSn=h7�xe�ڽ��[A��uc�q�����6�d�	�b�qADvF��O4�� �(~�������a�S������QC�,�Ijb�!-����km�۱��%{���%��Z`���7ױ]��<��ɝ��~J��G�a��N� ���ū�#V�����[�8��xM��I��@����[<�����3��0B�K� ���\ Q-u�uOJ�`9j��r���c%nz':����I����\��n�s嵎#�@����g��O]� �gݷm�$7�I�ft��^��a+1�3<�,��t�|jPo5�8IS�yiw��I�jY�ڃ��b�Y���n�K�h�@�&,�q��U""j7�UA��c�r��2�X�/�|�H{����j�]�l�5���~�
�p����m�O,Z�?�����L��(15�%WND����6�	ƹ"��w����#�~ �����L��]�<�J��H�ysu�l����.�R7rCY|S���\�6K��I-�%��}��&rw���2N�������SZ�%	��r��LE���P^!�����>�&�?>����8E����̆�O�u2�r���BL��:���m�������L}��=b���v�`	��@9ܛ�*���� �&a�
]�"�F�hv�E=�3��9p�œ�Ck�_���Q5n��S3Ew�����: �]���C���ܛ�.��_�%u�9���R��T��R��l	m�	��|؛4F� �H��X>��YXj>A-�{�p>��s��-�6�J5ί�?��_�J��3
>;V�=�����:$�O�҈��xQDH�ٻ�'��������z�ض�h�[����I�.�� �Tp�V�1��+yب�
�5 t4r�x�c �$�v��*��Cn6tg%K�E"�Q9����D��1-}!Z�P��c*r��.`C;m�s5�?��k?H��bc�=ͪ�/��W�|�Kq$�,&]O���{[���>x��V/YA�%hC��{���JH UuΈ�B͑�Y��W�W@2��$��~�Y:#=̧�W� =&���?����S]�lҫ���/&��Y�ؚ%�0�xl���A�������#9.M�j����{��������f2R@jvު|�H���zvI�}xQIhﶽ��4�.7U
��������|3�~=�CM%=�{��ilH�*��o��OD���Pg)�G��)JӨ���^ڹ��q�]�+q�fgjx����\�xU������k��M�ΰ	GV�C� �
�a$���_�aG_�E�PO��x�J���Bt��r���[�$��h��7���8�`v��˦�j�a�Tk�&�K*g��V�6WN�����Z� ��g��Gȅ�ՍW{m�d���hU��BML�L|�R��_6���جD)
��W�Q�>��#�l^�d0�'�&0�8�|�#,~��٦5���1z+�:���@�����=2�+X���6?� �����B?��c�?mV,�HFt�/�Ǹp�H�h��?r_vI#��D��G�R܀%Bi�{F�pʽ�e)�$�l��(��8?vG8�~tj�Wq� ��M0ej���^��i�)�0�>uP9o��ȼ'���!�qRZ`M�v���@�S����-oVeNİ�Ɍ��5��M���â|(�r���ѫu�i��d��׹2kҋص�r�-Z��`��d׋��.���s3�H�}z������"S�P�B}n#��g�&��xh�0�j���k/�_��Q87AT�́��֑�%,y2\�γo&px��x���Ƥ`X�����,^%��Ý������ĩ�|~�}�T���]H�g��,�f58)�#C��}@#P�Z�`�s��`���E�8?���x���N��j.w���Ҿ�5��*T4��`����L[L�1��j���p��!����/� �^p�����/#.{��*�����G
K��e��Zr�
���>�Z�k0Z���������e�k�g�e.'��)�w���W=�\~���<�~��� %�9P��v�g�M"W��oŇsp`"bEE:���4�%�Ghni�w����vLhZX>ٿ�+b�u.�؉>��Bl8=)��}��mA��^�0�l����ѱ`�;h�ÈH�D��c�޾��\�!���q� ���{&��L���������N���##�/���ή�-mEۺ�;��Ա�x�[ ������Q�b$��%Խ'�"�����`��ӡǍ;C�?���7�\յ��u<�T'�	c$��⑟� {�iyF�6��������p� 6���:'�a�� 7j���^�� �*�+Ȇ�o�yR��0 E��%�����0@���K�t0�e� 	��X�*E�·I�)"�l�w�UP3�wS}�f^�.ү�Y4�$�>�8<�Q��-�AJN�s5�-�s�tK4%: }�a���'s�VR
��t���,���P�d������Z�b�8{��ve�d�zGt�E�L�9�{.��Wk��3�X&.�i�Y��z�k�MI�Ҫ̉��S��x��с�+~j�qz4A<ݍk(�8�[E]����B+�~�S��ø�{} ���W��q����ќ��� ,G�e�<�C�m/zƶJt!��#z��s_����%�K�f���09_�W���F��aګ\���vT|E $o����dtC������	�y�" �w�xG��և��� ��Fj�rJC��h���"�o"�Մ@:-�V]��M��ּ�Co��]��������ŗSE�je�bc�&��7 wv7gPQ���(��܀��t���x����o�8�M�'�C��xO,Y̭��5%iC�V�,4�1�,p���`��B \�n�z�,iʒJǃi���EVm%���<�KW�o-�LN�/��?hWz��\^W���p�"���p� 7�r��^���l-�6<�*c������'��T��Qҥvs���h��� ^��n�p��*5��=��V����j(��u^_pn9�R�x�E�,q�K�����7t���q�k�T��]�!Ɂ=Y_�0Ls�uI�D}p��\J��������9Q�ke�!f�M�����7*������^So��S���R`[nC��D[��>ӳi��DV셖��5��OQ�թc"#�,^R#UvGI���ɗ�l��b�B��%��EԿd��~)k7����[)�Wy�����0^?�e�nQ�`��VtQ���=@t� zk9�i�%&t�#$6���y��j�W-
�qb����'�^y?�����t�̙5I����Φ-�._�zT:;�
��Z�:d�p��I-�����$�&������P�dlR����4�J/����F(�zc$��2,���,bŏ�\}� Z�L������gf�!a���v��yз��ܙE��;Jҋ����$�C^�&���kEy��ʤ |��tG��	9ˁ�i����If�Kx|�Y̛�3^�@�Ia\��d�K����9#�g�V�g7���`�j���Wٯ�W�5p�����}�?���k3y}�~ũ�ZA�֙���}�^ʬ�6��]��Vē����h0y��e�%{��6}%�P�c�vI=f$ԓ#N���\Н�߃H�����$g %�Cb�5���
�;L�8���|iE�)1p�d���g���P�8�g���y���ll���!v�`F��u���}��bu����O,H	0(E�� ���(V��q܈ևi�s-H#�8�����7t�VR���_�/��=F*��N!��AjMe�>�  ,M>GR��]Bm��B��&_/�2�>  �%�sI������5�`����lxA9;��o���"<�@��[�i3�U0��nũ�Iھ��=�n�!�\e��c��"cz�Z��/hf��-vG��j��=�Z�� �����j�K�U��e����Z9�ֽ����ʂO��<��!Y��,&j���:uD��\}�ͷM�Ihes�Y�R'�7�t�tJ�f4�o6�!t�ۀ��m �l��xB?�[\GZlF/	�ʀ�|�a���2��+7��?�,�Z��~u�X,�=����e��	�Ԭm�-��g� �"��[&_��#)��������v��?�M�E8i(b��Z˭pv֕��l5����f\��1�T�tc���VBnd���~��uF���?)Z�5��[4ߌW���wX�BD2���ܟ�d]�0'4�w+?�}F%~H�j��P�ǽ�xƭ�r�+�/F4��}5�g"�'�飙NP'���a)d2�@	��b~�
��0��#�VX-d��D ��#hJ]�)s 
�����Mu{��[$�+���ĄSc7�1tcb�XSf%�,�,��=�����\H��V��|�wyz�xH.a��~���8PB���s�&b�G厖�̯�/���#�F"df��q:ւ7A�L���6&iT�<J4ƍ�Ygri��x[��܌�I6���m^��~j��tl��{�$��+��g��ᙽ�5�٨�'KP5�6k����8괣@*)�	���e[n���Hab��ܷ�����6�B��)�Heʉ.��RF��	am���#mCwOec9��I�{BZ6��p��)�9�$������X-��i�3Z{Sc�[aI�RSl���\$lF�W�]G�2�E0��r�z��[��Hj/� GJP�jT'��.��6�F�৹
�D/f'V ��?P��Jk,to��<���y۽RK��R�-��?k�JK���P��߮E`�T�� �Ĉ�-���������� ��O����e�R�Ѳ��?kb�@�lB&�;,_o��.��L�-
Q·¯����o��k(Z)x1[�|N6�	������b؁�_YJ��:ɟ&'�叿��f#{������P�Ĕ��I�	�
�i��򿀻j��<#����[gM�v��{�K7���f���$�ҧޡ	��H��%�k���,����|���Q_O@?�EE?�Ӥ}'�O~���H����i�ph�k���'��Dv!�������!a�OQR��4��T���A�1<ja>�Ffg�*��pj3�s_��h� ���z��h�'� ��b�92#��gc� 2Uuy+yUV�3x�����֔����4�G=���c&�~�_6�FǕ�[lNs �+n���#U�Oh�� 5v_,�8� 7`=\Gh $�N,��Z+Pa���t���r;A;x)Wr�*G,A=��[pG�Ֆ=R��jQ�h8�����;�Y��XW�37���Ӕ�n:�<����1��!�5�9b`�B���ޜt�s��<�h锤>�\̬��!�^T0��è��`�O��?��V.�ēD��xc�߆��7j|�����}�0��NZ&<�Y��������(K�9L���ܟW ��o<ܸH^�̩��عͮ1��}!2�F�&\��5��G�y���c7Ӏ��t
��D%��=ۤK�:ofQ�/�7f���v���
]g��J�0<Fn�1m���ӵ!��0^�����k�(����I7��a�RѦn� n��i"�"��!���Y��Ď��5�S��6A�[��7U�,��z�f�,��'�A)K�v�Xpe���t6�r��xO���`���>�s�u���y+(C�F�:��ňn,!=W�窶��%&z`(G�0._���#37���u}S�Z���]�!����σ�'")�"r/{�C ���H�c~6�ݬ`��Ѓ�D��Pokx*['��;e��c�.Ņu$d\�h� o$7�F�u�$,�f��LM۱q�=�J��۴g���M	�mE��Ā�F�}��u�Y�<)0���}Ӎ��;��~����˕o#���*�j8�(�ጪ1�g;��S?#B��o�0m�Q��J,���5����4��9)��o��oU��'	��+���@;_�P�w�67�P�s9�iJ�[v ngb ��h�J��&3	�㨁?jS٧�&�T:�rEmy���a���Y�^(������Oa@@V.h�Bvz�p������~�Y�<��ဳo�C��96���ƛ��=1[�xi`����P�������C�(��3r��u����T�����8�?�+%ޗ����h�Ez0��M+?����-���z�r�B!n�/w�%K�{�����D�N�@�ԩ=&�"鄊C����Q���]�-���8Dc��LrQ�;?,���S��ǂ[�V&�5am���L�.�!�<?�Q>դ���n[�� ��G���!��ԋ��Ofx\���č�7H��W�H��YB�x��$1X�ӡ�U��W�3f��P%��gВr=�u_a�ԣ����~Đ-Sd�#��kD�+<��b���9N��wV nh��Ɍ���K���io��Z�7^H��ם���R��'8�(]n�C��������p���o���3đ+��&��++)`4e�z��6�lֈ�u�� ۠���#��y���̰�����fP6���߆V*�O�c�w���р�" ����~�aZ�Q{��汱J����CZ�K\e\L�𭹮^Vݕ�2�����y��({چ(�-�͜E�]"k��E�3�w�ʈ�3�f��G�,��w����	<ø�<��#��]9�6t�4'�1��� ;��	-xسL䴨p+9V���x,w��$��
EK�2�Xž���d�*��SuK * 
kѠ�.;q�b�p�iéw�!��Kd��&]w��鰶'&4�]X�����\���o�E|j�&��*���p0J�%���E	v2�mA�s^������_q���4���6=��uNӬ�5�����"*LyO�L/�[��g���+ɔ$t�y���f�m�x^2R�㬅�}�k�������b	������qi�y��gt�Ȭ�k��8�Q�!� �qJyޑghR���>R)O�5�j���2rJQ��c׫���F"��\� �y�[Qi-_�so�*f\݃3.���Ho�X|e�C��1��jE`�.��C�k\��s���3E˰��X�me�=,��<͑y��^%JL���Ǣ�t����;	������r�q��zR$܇�Z�!E'���_�Uu4�hپ��O'-S��0�4l_Egw��8��[�`�dﾮ�LZ� ���7�����,=T;�ZI���>�9{��F���q��40�'ǭX��r}q�"�l"K�ggk�H�Id��z��:S��C��r�Vz��D�0$�U$:b���*���#��D�b�A��z	������!��h��'m�c���9띤�o���
#�1��řsJ��t0`�Y<�!מ#QUi蘓�����cZ�>e�����9'5��Z�:��F2�7����(:]���]s��6����$'�18��]�?u��NXwF���k�D9��M��NgI����$BE�B�͟y]�&�0��΍s.�o��s���K������pk�gk�� R�S�jԅX�fTL�@�i�
 �����{:�t&�L��ܷ������ژͭ�6q��r�d�X|~-���4&j�ZA�+�&�L?ӊi��?!�B}� ��`	O��Մ�����"�a������6�aR�����v����8os�wc�����ת̤����������9i2c�S��Ui{	ޢن̏��4W��"�"�@fe��6O��c�ǡ �^�+ޤ@����j��4���i�e<�_�b�jY�|:�U]z�qhN�P��fo���OI*6ۮ,��KPȱy�/���ǘƌjLYdX�#�zx��]}/�Y*z�� �HQ���הd������w�Y��k��ߣ�W!�Ѧ�s��V��0�l�����q���3��EW��$�z�>FC�;�1n6����ټ:���O%��i�1b�q�lPG�]*����֯�5u��"?��NŏB�����Vdo�r���S?yz�t�PZ��yU_��2�:��N�^��R�¤6����Ɓ�� ���j/US�:�Up��@!$��/�n�uBL�)��g>��J���m��w �|n(P�2�N7��"�J��S���ߨ+2�)��Sԡ'W�c���ma�H �C)�4v�1W���mҟ� ��y��[l��p�i�L�,ZМ�W����d�4������yiF�+��A�*����n�NsI�,`�.y��״���I(��Hh�(s�&�*���Q�V�+獺,�`p3�
���v1�y�ޗ���0'�T�D�-#w3���ZGܳ58{b[.v���Ft�� n�!����V8H�5�Ln�|G �V%�DX	�b�~�o�����o�@�o���=�lF^4>��Hֶ���"�x�(��&��o��,��1GL��6�`�l�w���Eg��מߚ�"y�*�p?�zB��d�cb�u�YfL}��3�X�"�� Uꔁ�A�0]�<���N��}kB�qx`���3�I2BތH�ry����F��h$��h����	ؓ�7���.F�����O�KRӖ��I�#�����H��:����?�T>�ɠ��uï�Y'q��=�`.ge���ݙx~"�ҡӲqky�F�ĠN2�AN��NK��Ъf��tf�!�����\C���⯘�".|� G�#r"��D(��у��2�y#@��5�z� �� ���W�,��T��߿���fV��<���o�0�(D-G�0�\�d��<������s��O֭����K�̙���ͽo-�	���}���mӚ�y�{����w�O�Jt�<>V~��n�qϧ�u�pbj��'?g |A\|�:��i� `���r>��'i�sF�>WL��'V6Z��@�6�c�<�_ϟ��Lc�!PX���>L��9w������ U�wCx�09���׋�ע�LfRpɤ]2�x|SBx�‿FJ?�)��\����}8[A��­X�z=�� ��S�b�1j^�s�
���(Q�
�3�����#�k���g�3m�HE2G��l��uYXH�Z�u�2�o�p$ 5�� �w�^j~͈A+T�l�p*���1z��Q��I�&�JB�����i��U��j��ν�:�7��D��B�!����I+��3�t[��1T�ͳމ"����p���r~�&(`�:�)���G�e����v~D8
�?nZ�G�fSBp ��do`Lq��]qQPq��@YP*���Q�R�z�L(�f�*�Ro���tsMK�I��$���g��crn!�����=wd��c�|�h�Z(�O�"��o���ygtb��(�����^��;�+�;r��[�W��M���pl,�-���/���*G�#�����C��-Mhq��Ê��X%.?w�%�Y$��v�sd��n�ȭ�\�����Q�H�w_����Ҋ!X�HVB\�D}�GK`�䋭r��a:��\ZRSÑp{#���@��z���}�}qV.��	%�!��Qmjvc��~ ��� ��faR���c���}����^�^ݜ`*��e�5���GIS�~f;��4�K������I��T�&�Q�ږ�3Ӹ�)tx���^���t�Ee�.��3 ���Z\E����,�����z������nHlf�	gpZ��4!�9���>���?{c`y"-����kh���l�d^�3@����I��~��������1�2꫺������|�9��$�uS�"��Sܟ�\rL�����}���,�)n���
�<�A�&�%��u&z./�N2�k�?{>�}���5�1�Jb��