��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ���������J�r�d���¦[�!�)h`Aw�JC���.<�œ8���:k�zYD	z��OԅT/ur3e�,p��֐,�=l�G��ź>�yZw�TF�<N
�{��\;�uPS�}4�"�mz=�/{:��X��F��V�z���|�P���>LF��#�Z�P�
��˒Ut�R����k�C{[�~HDDc��?���+�Nz��W'����۔�`��d���r�C組kj��]��X>��Pپ!��ѥ�R�G��@�UȄ����K�c���e�9[��:d2���dE�Hd��r���yͿ�I���^������X��G��]�yo}r
��@rUgyW���4��������zx񕬛�C�blP�����nt�Y�6���v<Jq~W����I,��?���_�Ŏ��W7M[*�X��^�z��k��©7�u�z~��u��6��u���q�>O�f ?��-դ+����z��W%Jɨ��ДlRzh�7�=��N��Be� �%��=��,�'��
�f��,ՠ3�����r"��c4uхC��Tu:*�'q���ۀǓj_*~Cb�r�u�EI�p�G#K���]�p>3}]:v�L��#/���{��N��'ɞW��t�����Q�e��kX�X���,��m}(Q�Y��:ҧe���_1�Hn���|e�_Y��L����+0��U�mp84�y��C���M��=�6��]�RP�8��$["sq� ��x��w����r�փJ�8�.�ˁq�(�L�Hd|��ꪃ,���8N�o��᛼���j�Fg�5*�. Z���V��J��Q����}�1�p�^s�j�G� 	pLwp��7�����#A��K~x�I�C�I��䙕�	���U�U�\��<�i$W�ɽ8X�+o'NÆؗ���x� ZC3��c�NRp~�3t4�1��T�Ц���_�����cL^�;��]�?���o�e�]��2���7h�O�\ Q.��n����ȬT<d��4֟��+(�k�`�Z��h��P0�1-h�!�}�Ͳ�d�5lZՎ������b5g7:F|j�__�p21\�pC!+��tF���B�;��=��w���O� ��/��g�ʃM"�qjN���~Q;y/�#⡂V���Z��J���ݦN�CBѷ,��t�\v��aB(f���)&89 �1#�2U��A-B� ��'*}Y<����W�����'��$��~���*�Ps��Z�_�P�3w(]��z;P��A ��}f-)9۾��e��*!�9xqq�(�3ƣ聫��~x̃����O-��� ��h�h�0z(P���g���N=���Ӥ	������.Q�_urHk��?x��1����+��ӗ�b���_��)�F�qH �`�y����}:��t���ͱ�}�N]R�)�m7�����/���z`��o�Z��i /L����ߍ��H��X�/\��� k����'%'f	�ǜ��,��F�K�ߛ-�����=�M>�4M-4v�)�����K��T����ٖ�pGQa�p��
���D J�NXM4���s�uI��bP/�	���H�@�5�qG��P�̵t�Y��_��sWN�U�A�N&��ݕ��e+/���s �o4֧�-�x���E��-ٱ7�K�J9��*��b�m�`0��#�3��7�mB�J�rf��H]����q0K{����>�?#��%+ipL��%<�M�qY���;�'�Q4j�_����x��|5�Ɯgl9�x��Q�U�	��ֽ�~!�Pv$�X_�|��A�BG�����#� �?fWC�;cں�f��4��`E���85��+�v�����<�bZ:r:��V��$mAF{p"��r�"{��S���V!�a4��J�H[���I�za>���|�@}���(Y����Sm�+�3d��~� hZ�H���]��A3�L�>�� �2�����$����JG�تs��S�58gʿ)㫐�R��J�S�\8X�2��;�����-�����r�hI�o�]�>Q� ,�5x3d����`�!8ae�Kqۢ�n�{�Et�Cν�'� ��Gce��>[��D�D�!D����S�m����W�K�ɜ������]����ӛ�{~�.��upD&�
�^m+�BI����N@����@G?��z����q��2\�C�m���?t!���e$��*��Gpʍ�'#b�U�&�8��㊟�g��	�[$|O.yW)�N���_{8QEPo�P^9������so ��*8�����d���7+.T0 wc��8JP 9z�TY5��$�=Բ�C�¶��j!NCb�$H?�6EZ��8��07���Py��l2�+���?j	��2��ʹo�N���;u��n��.N�h�8K��Rq�fw۸��M��s��X)qdݏ7�C��s�8h��L�JR�>����r y,��Ȇ�D�!(���a�L��ݙ��^�=fV�8"��L�1f]I� ���,@�A�� �B���t��6V,�P��%�����:��QB�0Y/�Ժ���~�e^w��	E��Y�7�3?�@�g	�?�q��U,�ǖ����C�{��Һb"yH�9�Ʒ�L���nw�ߖ�h�f����e�ʺ��4Jv4�:^g-�4�e-L{gݍ�3���:�g�m�ڢ��$������[\x����
�@i��*�u���&մ�s�G�ߘ��Ea�N�ѕ��z2O������ʇC9�û�xz\GF��lo�q�c/.u�C3��.��p͆��\�av��]ȕ�O80��b*�gZ�spdK}}��[�ri�t����,c2֗|�X;d�d�,�CM��Y쁡�55e� S9V�?�O5�?}k���O�V���DX"��m�K*�ށ�=�V}�%k��t�����Qnʘ����_�����^뽛ŜV+�ct
�X�����r&�ƤFj��*�.4�g��G���:�U,GR�0�,?������T�U�������yY#\;��f�l��4�z�c�Y����?��>,���ԎQƈ�}�z��|�l��L�o$�؛ E�$�j}nu����Ce��P-�-4�/�p+< 8�y�+Z��^�+���d�-^�sJAr��d)�R������ҙ���S��v�F���1�{�l�����Nr\��S���o*U�X�9뜥�x,�R�ފ�}�_ǐ<ګ
[�W��q�p���=Yg��� ���h����߷����Ke�ߚe�N����$P�:]�W<!�!kI#�EY>����WA�7v)��a�/����Ϛ* F g+q��'�e<�����e��\w"��@�
P��p�����L��V@��+�ւ�n��ulN�3�Jw(M��O����o�1�Jǋ����TU�'= ܊y4�^E��	�io��aZG�uB�(�a��S�/�5����N"(M���q��J{��p3,�id`�������9�~�0}V��:�T��/��j	�@�D�s�7GUpOƱ����C�E5oږJ�D����}���K�CJ��u��y��P��>ܵR!^V�'�"�&�Xc�Arz�hf�!}{��UG���0�z��KN :�d�9 ��ɞ����l��^NH���̶ƞY�/���m��������%��9�P˶=��QҐ��8���zq<�����Z��?|�Dh�w@���.��1,�(豋��mu��Ժ���#)>5����Ji�&�[����zG",/v���:3�Ro<[��!A]�ʦ�}��U�Ĥ7zA<ٕ���A�`�֦4+�7�+�gN��'
�"��(��G�X��9��W6��,u��H?�������p�w=c�����T-��o�3������E���ʚ����c�L�ǩ��G��Yu},?��AK�E3t�m\MU�]q�GL6,D����
g�>��ᦏ㷅8T���Z�����G�6��� G�lsS�:��=u�T�
�����?��qp�,Ӆ���~{�l=�����`*u�o*��C������1�ҟ���w-6��,8^�H�Vi�y���ͤ���	���ڮ�����v*��yC �gD�x���Hǹ{h�Q+����ۚ�ʶE��Q,��'���D�\/K
�dB$cI0G;TGY: ��WEWx�>�{7�0������\ŖV��\=i�����<�ڝ6Fq?�rv'��ȇ�e^k� �2�a�|����_��g�|���tA�A��6�*��L�Ꟁ��o���X:@TV�N�ֵ�L����-�BWw.�.��S�Q<�!�d}P�H�(��/�y=�]TE��՟ˑ���B���+�][��L��n� g�V�T��n��.&ճ���^7�P��dVh1uUHj�U=��b�5���f��0�����ei��KÏ-*Z�
�<�*�~���"���@�K_�s�E�kp�vȱ�+�3����v��*�ÃO��.�r`�D
ٓ �� ���Z_m�^+������t[���*&S��Η�*Yr�d�z��l�{w$`�z4[����	)l�����+x��c�q�F��S*�{�����x全�:�	�G}ڃFM�?!wii�dB_��Z�k�����=�OB�0 e|�V�$ҏ�y�U�=�
�Ufkچ�.L3c|���К�cp|I���,��h��ȧ�_':0�ȧ��d���@	'H��)��[�Uc=��� i��ؔ���]���������`��JK�K���i��*��#�w ���o�� #�3n�р�Mך!�2T����zfw�3\��f1̇�� 	�|M�;p�;�j�k&�z��*�>��:�_��P���㮵�R>�(Q����Byi;2	��,�!�}��ON��R*���{�y��E��*�����F��}�{	0v��;i�t���ɜ��8II����VJ9ϠV��2����f��b��C�ǛL
�տ��=�.��&f.٘,w��;bn�X��'+�J㺻�N�| YT-J~7ա/N4}tSH^��vI��5n����r�Y �hd�N�CR�S�J�{�����V��ҏ�f�d�)��u�������i�X*�7�7�A�('ψ�a�F_a���
>MG�JZҷv���z�q��f1A���:��p�
����f���^{ͷ��t�u��SV��#_O�����G۠bxX���eܾ.0���!5U'��RP�F�`�5���$��5E��މ9��OU��K�)V:�ߕvi�QT�<]�Z����e�$;�a���i�V˵)�������}�Ԟ�ᘤ��5@�A���S9>T��߻�@�BR��
<dRZ]���¿9���+BoV�?�C�>�v�AW^����<�y�lǜX9�GS =�&*�(ky�S�fQ9�1l��.VT�Y��	u$�� �!��^&4��?���sC����#�C��X�!�L�_J�±рc�LFPB�����)�&�e�`� }��(��͓͞���*�l���6�8]V���L��"���$�~V#��
���hdV�Tܢw�3�F��(�3jH9�k��ASP�,y���J�j�I:f��#�����}	N���G~�Âi,���s��K�l�����xL�w��}��I�U>��m�V�x���Ԛ}]y���:_�wϙ��i���;U+d���/��(x1�m#m�7��Ti�/M:x�>!ѴO�c�a���@���lcT���0���jȔ^�A�5����X�5�0YT0SO4��Ǝ`�1����d��ȓr��M�&G(�'i��4eq�"�{C�ᘁ	�[��@]��%T��-�F��?����1/MՔ8�2r9d��~�]��7�N0j�A�"EUqرڳsc	�ybqxJ��J��=RgO��~�ߎ�@7��{���2sd��97�ux�+$Υ���T�7�{q ��}��L�����ӯ��x(Օa3�e���)��8�"����=Wɮ;xI�kg��`m�}|S���������kr�,�d�j�Q�9��F�h	w\�1�锪�Z��O>�|+2Z8��g���P��3[(G��j�w�	�r�|O�^i�:�3�NZ�i%�	��?Lo�w��{u��������1:�|��lC6{��&�ZT�Ar�{����^C9�����ES5�o�Waϣ�U��'aS[T����\J���@�S\f��n����Y۷vz엨�}����\KU�f�wFw)ʗ��F� e���T��.�����#F(C���[!�!�F�@���yʛ�:�zf:ʸ���j%q�����\?`�o�!��)�o�
J�\i��ʴT�Ωk]"���AW^L�^�������h����3�:]ю]p{��Q�5�ۡN�_�b��?�3b�?���4�=��Q���މ�'� Ǹ�E���07bL=���I�i�v��A��N*�G$DmSB��~���
7Fؕ��׎��&u`[�h�T�?=��8����Th���h?%?Q�+��bGW���l���Ӿ�U����Ŏ�eg�����A�>L�oV��g�� v��?}}�����}S��\����2�0Y	:��y#�]K`��Y(<^��͇ls?~p;1�2RڤK{NǨ7�ݗξV�DT�"�f\ bp���C(A�����B�
P�,����E]Z
���iIokowg�� �Z"�̩�pF�����K�F��A\�k�lU��
BS۰|��֗�� �W���C%�|�H_�RƵ���7�n������&� �Qr��}��S���{x���"�\�l�B�v^���V-"�	��o$ќ�<�Ec�n ����B��f�M�����Pۊ�C:�/c���0��x�FefS�~n�矎��e(#07|h�+�;�Ј�Y��G{����TJq:�w�Q��[��J�A9���	R��s�c�F�~^�{H޾��8�o�xTC�������r�T ])Ϛ!����2PiHa��h�1�4��zrK����{�pfc�#���;��0	(+���z��pfS(1"C�����KG?��X��):��FM�w?#�mf�ۡ8�����˜�z���n+n`�� 1�?�Wg��p��#r�:"�Ӵ8�J�3œy}���o��F��Y�������)T^�� .ݏ06����I�k >�B���dp�~��̀,��81e"E�����}�9q܇R���Ӹ��"��ȗ�yф^j���E90?&���K�M�xMN�Z/͚�
���&G⹨�k͌��~��~,�8�����?���>�,v���$D�m��	��k�	���ukl`��M��T*� Y���o.כ;��D�Y'��ǃ:��Fe��2��hz�z�/�y�vL﵅Sk��t�.BC��x�����y{���c9�ˀ~E�))r��#��3w7�}��H�ץ@�'�k��V���$�'�6��#�b�٨�����ɠ^�|(#�&���A{��K��Qr#�j�d�ioȻ�1(Av;x-4��L:��YΖ()��Ε� s�=]�֢>ق�xVX|��^)�%kt;j3��b�'�j� ����x�5������Pm)�Ȗ���󆜽	�4V]���/�L	m�~�u@@B�S�j�)+�O���M鎍��B�{\&��PKW��4���F�IAь;O�6Y��bf�k�}9�=;ѧ�0t��Wu���"@.��r�bx��\����O�'