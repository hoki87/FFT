// altera_fft_tb.v

// Generated using ACDS version 15.1 185

`timescale 1 ps / 1 ps

module fft_tb (
	);

	wire           fft_clk;   // fft_inst_clk_bfm:clk -> [fft_inst:clk, fft_inst_rst_bfm:clk]
	wire           fft_reset; // fft_inst_rst_bfm:reset -> fft_inst:reset_n
                  
   wire  [1:0]    FFT_num; 
   wire           CP_type; 
   wire           FFT_type;
   wire  [15:0]   Din_i;
   wire  [15:0]   Din_q;
   wire           Din_h;   
   wire           Din_s;   
   wire           Din_v;   
   wire  [15:0]   Dout_i;
   wire  [15:0]   Dout_q;
   wire           Dout_h; 
   wire           Dout_s; 
   wire           Dout_v;  
   
   
	
   LTE_FFT #(.BIT_WIDTH   (16),
             .CLK_FS_RATIO(5 ))
   IFFT(
      .Reset   (fft_reset),
      .Clk     (fft_clk  ),
      .FFT_num (FFT_num  ),
      .CP_type (CP_type  ),
      .FFT_type(1'b1     ),
      .Din_i   (Din_i    ),
      .Din_q   (Din_q    ),
      .Din_h   (Din_h    ),
      .Din_s   (Din_s    ),
      .Din_v   (Din_v    ),
      .Dout_i  (Dout_i   ),
      .Dout_q  (Dout_q   ),
      .Dout_h  (Dout_h   ),
      .Dout_s  (Dout_s   ),
      .Dout_v  (Dout_v   ) 
   );	

   LTE_FFT #(.BIT_WIDTH   (16),
             .CLK_FS_RATIO(5 ))
   FFT(
      .Reset   (fft_reset),
      .Clk     (fft_clk  ),
      .FFT_num (FFT_num  ),
      .CP_type (CP_type  ),
      .FFT_type(1'b0     ),
      .Din_i   (Dout_i   ),
      .Din_q   (Dout_q   ),
      .Din_h   (Dout_h   ),
      .Din_s   (Dout_s   ),
      .Din_v   (Dout_v   ),
      .Dout_i  (),
      .Dout_q  (),
      .Dout_h  (),
      .Dout_s  (),
      .Dout_v  () 
   );	
      
   ////////////////// CLOCK & RESET Source
	clock_source #(
		.CLOCK_RATE (100000000), // 100MHz
		.CLOCK_UNIT (1)
	) fft_inst_clk_bfm (
		.clk (fft_clk)
	);

	reset_source #(
		.ASSERT_HIGH_RESET    (1),
		.INITIAL_RESET_CYCLES (50)
	) fft_inst_rst_bfm (
		.reset (fft_reset),
		.clk   (fft_clk)   
	);

   fft_source_bfm #(.DATA_NBIT   (16),
                    .CLK_FS_RATIO(5 ))
   ifft_source(
      .clk     (fft_clk  ),
      .reset   (fft_reset),
      .fft_num (FFT_num  ),
      .cp_type (CP_type  ), 
      .fft_type(FFT_type ),
      .source_i(Din_i    ),   
      .source_q(Din_q    ),   
      .source_h(Din_h    ),   
      .source_s(Din_s    ),   
      .source_v(Din_v    )
   );

endmodule
