��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ���������tܹ�< �E	���Bh񞲠Q/�T9ÍJ�]͛0�S硢��m}�[6� �w��E�w�ӆJ|o��>��	Џ#D$Ħ&z�C0z�����ͦ������K�=��?��Z��_,��@�ZR�ͼ��ɛmF���� �H*���j�P�KH�u�����33����K)>��	�+=0�������w��J0���N�2��G����$ߨ��K5�J���u�L~�;�ʢM�����a�T�GJD�6!�A�E�t4!��3�a�>X��/����`@�ᴹSP�gR�)���PV2�x$n7y�qSԁ�De�l��}�,X#���9W����n��p��;���q�Ӻ����xQS�'��K�a#] 3�a%("�C^?cS4�{!������d{E�W�T���x	Oe�����/�odS���4x���vp�����u�PW�p5f�U[k��$���UCM̪%�֑��>Į�%߸�<�3B��)?��}8T~'�"�c����3��v�����D�V� ~�.���G(ޏ+�A�?��#��ݳ����Ji�^ԗ���W�����6k��q@�nP-{pD�M�TL�#p�;3ǁ1�bD0ǃ�IÂ8���AWэ�
��j�y��P��.P��_nv>��*и�,���s�����{����@I�3�;��L%)������8&����Qu���G�=��Mg@Ì2�[�L�(��`b\x�Ë	�T�ː�7�Mc��|�P/�*�J��I
��2��[&�=Nߗ7�k=�#��=�����օ��Ҋ�q�~)6����������D:�+y�����|��;]�N�-�t�X��؀�	l=��(�}Ux�WOG�/���A�[�2�+jr�]5��y����|��=��;�܌n'�q0��v&���@e������kz��x�l�ԑx;�YjQD�#P9����b��w��ö������F�	���������VN�sgp��Ki���~*��z��l���w��t�Rb/d��5�Հ�r'R2���O,�Wlxl7�ܯt�o�#��v�?|��q5����hڟ����|t�Q�A\�f�PNH��N��x M�����O���$�9浘��#���Q<�,v����Gb(�	V$�f7�2<��:�E����T���Ï�b����EZ꓁���*G#�D��{$������Ǯ�4�ɻ,�ѡ�u:����c.b�c:�&w�����_nq�s����$��)�����~no�X-��,�B�Q����
6Rʾ�>��	�:����w�j?'����X6�ĳw�����{7+�w�_i�?�Z[۱����2J��)G������0�T�$Uُ���N���|�MF:�#�;�Km��Y�=��oͻ�	+J�r����l{��|� �f�k��*VP2��%��c����ᴼ�!D����E��k9i��Z0��	�b�T�se)����1OKϲ�5i"�ef�������I��kJI9��D��}�?Vy;.��È�O�	�&�Ó�a8eҦr�Լ��T�BXR�c1۳a�ם�M�I������_5mPd�`��a�T���"@�tl���5c�e���Ѿ�n�"��^U���O�:p��"Uϭ�Qn��}�ѯX�}=בf��܍�`w`M'��a�	ne���V�HT��W6s6�E�D�{6��>ᤉ���-+�n�Z��÷n�$nFX���ZläK�	�Oz�y�p�pGzKq>������f��[X�шgO����B���,�1�TzF��c.��[7���}O�c�aȢ�6�j�%�T��1�o���w�_R�)�9w"f�lH�ep������-!j%��1Z��C$�r�2�K�W�˹��skY����b%uΚ�xv��s�t/v]�7��J=i���-�-L?�ZF�hm�<��~�;@c�v8�hfWw,%B֒3U�3~�20�<�OL����p��~א�l�Ev�B���'���ܽ=B� Ekʡ�m�**VN*e|"p|>|�,Q��3+�7�-PrY� w�QǦ}v�Lf³Q�b��ǰ�A�$\�s[��RS�1��T����Ѿ]��e�٘pa�^k̧���!�JC��%�ú*��>q	�����w\}�K
z&�W������
�tE�m�b�OZ+ܔ�s� ��ٶ��9��ՄF�[v#t��W�ln��p�G�Wj��0Ʒ�vl �g���[�ѽ�֜ /�Vݖݔzx���B�L�z�����V�ի ����l�/���P��זD=:��,�� +����u��:�C��;UZ����FJ�E�
I��E��i��t.���j�o&s<���,�W�"��]���:�!��:���a��z�썩	.ͮQ��"��ٸ<׬/t��UeR�!/_�/�є� ��i-�Z�Y׾�2�`, )9���� /��:��S(�E�/wܤ���H7��F�w>h�e+s#��	�o�G�4���;d����=VJ�\�N*�R��>�ٜ�r�4l��}M?��%�O����:4DgE�ͩc�<?K�s_��sI�ܟ��I���%��xx�פ~�\�8�_��J�t8��u���,�)a�#��7M�
u��Pj�fb��B��9�D���K�4~UȾ,�oK�R!"�r�i�����P�`N|M��j�K���jI`��g�'F�:6��%����3�9��T��]���cV�5 յ��_�6F\q��-�O�5Ne�p {�g��'[$Ix������ߤd)��q^��w���-��#���Aa+EKl��}��ft���3+b��U2!������+�2bC�oWCHJ�掍cjU�7�3�I�N_fW"�0�o��h<ǌ���/��8��U/*��Ȉ� �jK_��_�j<�ó�h�@��I<x��n~G4П>a/Md)��I�m���Dȸ/�%�}��\�h���S�N�p���>i~���k&�3�cØ���ӡ���ۓ�Q�\[Z���:�rƷYX���qO��K9�����(-�v\�}E_�܁j�+���/܁F�Kg,�ɽ�C�h�>�	}�-�)d�9�긅 �(�ߠ�2�8���LyIOG�#{i�����D=�^�sm&���=dn��ܖ��פ�{�J�S��v�.	��2PU�e��2�c�	�&�|��Ne1����1�Ԗ�D�1O֜L�wt�ws<�r3�3�� ��N�8��S�읨�6���.�p��#�͘ī��=F���-�J�ibH�B1=�*�����X��T��4A��"��,����~������9Zb��@[��̔Zm��p�5�#a�� !7x��P]*���N��f�И�T�N�b�`!"Q�3���f=FEB�۟řWK��Y:�p�~w����;t��j-��(S������s�>��+���B�9?b��090㔫=H7	��,��8�ڲ;�y��-6����DT���V�����y�I��`�5$�������E���G8qnݪ�BH�����$]c<��g��0���C~����c��ԇ�:42ǩ�'�wQ��D��&���9/t���� U�8 �2�1�x\�2��aF4+�0a�h�n��)�T\�u��.�6�@��Ѭ��As�t�94b�i}�oĂ�	�	F�'���O�D�/.�Q���H�^���%x�{;5k�ngFZ�Ɨ�dPQ��qe�aL��ܟ+�)���������U�C9��$%!gB4;�%yJ-��	!C�a��ɚ��gڒ��u���e�2e�&�{>1;f�a�ˡ)=�
LV�p���Ww�ꓲ��G��0�iE#n_BJ�k���nO�e2�)9��j�e�C�D��8K�\�`:{l�e�*�_��Ȓa�C������>��;'���<U�/�[�� H�a$﨡�ۡ�&�Q�*�]�ѹ}@�2o��
W	~��T�5��iOd�U\�ho/��B·��R� �b,�wB�f Qn;��S``6؊�3�j����fcJ���{-Z0��TU�â��%W�w;5 2��-���R�gv�����Z�=���u��-��l3�싋,������X(f�V�%�l�h��4w�ZӲ��_d��0m�e$�܆>K9�[�j&J �T�끢���,(x��K*%9� VU��
��D����E/�$�+h��B������i|�U�A^�?�*�#�A�2:t�LX�K� k�V�
��g�.}�Y���]y� �?U�C+��0�f'�,ᰣ٭i��>#|�3��xi�+�� ��Kއ�ﯼ��\�|g�V��s��kυ�k@F��V�����r��h���r��D4��w�e������cϻ���jSΩ�s%a��F@KN7a�Zr<�kD�������e�$���DU�K���'�N����HܟB���/Hʒ]V,Sy[8���^< h��]�&��g����E9�&6��Wz=Z��M���MǯP����3>��K�vˈ7�IMBd�FU�$�$ cF+��i͸��@7!|�a��<�Y���H�+I��y�kG$'��8_������"����V�bڮZ���BP�re��x� �����`m�58"m)���<�iJ��t��Kf%��.��;�f��;J��Y������'W偺ؙ�(x�O���,���֑�&�NH�*r���]�cq����Ҙ�����~@�t��� ��Z����-v^G�������P厞���M���X������!����-�Qx`W�d�9zf���o_�LN��7B2��H?�h�0<ȡ�g6)W�	�_�4�F'��|"A�ykD��ﺗ"��Q,���'k*w�0�C$���S�)�E6��W��' ��F�1$����6�L�ILT�R{�����O%�%"j�k��'w'�<a���3PM����,ڟ���A9�џ�۰͈qyӇ���,��'n���
�wCx8�OU[���%�qy�ߊ��5�*t�_n��=`z��&�K���Kz\h�}��d�(��ᗄ����D����L�.�x�1'�l):~Y ���"n7��3�̄,��W1{���ss�y&�P�7�gg5ż%3�[��Z�9�O����3��fЩW�!k��ŠIZ�}L�e�a���25�Q����&r�M�z�a�q�#r ����sj�7������>m�{K��P8��Z;�X��v@Xo-$r� a-]豦 �^�{���EjRS�5�iy}�������[�b�m�QQ�ZY�ɳ�1�j��{�Er�!�>���佦ON�UF��Mcf:�l�7\3���=U,Qk�)��X����t���L�t�G]��V���V��fN���g��AF}j���wY�F�Qn���Q���MY�T�圖ZI����6�,��ޙ�˅@��#��|MR�#�
�����[��w����SK��c���.���
6v����9\Z�6H��BRq^ta%� ��������|��V�\������uZ]�f�;O���jD*%\�6�� 5I�g�?4�m�I�t��(��JE�(��IC��)�%H3�{�^h`�2���!�nJ\O�?���ağ#1�M����Ur�E%q#�m�˥�:~p#�0\}[�X�F��W2�II�X��LS	)���k�v3�R���ӻJq���>�y����@�o���Qk������dLalC-�e_K>.O��pz�Q.;�h���N�gh^����J@�t� ��H~ա�5�8$�)x p�t��tpjr9x�)�Ѭ�:��O���X��%1ۉ��[`	(�M":�	�o+�W��:ԁ��7�|�">J� ~������%ڧ,�:�zK���ाA��qAu_�~��G(�����?��%�c�]�!���C�Ek��m�HY� �\�։�5�f[�!u�l���\���ဒ��ek��HFZ��S뢸�8s�3i�ZuS�"9ظ�x1���6V���?B�O�qMCrs!���噏B'��堔ϱ�#� �Sr�T���,��+����,��ڟ<����,��2g�yI��~����n���	9#��4���.ΜZ����M�7��a#��lH%�<�-��#y�P<�Ն��Ή�Vՠ;[�	�	��~����`� �|&�e����քe0L]��rŲ85s\�����qI�t���c�v���/N.XD&y��Q�h�)�v����e�PY]c$�=�?�*!�1͓m[P�v��[R��T��AG'����'孴'��C�o'�"8ğ��yi��.���''X	e۷�:����������9}�D��|+�~l�*����D� q��RJ �k>��_�"ār�'fw9��9�u�/��뺴8T�r�Ĵ'U�2z,!��V�!���}f�)�3P(e@Z��c"��Y��!řp��*�~�+��خ�bu���ÿ�5�ԋ��R{N�4�\��u!4W�5�co�����퇺����+�ȯ�Ļ�/vR.���b[v���*�g��ˎ�0G\��/O�F���I��F3�1���ä^�f*��Q�GO��a+��kAsfˮ᫤��|��,"a�� w�Y����D��%��7�����)k-�ɥ�\��pR�ZSf�^9/�c)t��
z���m&z��L��,-�q��;�P�����N�ҕ����I���d�A|*U ���J$7���v��wè����4Ky�����=Z�.��uC��O����h�7]�M��-��M��}%ɵw�@��p�zk `�2��
�p����|���rTPT0�i���s�q�e��K�������`����ET��V��\F�O�G]��xP������N�A# n��� ���d���S�>��aX�(�J�[3�Eug@��(i�Z�@
��Q���a�"��U��a�e�	%j�\7��#7�kPa}P�Z�I&k���5��̀9�nkR競��R[�;���w�� �mΏQ��)�J��/b�L�R�6���Ѯ��\	(L��k5%�dWS�1_^��j�����?54t���U����X��ScT���3����d́/t�٬���W��vN&��G�x���=�� �fSp�F�M�$�iZ�"����<�	�h�6}ax�匣��w���Ƈ1A��%z��,ƉW�~ȶ�k=UR7#��r�R�]��P�u1ڵgLH����?�ĀJ/���+-Ao�0"xhI��|I".��H��E�z>L��4������acU��k��;�d�-ݧx�7�m�KeyG��X�@�>ɧ��+1ɽ�N����~LNgYH��u/��'W��5�k��ÿ7��nćc���wl*�Q��uW�~�ʕ�U��2���ǚ�^�>�c9i�[ 6�KS�rSۢ���7*Md�\��V3��<��bƇ�"'3��3xt˞W��P���t�q�'N�G=�#�,Am����r�x�ȜRt5�e�v��b�s��A��!�ҁ�-̇��/� nx2܅>%���
*9.a�����p��H�${t�ޠQf��]����ė�2�6�����7�z�F6ԁ%��1�~7fp� �X%�ux,)%ظ[�C�Sd`�n��e�#6���H�CV��x�z������Tͳ?x< �B�8�MDT�����M�2��������*���i7�|q�vG!H�5�8�%Bd�nE�ZG��ZI��Y���ʓΪ\���!z��M)sZ��a��"T�	O��H��e�oı������f!]�I�������y�����l;佮
ɕ�'�����|������]5;�R!V����lA�Җuko4�F�z�
w�Rx@��Xc�ʪ�R(���0*�H�.��pjC���r�"�����5�D���[�Ս�ȗ���`����'�1n���e�Ꝗ��N��y�sz6�Q���r�����s3#�W2���Jry�ᶔ4�U�!�,���~�,-���d]/�d*钬��/*R�5q��_�X*HT�*��'?���|o�zԕ-cQW�𯯌�cXY{T2�w�h�X���`�����^��eVq�[�@)	:r�9�`#�V��">�L�p�/��Ћ� ��c�ݫU�>-b�w�p)8��!��{��C�����jq��'��?K�܈�J�=�XW3O"���D#���P���o~�~uro�;�䵅�ojJ�j������t��_�K
��t�8D�i����"X���|N��ž:�{Zk�Ʒ��g��/��c�6j���z�N*m��2���g��sl����bw*��t 5mΖW(EF\`���IW�z��v�OC�<����c��A�,R����}�� �Q�һ:�y��Q���PЧcu�g(���)ѭ΄��@���	�=�Q&t�[?k�.Lgƽ=��� �c���
	�����Y+6ᕦ�'�ۣٱ�]"з�����i�}���DV�PII��B>ů�6���%>܌��}��C�L���\K�A�o5,*e��y�d�b�AD�C�l٘����"q	�7�YU7;���� zF2s�	�q��7����+�����Eh<[��y���X�3�:F�l�˵�
�g���Mf��f�a��٩��HM>j~����� �R5	7}C�f^�?aj�<������%��>	S$R� ���͖�;Ǒ�����}	!�LS���4�qTi�;�[?{l�nA����j� sѫm
�<���~���W��
�
H�0ݸݑ~�rZ�:�o���>� ��&�r&�O�SaX7N�"���{B���#˜�a�b�����<Ő�_)��`�����0C�{%J���L�w�2A�∭�Uf�� ^?o�'2	$+JsP�8aF�Z�T-.�:K"蛪��d���R;�P~R\���=����'�Zы�nE�>F}���j�۽��w�u��7����`�������%[�'TvE��Z2�Cv�D�.�(��8��^yY.�ߡ]˄��m�����bL0����I�W�/���J�T�u��}�C� �M
'x$�L�v�e�(���@�J�Vc؞��\kYiDw+����s+��<�M��`9���`]W�U�^�]
@SCfd�鷮l��%6�x
���2}\up��#J��X�)��ۃ�=o��M0s6������/2OB(�&,x���5�Q�2ĳ5�"P@�>*��9��V�bS���Oa�Y�<� P���!���
�Nc� "t���RꏛQ!4z���1��^�Q\ZH�{<S+���,�����9�1���S6K����[|ٻ�Mak�N ԣ�Wc�ʹUF��@!��S�W3D��a����h��=��u_�NF�K8ŚG��ky����ɉQh� K�$GJB_�L�fIX>J��:�U�p��dH:��f�6��Ȑ���L�5��8����{N��! ��)��,ݻ� k�C2��:��+3i!.�ˣ�> HpS�C�k�&���2X���~?�I��B&6A �֎�8av�}����x1�~�O�����[ɢ?)��m��7+��I��pW��P�ݬ�l�W�@{�cݟ(�/��70�&$�(����x��G�a�n��M�6W<��r��D�[�����\]EK�RF:#���p���	�ݯH�|Ag2�W�$P�w&�B'J��Ao��D���t�����>.�mN�y5;G/�#@Eؗ$��;�'�DH��4mﶴTh�-���)3U�!q@eB���;7C�SP{l�U{���_&�0=$:�A$!{ď��?��?¯�I1tp����I-�=�y,N�S��: ,���J�o����ql`f��z��#�-Ù�)%L�;�e����ea��KW��)C����O���3�b
'��aw@)AW�Duߋ�ԣ�$��vN��b��loiD�
/4���F��"m�j<ۧ��IZ� H-`&T����/|"�/���|W�0n�e6N�bc�3�7�XmSS�:�Xbn��C�:��M1��^2e����pe��1@0�LY
�y�!�U��@�ʛ"�m���Kll%<��W�y$�J.���=!�^>�iW,�]>�W��n�@����uO��@O͉���r����}^M:cB9V3/���l�=(�R�j��M�d<�-�-Y��"����q&��\0.Г`�)ƥ�ȍ��������OZ�l,�p��ԞC���Z�O����)���I("*��^N�&�(��Qޗz o؄VF�D�|e�p���ѯt�>������g� jG,!n<��u�N�_,��)Q?��DW�5�PlÖ�PS�����$Fq������L�G����b���
�.�Rg�N�f\>�,�Z� U��tP���̾"]�V+�%W/�:�'���ig�Q@c�ⶥV�}�f���[��q���*���l�a;?w��`*���p��: �&�͘ߏ�V�2H�=k^��;�`|"�F{�+�d�[a�U�����4�����a=ߊz!4�6�yZm��j����jh&�H�2���ḇ��I9O�,��ƞ�h|z)���Ԕb��'�%n)̭� ��s�6c"��[g�|pm5�B�r����SUݳ7����&��]x����y8��SXd�v���lX^ґ���#�����(�5t���z��өEE;�n�_����r:�����a��.�QF�z�@�[��Ѱ��]�L��s��r���=U��LO�DH;�%�NX�,:�?�6�5PR�����^_m�2I�X �#���y�Z�5� ���j6��V?��a7�IAN%�R�� ���_�\l
Z��9��-s�Ӹ�^�?�-�2r�I�#�L����^I�6�x�w�t$+����� Ǥ1��╳�Ҽ�:,�W۷���p;%aP�[>��N��0���G'�֬2��S�8�N��{�������1muO�o�\�\���Q�hlv?4�̧ӛ�9�횱U�j.D�����UP��)VZ�j����]�kP�+J�h�ѫ�W^L�l	�Dt���
.�I��})d��}9%�w��qڹu�7��%�hh�<���1C����zG�X�8��%WQ�N���P��=G�g���CEӨ} gE9c��VI��` g{\��N2L�ہC=���9���M�g�݃�>\��z�/���-��\�5��B>^���Պ�G�0�a��� ��U֑s�m�FX�$�B}��<��;�IYF(m ��Ƴ?�P�z���ed�j,������j<G�|#���t��X�;��y<B��|�ʗE���5���8y��,���(�Ȩr�J��:� �Lx#!�N�t��-�dB��O�+D��#_���q�.��#��iJ�?Q��tԕ�0��pw�,�����u뗖2����#�0{TzQ[��n�[D=��� Z9^������2�X��kA[ׄ9��@��������9��v��&+Zy�� �`�n��L�������U�G؊��
e��(6��h�;�%���$i��ey/��@5���<��B�'^�A����f��}]��I������7H�yw�"����N���e�Yw{�Z�:�����\46nb��p�������g��>7�K�:}�E{4Cկ�E��܃ܸ5�@K)��~&Ч�5�\�bC�l�5ţ~�L�����̩�β+�D��.���L���V�U�h�
��(.VE���`9I{��E[��E.����C��ect�{Z5S*��R��]��%N��1�!V'\�Od1J���ʹ�+짌���}�������{GBX�Ŭ��~�:����q ��E(�	.��[�!D:y" q�>����l����os����K�f�����(\~��,�o@��� �\ж����	���߳��%6�o��Wg���(�6$4���W��R�0��%�r��Wh%*.���׌��ɥ 
��aa��R8� ���9S��!<uA���՚���ɳi�+A�U��fE�ʃy��y+����~�=?6���鹍Q6�e.�Mi�i�RR�@�73�qcRዅ����ٺJ*Y0��s�R��du���"��x�J��R{]��F����g��b��6h��IT~��щ4���l>c�&x�a���<�p,�q�߁��|�S�}z��x��B8� ��)�!4v�z�* DY�.`%�.�;eJ4���a�Ȝq���$�+ �/'�������%/Շ9���xx��{DJ�S�Q�;%����O��+�])�,4�T���3�̱L�1�;|��`*I0y,�6�;�u�x�zƝ����fͶR4}���у���ϐx�dۿ�D�M)���-I�:������4�}�S\ӑ�%�~Er��K���]@�l��W[�,_��4[�����L�g��e����ަA�g
�]�K�:}[=���>���h
f{�~,�Uz��j2��l��]��l�F���s@yR�t?t5��~0[���.�*ﺆH�4�ý8��)�F�ˁ�_�b�AϫX�#��o#0�]�a������A�[^{S�s� ����ݓ΂UZ�����[7�h�91�B�g˫~��e�6�fn��?X�D8n����E_OnyGL�{����P���\�ʼ��� �e�
W1� 'uܩ����mX��9Q�bB�ܘ����܍W0r�l}Φ���/u�l+���)�n�\���}
+>ڱ��Bm��p{a������2��bAa?�@�D�
�%� t�2UA��N[�Ԉr.$����~.��-��h���[�h�yU�ظ�ϳ�Mt�c���B���y��a-��~(�����Ąe^˫X<{�D$��Q���~���`m��Eik���U���Ce�� �%�6��G�r�����;��ɥk�-�[A%נjktC$ĝ��<�HJ�{�nQ�0}"��&\eO���3� �w�	ˍG�Yn�>��{��j�K �eMƌ�Yi�� �mՑ�G�K�9�jwR�x�e4�;R��kc(h�r�Y㽳�T�܋��0����S�N[i�yx�ISmb܏�-}����<Qt+/��Fnɿшv�v
IU'�D���4=���I�&��rۭ�u��D��|g�m�-{n���a�lU
�!mM1���Uz�D�Qh��04nw�3�}�8��3��GU�����eiyfz{�گC. ��z�Q*�A$�����`{($��2��n�d���V�?�.���亅U�bB��~�8͕�d�o�tP�O��n��5kskM?��t[������ �|���zQ�Ʌ�Wv ��c�+�扡 RH>T˩u�E�}u���7`����>l�l�ݚ��)xBF�$�;�Co���9�:2����~XM�	��.����w�8h����Z	�Ex��"*̛�qI�c�+��89���_|aG/�ۂ��e+�f��-i%��o=nmx�X����+_wd��h�x7"iH^�x�$�|;x�䗷���!P8-�q���Co��F�� -��	L�vm��<�o����P��[
v$���S��m�s�v[����!F��4�%��wx#������l�AɸR�,:���K����
��d�X=�#�UJ���(���I|`�_V)5e��bBfJ1��gỸ���j�9��uˬ�⍱��I�7TK �3�VP�dǊTzz���h�����N�:Z{3�[ �v=dL�$2^�)]��Ŵ/�@>�ٲQcm�=�.KY���x����������e�%��t-�]�l��:���$���q�s�1g} �2��}c�䋤��|��L�V8G���
�� ����yƈqF��$��I(�Q��i��z�r�����T���eY��N-�6Y�P��[�?뗔�P�MЋP��ȍ!t�aO6�#<�SܹbH�p�H�9W�	�o��p\��7<۪(���Ah8�(�"&C<E,�T�hܮ�=/w���m�NF�N�Ź/�POGlJ-^��-��5�v2���)���:����'�ؑ��jx=ωE����[d���4!&]��}��8�ӹ��E��9��L⵷�����o՞oL^���3aB�E_D�A#�{.na��>0V��]���ÊY������=���� ���TV��\���:���kl� ���|;�P
�h�����G�"���Aק�/�&V�⻏�b�_���*�*=���`3��tu}���+�������'��W�*Ki��e-�,(Ec(���� {��Ę&0��t3@3}�A>���d��K@ٲ�= F�T=<�#:�t�K9$��kV$Q
&z���kv�&���H����@��>��{}�@��P��
fD v���$������a%�\/�� AL�WV�zh7P��R�&L�@QhjJ��8
mG�۝��I���l"���!�3�)�o�%x�ت��p& ���/>GB`����_U� �W-�3�����!�>%�.�_��D��zENTu��ά��@���)JՀ]�����S@�~��z�)�M�ϱR�%-�`�z�<r��j9�>�0� vS�s���#��}4��Qm��9�C��y�^��7�O	�����!3�Ԙ#���Uq��ɺ�f�1AnB]�,����)77*U�����3;��F�ˋm�㗲�|�U��ݢqO=_�?V��{!9�I>�EZ�A���EZҴ�ݙ�3�Ad/W�����r�6K;N8�7,Q�G�n�l���� w|��׋�Q�����1鄕���ƶ��pp���_*�Y�u����m������3��O�d8�xV
�aA�!�1\��r�M�!'5�W~4�$�N��$���Ł�lz.�u%Z�����9�>�k�`3���1z�ɇ�C�̂}@����m�eiu���q�+�yL�'��V5}����`�X�#�=�q��#���T�$@-*s�	t�*�^����m =[�Ź�*g �f��!<D	��� J%�ZL���G۠W�Z��	MN*�sݫNd����kW����h�(榽���l���]�c��N���p��E��z�33|��/BH����B�&A�>`�O|][b������s����W��*�������IĠ�H��r��0!zwB���9@y��";Ï���W�W?:�%�6Wkwz�[!�H�lIU�@���, ��Dm�a���"�[%f;�kf��M+��-�Ώ��f���F�y���� �K��u/4��,�xg	z2��E }�1�(@R]fK:���#��e�P�g�-la �0��f�P�FA=��<LC�.���%�ZF]�H�e�x
��P����y2Bc�I�(nӪ���*��j�&�ZZKQ]ɶ	O���ʃ���(}�Xv��i퉰q����y}�E/t�w��k��$S��̇�Y�܀
�R�9�F<gd�R�TJ�߇T+)R�ot�I�BZh^�Zv�K��Iڮ�͎�}��)��J/�$���&/%q>�r�+%�ߎ<���G�S��6�y$�3sԎ�Cɖ�B�m�?v�d�k�"Ib�s<ߪ�(*I]�!]��G����3_�r�i�pË.Mv�@ܱx"z��4yÎE������Cd�.�8D� 1Cf�}�x�ۍ�<�Ȍ��Y��>�Z��**Q��6Ƙ�l�N�@�\�b>��� ��-�[p����N��̪��&
&�ġUC�*c>!A>����-�|���;��vjGl�{7�1q	9P-���������`pZ�Ч��H�z�}�����p��ڤіB���Ѐ̿]��yW	㳡��r�����qm#�iM����e�\���3�1��	m$�6�R�{g?䏟�m/[�5Q���*��W�&Ю��L�W��:d���V�?0� �xڜ��:��"�$�|�M���\�/&�}���g��[)��F%�p������@�D� �^%%��|�Ѹ�`}Rsv�uM�)��軏c���si�偠��`�4�c���T)U�u�e�6��a���L�n|Y�3�e��P���p[�NZF�4E�#V��$eI�3�^5�VP(�iy���~��`�YO���|���/\��@Ƿ����5v�68�,�C�(*}����1nh7Mu�Έ���å��J4 z�.t�c�9_�RrWp��WW��,������SZ�iѨ8R�s���>��[-~��/m�����B�?J�{�d�ɧ1
��gG��3B�����X[�ۛUacunGe8y{3�'��'ͯĺERs��^�K�-ßa�Q]�诶
��&nv�Ϥ��#���Zi�_2l܉���L�\E7Ԋ�,r��)�
�0����RG�9"�ѱZ:F�>���?E��W��u2�0�l���T�$$|�7_|���q輖���x��d�1�'!�����8L}p�Wuvj�w:�� }x�ڷ�D;�=�$Mב�����p�rw�Y��v]���Bk~2^s�G�����}�ޟ÷���HNo�E�)y�N:��� d��RG@�M�0��c���YE-{�0�6{�����9g�M1�,q2��B��~�|K��$�~�H�o�;q�:��%�G��a�l�p8#�J���D��o&k+�r+��g��.���vӪL��J���-'��}>�xtX�l�mFL��i��S�1m��8Hf�G�������E�_K�n*�ѩ�I���<���g��D�����j��8�i"��GX�����'V7/#x�����Q�]C:�#�B�4j<�4庹�6
�S	�f=ns��/�ݔ��Z^�\��`i$jݿ�t��-낶W8p )y#��h���L!�5�,��y+�ުCۡo�6����p���%o����c�Ok�@�d)����F�q���" zp������<|��Ȋ/���*`�VI�\N��`�������s%]�:{O�ꕥ�F)ഄ�]1jy��ǋ��0�X7��Q��pp��4�Ğ�>�J>,r!B�ɐِ�E���0�!�g�5g�T6���.n��ٺ����|���Bi�O����/hV�&�*���ؐ��mHw�\ƴ@]UX�����\����C�O	a�J4_So'�W6����T������ѡ��p�Q]���%���lV�B�<c�����8��q�*�z�_[���)���.��?�d��������8Oc�^����a��Ǭ�G�v�^ؿ�d�|;�i{ً��fOl�v����؅9���Ѣ�T�K|���������7i�W�o$&���˻C��6�i� %�p1�i��|�3f���,`u5��v�gI�/�f.�E��0�}�Z��( �o��_�.�'Fh��Uh�� ��
�Qb�7� ��AU6���_Av�߉b��R����^����/Ū��Z�
,��|҉��W�5|�"+�Ɉ"��pNIB�H>-�D��`�Ub24�����\�cBA������\+��*�\f ���[Ϩ��F"e�&3h��b���~�+��D+V/��v�!WV�wq�,���iU>��<�7{۠�2�pr��rMX&����j�T����f�#v����mt^��qeU����1�*}V0eVhb�y������FX�jA�ǚ[	�ȕp�#�(��$�}'B�`����#�~����̪o����_�dK)��B%�k����)��̕��u�+��AEV�y'e�ɷY~����a��T��S's{��z���(7�� ��@q3��h�����%P�ð�����\��\ޱ���x�֘�XPq�;L���7�LL�J#Y8�/��S��TuB�<�{1!8��B��L����I�������aj�';k7�q;$�BVF�x'����UT�dm�8s<#�<�����<�st.�J>/|�_��($��a���N�z~��`�%�_�橎�E%|��P�$]~���\�ݥ���Z�04�h���ގ���z��^���$���6x���g�j�5_�)>3|��/)���Y��x�|*�'�%V����gI�y�:\��Nm ��{hg��@��\0y�§W�h> ��>��UU4�fYWF$7�b�׻��tEQkwqU;�x��n\[Nh�OEǵ*u0(��lP%��>PiI����`O����rŗ���G,a����v_^KAm���'T�1���ǅ�
���´g�c "@�1�e%c@+�Ȭ��8���F�ϣ�⨋��A"R��mF���ILL"W��i�#�*�Vg%_.���uSևq8�A���o�s�f��5�c-�QL����D6 w|W=��Wf�+���=��YT1�l}��>{N��1|Z/���o�6NylŅ�@����:|$���g��2�����d@�o���>�v.Y9K_�GQ�M\F]�aX,� �,����^��x�X]M���+�{��~�3J/0�)�T��i`�B�QK����u��Ǆ���t??��H��Og�E{|����e
]��+��$d�m��c�M�w��H��e� xӳ�P9~#e��ՃZ��a5�f�5�b�d�m��~̝[R"�X#�3y�	�cq/���K`|���|
�l�`���?]&Ѣ'J�b�kp��ɖ#�	.-܈����j�d`��`�$��M�l�)X��r%�Q&���q�ƣ����{�����S���f�]������ч���}�,���2y���֘
�^<�DZ���E��������S�$�8���Oc��������?��%4ҏ����'H_���j�C"\���|I�WYZ�[$��Q��6��XW����Sw`eU�ə8g��6D�g��:����}��~����K�A�O%z��Z�:��E@����csJ~V1�dƫ��kx���Sbe��?g9�$^�YD>#�r��%���H�l���9�H6�߮�^G��d��=<����C����	��m�zi��?C��>��v� DQ�xQ7P�U�aH�I���!?����J��t�����g~݋����gS_$�B�zu �� �"-9��{oy`�H��2e�u[b{��;����/P�N�ab"v�x����D�u��'/�W;a��1��r����И�ϳo-#�z"�dN���>�8 ����Ղg=�ϿL:T�-K�n�e3��Љ�PY��s"����.e������ͪ�����"t�ؤ�e�)ـ���Ɇ3�Mum���>	AX�d	.�%��?W2n��4����K·���T�ORA��2�^�JPj:��O���"> !����j�P�/�0�NYMBԇ��@�p������`�O7�, ��D 暍�g��VS��J}#t^4%o׺���l[n��e��~m�T����ƚ�"m�6�4�����8��8��Y�5���=�l��s�R��n�k�v9�l�e|�Ӥ,ZEjn��o�˖a�N8����$�_��}���~~�]Ƅ�KBH����"�̾�=8���!.��;��Ϡ�� ]�`s-���9q�i�"�s���]'����7�`�	���7?�J��?`���<��6���A��yy�Z��n�?���Ο3�D�;nQ�c�����l]Ē�8dpＳ���_,�	�3��c�L�)Eh�)����5x�!�	�ٵ�_��6.V��o6��X�����/D4!6q3N|PXƸb��4�M�[�8��ߞQ��Ұ4�~����4tA���V���Y��tPn6���l�h`�/\�鳒?�v���n-���Oo�"����d�tZ��oy��`������`�O��3%lQu�<r���'1�A� c��X��O�Gi��'��d�8�W�nt�kI�f��M�(�,#8�mፀPX�_���ؿ���X=��U��S&S+�ҏ�ֽ�W��zy��ރc�@R���Hbt��"��Z�6����H¦ R+h��θI�r��AwK���%��k��w�}L}�0Röv�@'���`�O�,��Y��i�������	<�-�Y~�k��c�������I�f^�m��^�C{p(��<c��3�w��L��0|��@X�-O�&��ח
6D��V3^ӮH��&{��?�yڡ����V]�v���j;���/	a6���{�qJ[H���"������~C��'0�Γ� ]�i��}�E��1��`"M���w����Ӄ������)^f����������w%n+ܲQ&��S��*f�k%#9�(�����־�O��W{:��q5^iHk7�H���'#vn��9L�\:�P��f�u��U�$$P�
�&����|�E����ԩ��R��;�ň@���$���
�\KS햑�S�ƹ��b"k�a�������������+�4}�.��9=����t0��^k��������>d�7	B��X���p}c�H�ZӡoNm������q�:Lϒ����~l�V*��(�A������Ą��)�Ɗ_k������߻����@���+��D��ٔ���2�(�y$��c�g�T���G�$���s��nN���-&��F�Z�_�ehN��)�W���mw̖�Ѧ���� $�*��(]�Q� *����G�M*6����v�m猚���W�4��Gs��
z_�÷|SÝm�Pj\��5��N��J=��o%� {E�QXBgb���Z�m�M�fuW�S�b�y'_��}I�32�βx�c�$ě69�G�[�
9g�NZ�/v�J�8���	O*
�P-���OÔ V�e]�����K&�9H�E/�-OW�{��PY$9���Ʊ�l�S��Ȟ�Ze���>!�'�gt(M$]�>���#��L��>���Y����[�~%�d�0�NQ�	�k��=5�����|�^��գE����<�aNK��_G�L\�.�MT}�g-�\��cngɃS����`�}k:����sn[k�&,��cc��(��5>g���g�"�ܠ��	�2VVM�R�����t8��@*^�x�6܄Ay��-m�Ʊ#�!%����glEF�f��NuL�i6���p��WH�wH� b���+�PGA|H�cs@�g���9�,>��1a�ܔ�`+uo/UF�:�����y|Qs{x�눹�ZQU-���^��:ܪW�<���{���P�;��cc�w����r�i�==�&T�bjkҎ[�2��8����1�9n4v��;ð�mz����+�e֕l�xu7;k��=�$���=ܖpz���s�dx�~u6
����8��:V�U�u��H�!�Fj܂�513{�iS�����PA����x@F������J�s���"��(u�<od���J)�>B&;3]���J懡a�U��>��bfVtL3l.)Ou �q$>���l���������mG��-K(_(Ƹ|Q���N�^�Lt(���"�q{w�8ӡ��d/�Ӵ}����S�on��¾1/l��􊑮�3��k����}�Ī��-l��|0�]�G��WϜ^+�R�g�yX��ʦ�"�绌���9��)Uhw/������w��?�f����.�j�ωC����R�\w�O�Hx��)�|��-�eAp�����U��#��eS?�)O�A�&�!o�JG�d���`�6�n*]�6a��������:��C�<�N�'4��F��� S�@t0O�w�s���h�f�H�;@1�f��
W�����MA�d�1@=6j���x�Z�i�����)z-�B6>���k]#u܈{S��L�iak�� 1�%Z-,q�*+��-������Q1'�[䃗l�f��[�z�$��[�1�֣����ح���O�u���0��|��n;X�Ar��/��G@+�K��{u�<3�x�HW	�y�o~k��tp�oGֿ��A����?�p�Sc��볃.10�/����t�z?gJG���~;�����mNJS�w:�hX-��3K%��M���`�l
�,�W��j#˗����W��z�������h0��i�Ē�Z��l@�D)�\@:1�w��0Zg7U�Z�M*�T���rW?h�!��:���b����%�2�2����r?��$��bH�%��)ݿ���\R!ܖ��"��Sa���}�����3k��M-/�����W��O�d�-ݯ<-pI��n��M�"Uh�H	H��pap	J�lqs����E�Gdx��L�ݿ��`-�&�
7��*0#r����J�# o��/&�����*bxD+����L?��:2/H�q�&�#z���o(q���Q���3��"Rp�]\~a�4`��#�v<��]�p���u����n��y5�[BhTf(��^j;F�J�����;�=T�K�y���i'tܑ6K��mi���a2�7�z�+���"=�4�|62ա<�H�UĬ��o�+?K�s��-��%́��=�S��<�"��D��`l:�@Z)��3����z��h���R�1�l,C��G��քQ���8�P�_ӪFMs��k]�R$ڞ:C�"�p$�Lʴ�6 R�*�J�m�]aq���^K9�H�W춚�OUf��k�ȓ~+�8*����&}:�\ޘ�J�E�A=�.b?)�<?��gw,�PI��@�?�}��}X��'�;��gxR|��[�Աy}��X#��Y/�ミ�!�(��ed%�����7��ɜ�Z�) %P��!ӯ�
ZM�Wt0�i�!�1�a�.�BI�aC _��V�!�T���M4z�e��e����^e<�{���*��#��K}r?ʀ�+�s�0g~;�	n����L˒�-���u���t2�"����5$;�x�I�T�9&.{�W�y�7��9M��Mؽ��I��N�g���3r,�Ǖf�=�4�Q+����_�1n��g���%����'���f|�[���Sκ��hkrsCmh�_�<�CjNj��~��d8�s���ڣ.��j:TU�z+��tgx��"F�؊\�'���֫��HQ�Sn����6������D����)�kۢ�.!��q�=N�7��㨣��_O�Z�������V�����jw9�A�W��GL�Kn&����c�3h$�+�_���n�4 ���b�TW�y�j�
�+�}�
�N�%g�D6z�ϳ��b�͕w+����C$Ԋ�ȼvOp�Z&t�����.�ׂ�\V`��-�d����/�N��b49�Z��r���Z��f�Z�FD�<f���m,�Um�.����2zHFK�Ȝ�r�qF���A�kc�,�_ α%U�V�&�8m���E���V���W��m����S�������7%����@�u�r�5�o&��������!I��d�z>Ȳ�z�Cf���c`�X�P������<�e�����7�DaD�w�..p����=a ��:(�E�v�H��C�)�3��E�t�|��<�{��_�o�2K57�W,NL5�jr���d2�KCW���$��*�YW�ʜi�1��q&��.���_���>EN���T�
1E	�`�# ��a�Ѡ���&㡇S�c�ʃ�|erY�s��C&��d��-C��'�|����KY�����BNù��ƚ�k^@��f�r���(#c��"��p���&09���R1�Ai�e���f�[�|Wt{iy� ��ה�0 i�<jŶ"���v��:��JW�9#�@ևA�ѵB��Js1����,(�~1�׎_�[ ٶ8�WhQ����~H��<ӭ��/#v0��\aJ9�V�Dk�b7�S>��� K��u���\X��h.���o�Ѥ%t���ۻ��䯪�������NyZ�!B�9<>5�]됡�̰%X����~�i�~�Yo�8��;(�(	����c��Z���aXzw�E��=(f\.��u68o��0���{+T�p� �הA���4�i>�@,R^�I�-�
a
��g㯃�+��6d��On3��sÆ?�F�	�]B�2�4I���*e�H���v���cͱ�q'
?j��ҒK�;�%jvl�ܚ��7�Eh��nKC8�\y�N�k��(�1�r#Yf�S�0�'��g��DFό[6Ny,�1n���.�40M�7�e����?m�>�l�Ć����d�G�5KA�#!��v��L��Tr�t�r��K��
wN��z�<&%_)�=6e�Xk٨�#�/�������τ��o�yNE�&�� ���[he�?�}�92�ѐ�M-1��� O�2z42�l�BRY�_���h�j���G�j��̀��(����t�29l+�}^"���[xv��:)�È��ѵ|pyc�6��f�V<û����"���p�x�z�#��"�� *�g<��+�qρI)�[05Ef&r��N��ۄo��~������@R�N�IR��*!������q�bvj����L����^����B���h}=п
q3T�w�fE~�^�Z���kN�O�L�8u/9T�	�DbK��c�����E�����s����=��M0��װ"��P ��0�!�z<ȵ��`G�R���H�Q)�YhC`,����?y��ӗ{��חq9-?�T���n���cY�_CT6��k-΃�T��6M�m2�Jr4K�Ō �7j��0AZ}������fq�e�jcTnt�Vp�J��(�g����j�����)r���8C��1	�U�s4�TW�0�@�^D09�j�#���=9L���@h \�q|�Χũ� 8��W~ '����p�� Aґ�3U~�(��x!J��:;H�֎v��W�-*���l�7��"{�㜣�1�^�:0�\3[eG1�#>��vnmF|q��g��Z�m[��H_��װ뛃����F#�T((�u��ÿA���^�)t��lX�#���s�g�Bj'U|��b��͑�UJ�v���3�X<ߣ��s��{��Q�e��rP�^ZgE��/l!���[�4���Õ稹�3MZ�@lk3!ѡ�[���_e��ϻ�R������G_������4���I��|�[�(�x��	<�f�:�̎6<i>�;����=����]L�^�>a���Ff�J���L�|-V�����,������;��
� ��g�I�Lc�驏��K���6�ù�0�Pі_:�������β�b8�S}�/�6�+�9�� ���+�)�o�^�x�7��D2�^b[![d�xyPN$H���OR��'�t��X�;�}մ�h����"���G1�m觐��`�xp;��-_�"��Pȹ)V]|88�eN�r��U\�w`U��.Z4u?cˇ�\���"���&'*���ݖ3f�^)�l$��	D%�Zc���/k�/�$Lߣ�&��&¡�]�� w����:"$�ۥ�t��4�[��ǀ�jSw�<��2:u\v�Gp� �in�%z/~��:sA�g�ygH�;���k�<A@j ��|��vZĳX���n�����9۫�+8Vn�R@z���JE�S럩12�d���-db���í��f廙�9C3�aǳI/�XKB��vr_ WW N����eV9CmHw
��<C=��N����c�)����{C$?���f
��-����1�,><W"��Ѓ�]�y��/�1�g�֤��7�QaU��E7
��T�]誋Ug�f�"���g�&(0#��o� r9m��E& GgG��	X��$�]�����������������a� E��n�^��71�.q��aoսΉ��A(�^�7�+h7ł�$!R��n�ś� p���9�6^A1ޞ���B�~���^��ؗ���708F��iy�WFd�R
�o�(�Z���I�L1�|���dJ�N*�ׇ�pVp[���P)ծmƢ��*�CI\{:zŻ&Y�3����k"�%�~����|{�&8^���([��o��t�����a'"r)��#�^�H ��i���b93ͧ9����ĳwYB/0��gҌ��B���Á�����: Ǎ�Ki��P����2�V�$؂+�s��,x�Q;�R���q{F9_��969���${GV7F�ʛD��+|�����y�҅�2��	�����y��>d&�Z�J�,�eC�;)��Eߟ�u�TI����F̱zس��R~8䋱#ћ%�V�e�b���^̣e���-�s�YI;i�6�D�:��Q	f��&��EQs,��%���"?>�E1����ֻ�i\��
�W��И��O�$�T�Hn���3���8�79���&Q\Qc��wxP����꾧�!*T���q$n��́��K(�D~Ͷ�����џ��?���@78r3G�K*��c[7��T��	�؂w��md��d�8W�R�y��{�i��T���
R>��u�6��O�99F�]5�$ṽ�x\M�E 0��k�����
L��P�$@t�ɩor�>p�UD��_�x�6ŸHfw*��`lX�5��B�&g���?2]��?Z����"��ry`b�v
�(��*�o���m˅&UZ���w��������+82o߬���?�ԃ� v����b?�L2�3����e�.�?7:=q=W�߮���k:u�!�<E��OfŘwK�7��iJ��2*�4+װ/y�`��Τ[C��y~#W���1[�Ԭ����)�gVcVz��Qgk!��аH.�a��R��\�<q,��u	���7Ѽ�0&n�>F�*`/�L�O���O��8�+,޷+��;��y3�� U8��v�f�*5sQ�f�'��L���Db�_��d>��#��}��-�J�9���]��ҀV�Ɗ��鉕>SД��=%����y�1`��	�V	wL&5)v�v
��'��Tw�#&v�����n,�8=�I�copj[f�n�6���hʠQ@�י,�6QH101"�}n�o)����֖�I�X Q\N��I��>��܅�lPX5[h�����bR5�m��q�|YYυ?H���S��*ȉ�w�xPm��;Y�G����qX�Ή�YW�4��9﷕l���g6�MW;����`�pA�N!;&JaS��a���逐rQ�tęyX��Z0?Kj6�<�[�|���2�񘳂���@�D��5�;��)�80br1@f�AYoy��ܖ�Ȗ*�f��3�Hid����U�n�D�3���{} ,�@Ͼ�N�{ƞ[D����X�g
#U2))W}�C��ߐ?d���2BP���a2�Z��Ԙ�'�V�\v+غ�1q\G�N��ܴ���Z/vί���,Wz��G��ٝ�z]��ԯ�.�>�:�l���rd]Y�t�������X�7���Ww mc+�u��m�V/C+=T�^�<���ՈnW᷻,���"�Q�:��C�FM\�R���6�N�X�L�>�z4fٱ�����/�X$����?Tuz�0��YDWJG�O��ܹRe�͕%�xI9�_ɗײ������{Fޗjk;8�bq����pEo,V�Kdlџ�v�;�<��LB�s�w1yEb�����k�FW���1v�ćZ�/��'�c�&�����)��8���s�
�m��z��zvW���ԅi�Z��De�aT�l2�䄕p�J`K*�����w ���q�|�O�1j�����l��Y��8��;���G�@rã{}e#-�� >Q� y��^7;�k,�@�&���%�@�!����e�+v_�`�Q�E�L�#�M��D�afa���)y.����󍂒 ��g�ح���S��|L�N%s)�į�{w��0��ܵ�h���w�=q�mO�Lh&pi	:�N�2Q��E���ngC����
�
��D�Ŋ(	1s�媛Ijue�♇q�7鵮M\w��I�y;�QpLz̤;�$E�AQ�_y�)�Ѻl��1���� �h#F*s,������qXc��l���'U�����yƍ=JC�B"&����N�/~�2�Z���Ga���4wrOW�>�h��%�>��[��zڌ��Ԙ	0����Y����T�}|�dA�O�MwKi�T�/|�S�Δ���~��zZ��ܹq.vw��9��.~�)�t��<K�v^"�R�$@P��f! O`���A�/�h���g{�c�pEn���d�>VM'ѳ�Ͽw��7���5
l�LZe��Ƒ� K'��&$ ��j}�/(��h-�_<�G���9���/��k^Z���%!M��7āL�)-& �11��� � h�)g��4�����E�{�::�+ni��?�{G�Q.X�aS=��N6���e��,T���Y�hzF,z7�d���E|�7W�$g������)h;d�^��2W���������K��t�W�*���z�k�5�PgG����UZ\���j�%�Έ�@������~ŷ�Y���m\)�CT[.j�N�^��F���7����	�\�t�Q�i1%�Q�%���Z��c��Ԍ���6鎃��,q��~��QA?,d���4�1x?%ʈ��T�q]&)�Y��"�y���*�r���@���NW,�r7^�Rϗ$�o[��$���Lt���` T��� �2h����D�Vg��ڦ��|��Sl\)�ǶxyW2��� s�I����^K��N.�lj3�L�R-�.��*	����+���R�{0A\��o޽p[
(�!%#=��RU+�<O��- "��|J��KL��uQI�(�vu���R�xuТL�uj�����y�D`��Eh�AG���S'��pA��qd��X_+����B/9[�'���a�3t� �S��(�Npr��BQ�s:ՃІ����j��9p����Ϊ1�G뜇R�ݍNJ�@Gu�d�Y=)���-w]�@ uJ�$2�LGO�g���~J��	�o��9�A��Ѧ����0�6��X�8C�]��KO�C���G4�:�ȓ��s��]Gr«���:��F���'�Lj��S�!�U������1��G���/0\\A=@�́��!F=24˔[���������>����8KkǭR�aSq��섕&�u��2�T.�����f#�JYU��c�G��%�5v
ב����rd^K,W��D��w�p��o��*���#��U�����r���\���P/ߩ/CY�Zؠ�����j�+ssX��~|�cU���lX����+v��3�d��%ѣ��O��Yk��+&Ω����m�� �D�k��/�5ƴ�&o���(u\iBAfA*]�X��i}r{9�g5�uGj�\hJZ���+��� N	���w��[�����Xdn#�`AM�L�O�9�hTi��"�����(R��t����/�}y�}fÁ�$X�X2��N8"���+K�6-Q:2�D����<���+�M�k���މ\���גR�1,v�o��K�������� #T��ㆪ�1�F����a��s06��OX���؃o�L�9�ۙ�;��KE��K[jގ�����v��(}����M��W$XN��Pq;KQ�C9./�&Ň��eBR���"�*���pv�zO��%	�v�����	� ��EER��[-Q[N�p�>���-z�j�{�0	&���l�������m&�_-�ֵ^�MN��k�x�vj��'>,��ҷ��\�*���.�Zf$�c�1�63�^�w�gl���^��q�����]-�2a�8�?J-�'qAA�����3�ܹV��EJ��`$q��!�
~K)m� ���~���#t��|�gWsR!�5%"�Z���c�ɐ3h�M��מ��k�ձX�u����1��fo;�a)G��h'����;;�Eç.���C �l����-�9~��7�Ye���N�o2�K�ul6�CX߷@��d�w-L2���WY��������W�s�����վ��+(N��/ބ���G_����Z��%�&�@'	W˼�D2��4��T2+b� l��p�\���:���u�b٫7��@����ǀR�T+���T#�K�`8�&��h?�aNvAu6żt�;�=�����t1T�:����H�tY�zd�nϐ��~��I;�1E�D����0�.s��P��ۻg-\��@~��	9���]\���A����$����e�W�a�\h��� Q߼���a�t��;皃L�<s��nm��� E���n��ںcu����x�VM�y�>͢����IHJ����Xk��H;
����H3U{�S��}�L�4�8���,�t�}�
 �W�ǭS6��a=r�v�k��ԭ-	?�d�����L���r
��ݏ��B�������� ���(P��~!W2e Z���qj��ۀ�B΅X23��T9[r��AD{X��DV�}A�s ��ˍ�O轝1�Su!�=t�Ō�}�7"�-E
�E��gp�:�"���W�V2�HtF	�7\e�]d���|�Җ�h*��������7���;�9��5򋲰��ܷa3s �r��hT_��ۻ&M��!¾R�|+���n/潧;�^T����i�>ןf{�_�-����Ҥ�i��%���춌˳��$�I �tx��פ��ջ�O��9wA���P���MH�n����lkB�&���*��Dn�ƪǽ��������X訔��"*R�����XH��wip,RG^4�/��q���`"����ɫN���Ώ��@X�$�֥� -�E|w�H�L��ks��W�M��`���Q�D�m��K:��?2�C�@�ţ.�I�Zڻx��(%mgDRFdd�mz=`w�E�¾�Ge��h�~��C�\��i�F)��z�D�H�i�l<�b��Àdr����d���@+N�\���)_MS��[���b�_��$1�:�
�
��5�]  &���zݔ�7V���j��b�K.�Qk�:%e���V�����i������[�4�%	w�0�d�C 2�I˸f�ᘺ�В;�Bnΐ/���O��+�G%�Qׂ����'�fG)��ņ)�+��/<l�%��!k�υ� 	�}�N�j�i�����Ͳ��/x�"��9�q'kk��Ι{��X�1Ǫ~+h�-|;f�����֐��ּ%�j�:Sv��MN�>0�v��d�8�W�/��h�@{���r��J�3ϓ�4��Dk���2O�Ѓ�dZ��]d���/�b�{I���RL�ldq5@=v_�qV���۸����d`�����ꦻ�)ز��ÿ��JC:��S�6l8�Y�c� �=�#_x�%�N�(}�˻��|q��ܺϧ�w��}�Y���9Ċn_�g5S�p;��q�uϚ=���w�|�n�ս�@^�RzN�4�D�o�o�"����>z)Aq�<�Oi-<j0l�U�:o��k�I�������DX�i��/#�����*kM�#YGj�b�����);tP{�ʠUr��s;I�>�)�fM�p�T^Y�犪�M�^f��j��Ӫ�xS<���z�@���VY/����� �;���:��%k�h�z4���û[(�C<IW�g.�Z�ZJ����_2�2�Vް���ʘ�"h�&�Q� � �vz��b0�� �t�a�����[b��z5����S�9�%�Z�z�֕F�=k����G\F1S��I��?�N���9�L��k�){�9C�p��(�Lǣ��&ڄ`*��/S_���k��m$d��}NT�`#g�����F�*8&$J����`�[|��Q������>�����2���k����|b�1����C9�Ι���c�yZ _M/.:�{s�r���F����hbB����x=�P~��'3��|�G��B'�S;�"��ee�u��$F��P�ƪ���+;R��ė�,��E�G�%,m����C�g��J�ӥ�a M�����h[iϢF�,��0n�������oԸQ��F\��j�TQ���L����1辑k��]L�.)�9u��D�# 6V4�y+��4��f��p�%���{}�C�7XD>3��IZ�x�ܽ��n|�.Xy�g�� �㴣��a� C����%q(�k�PX{��ގ	מ�����M�\P��Y�g�!��Ͽ����l�}�?Ħ�锚�� :z�css����VT�Hc��R��������K��_�UA����+���1�5��ݪ�u+|�x$��{����9M��D !]W��e�z� �HSg���������*Q�A+8��*��:�[H0׹S�zH��x#,�n��)8�W��:�%��d�W'�c����t�,<ડ�e���K�Ҩ��A8V�m8[�l��m���m :����Q��B��>}�@�QvX��[&z�#=g�%��:I����d)f틛tJƱq�� r�mtр|H�q�%�+Y�̈F8h�h���N��B�2���
y�2��0گ.�68��B�{�
O%A����R�U��ۼ�H��O-2$�E�Nb����z׿�#����$>VFp*^[��sr;U�T�ɨ�S��T�'ɠղ[<�U�#��fG�y�.�v`VY�>��#�O��.tQ;S�ln�Kh!��B���B�;�fX��9+�d���ڒ��a~�!�^t���N�6��qcQ�v�5E�}[y,�J�;c�x[j�PQ0��P�@�~���@���ۃ���t��rV3d?K/	�f�|��8�m	�vc?�qQL�J�v���~�g�G�V��D�'��I���x���ZG>������vS�iZ"�v�M)`4������"�x���q���=��h� �B�JU����
�4��f��Au�e��}ӧY��O��"0��K�	{c���}���:b%�R��55�~_.~�H�l�[��Ã�ڍ<��.6�#� �������rRB��X!Po�l�O����H�	Uy:�)ҥv��S��o�aa�∈��9�NF�"B�MK~�Z���}��1�=.,XɱY���o/��)�;�e��_1ӭ��>o���Hl���c����?�9�҈~��&h��\��1����=�Q��$��\o��!����r��y).���j���(E�i~�~I��&�	 �.w����������	9]�p� ��lZ����L��QN����Q��V���Y��Ţt�-Y���"M�A���{��7�-��v�L�j;>t0UΝX�_|GNs�p��(sa���-%/Q�{�*�|��3��� � ��FXp���oʑsh-��u
n���ɽ��
����}7��T^Qm�g�l�>.��5�
n��x�i�����ڣmcE�.P�>c�7�3��V6�Qh��)�TS;WptF�kN���0�H�gI�b_���(�J��ou�T�8k�x�������u�0�vNb"�l�R��kkC3�.]~>;�;��Ţ�ǜ^���|����_�� �y�� ���W�7C`��#�/�݆��b|;Ǒ�1��X"8�]8���ޛ� ͗y	��I���yrH\�h����(�6�=�<h��~v���=h�&�ݹo3�j���i�Y��r����p-+qy�����"�[!�L�(='�Uh��[�Uj3��4у$����
��U��J
䇳�46�?j��qrc���K	W�u̓�Me_�Ǳƍs#z��`m�sP��>z�&��c��B@j�N0Y��
���el������ �����������z��Ÿa���ˢMrH�G���_��׬q�G�����-�V�l�o-�]�.ǥa���ƾ�텊"ŗq�%�{1�w�mQ�(�o �Q�;��O
iD�<d}��Wq���K�s2��� ������֣����&�m�a��%���"Y����a����^�#�������ʹ��BJSU(z�����#�;�+�'WѾ;�7k�����P��A<5ɲ\VwR���ʉ��u �l<�WR6Ѿ��i!�M�5`'�ԡZ�}��O��f�,z��{�jS4�Sy%I�RjD�,�bV���m��\D{��� �#����9�Imd2��iW�V��B���{�F�gŭ��ts�<��Ј�S�T�V�<_O�/�*s2C�h-�-��l���3e�Ri)��]���B
�ͭ�+e��W	Fc�Ia�,��6�YC����K�ħ(��s'\x�C1]ۄq���f"b��Ms�eO~ƺUk10Q��O������Co���Ȼ���<l���~��٩迾#��>GQ�Q�E�b]��/Ta�@h��WY�Qѱߘ��_Ԗ6d�p=p��c
ۀ��`�r[�M��
ݩ[�3�Nl����e��+2���C@�����m�)z`�9V��屣[�V��>"��-�zO�,q?ܭ/Yr{��������mS{�"�[�f$��U�-V��:++�������#�B�60�/�Wt��*��O��n�`5!�M|ٱ
iv.�uX/����Ň0F/?�1���D*��J��ơ�y�����6�mS1BWxi[�`X�I��Ջ	�^h��A��PN�?rH_0�s��늽!�LX&������]\M�2PĊ��x[\��e7z_L���=��Cv�(�6�����}~�S%N�-i�Q���B����;"5~�#i�����S�Y?s��&�+�X�Kf�j��|�(��x�d��#� �&���B�|��з�L7����t����>�w���o,7+�U��w�����$���t����x�:����˪�c��3ׯM}�>�T��jxmW����<e.�:��^��~��E��F�Kl���̃�◴�E���cM
��68�BV�R�����fh4Tw��>H��.~@�v��3p�&�M��n�о��V2�RO�>�vy>	�*4�s�_��A��������Y+�� 3#�o˂؍�~1��n����"FˋDv����}|-��*�JG��d��٪V4�{�������E�{PG'V�dA��t6 ��Ȅ��>��vn�3��mQ�WL�nC�p���/�
�V�+ ¼H��#��s��8'4�;�t�w1yG����`��^J	^NĚ����.bX��(�Z�6�A���X|��a��́��%EkS-��>��o��rO�+�j�=/6K��J�+���X�"ƈ�=*𾹌4\��g6n��a�kd.Y\�^ �&}��b�nQ��
��GC�?>��
��!4������D��(ھ�g;\WO�P�$xضJ�-��Kf�K�Z�h�PSj��:�y����=��j���Ȕ�A�cF{ �c3I*k�{2�_��=�T�B�b]���3/��_���(A��[c��R�M(�A$e�u�,�@)��$���%]�Mc^'��¥�خO'o��Ke�Y�Z�Uԭ�7*qY)��^��k���_��a'1�7N���%rPKg|����@B�&�U��F~b����<O0��*����ȝ�Ҭp���y*���I���w���R�� �Rø���F�
0�7��B�y?�N"�|�����d۾�
O-�|�� ��T�oo2����V(]��"_�II�� R��(�,A�i�X�3�|�|��"�1�%,��8j7��z��l\����6F2�[`ř1��ȳ$|*��2T�(��r�tK�_�̝�\]��G\��!J��!u5h�ɣ��OR���J5` )���~�OOj7�L����1wV��AJ�h'�O��l�/�����ۋ~%���1v��Ch���KH�h�vM��DC,FA��Oh��s;����VB�_����xv���R{��S��;��^���EQ��L ��G|R��]w&k�p����ۼ>b��(�#��d��9��l�W���q��L'��08�I��3��v���N��jK N�	���7:WA��%���UF�{�ߒ%<���'�&�X�5R������l��F�r����S��KYlWF4ݒjaB(�n _��af�*�bI��^���2���,�Ke�?X����w��L��u w>�RXAt�Q��P�/+a[+Gu�M��Ŷ�PR�P�%��d��kb8��� ��ٷ��s��`�$#jJ�_=۶���u�!cYx]y�� *M]�;�5���o��Y=������ v�31`����D
��P��=��_���W��!�rM�Q����Uo�Lr���;$=&f|��(�C� |\����C�Ŗ#����׹3�OM��������e
,%"fF��}#˕r���y�r��W_D�{K˶�i�ּIlҙ��ٜ֓�<;�JZ1�+O�e�����>�x-"=��bc�V.I!��X/|OE�f��Z�<�/aժ��@
_[Qm:ܕ����I\��0�Y����qYT�����j��GxC�6�s^��̀��M��fؕ�f.�@���R�dU|Ä�l�@�s.DGM�J0��	C�;+d�-����tbt`�2��3�(n	��_�5��/Ou����P�RT�̙��walbqH@h	�u]ҁ��t���� �m�����\8��Xӳ�lBF�R�*���/#nY"����oT����' Vfۏ"]�?%G_q�x��y �7�>0��fz�-�D0W�>y�
w�<E��F��uc���[՘�W���Z��:��,�IMO�Ђ�~ ��k��{�:q���N���O��=g�!k�[ol�}I0�P?T�$꽸�Yof�5Xi̐��>���J��^x��3=^@��.��ע�p���"���-Y8.�@��Y8Bk�I�����̫����'�64��"\%�ȋ�J3��2�=]"YA�Ԯ��U�`1������%�'ɕ�̞�#��R���#�0*����2�`8T��P���M�|�Y�W��b�_\�а0�>Es3ò�E�{�&:V,:Լ|.0�W�Ř��Bs��g�����;SM]�;{��rF�<E�f=ȋ����0��5\gE�Gk<�-��jj��x.q+z�y\�;szy�#o$d�J-c�	_r ��M{ӕ�����?�oo:~�ҁ�[kO*�����ԟS�`��>ǋ��ו��]r�:���&��F�J�`�\�so �����pK;UE�yG�_6�i���Za����!�� y���9z5X�h�D���u!����QO����E��7c缕�Ʒ�t%�ށ��S7���P��ݮ��[!ā��f-�/��h�c ��1���+ �������3��jC�������9F]�^�T���\�iT&Nˀ����w��	�����30
�!.f��+ml0����� d��W�]���â��:������4�ʞ���-RٞΟQ`����p�62.���F��ԛ76q�*u�)�$F�`ǿP�����qA�ݯr�WCKM�oyz�:Wx�8��T�D[����X�c&� d��=��U��J]Y���
;t�ɡl��\����jI�*��:b7�$ɊA��Y�M�Y�q���f&$�"�1#�*1$��+3��?Q̳
K~{�Q6��7)��Lmw�!-�v�<���ߠ�b��4��&�в�&�B�O7�iVZ4��mw��{�c?X�p���/�LТ-��Et�uI�OL��btI�̄Y}� �$�.: ���.�
�;kr��CEJ&q�n�Jp�؏0�=���o�T˖�I��;|.@:}^^�
oC�@��E��S����7V&�>fL�ʚ~� �.��"g<2gk�ͱ��+ˡ��K��{�}�n�UWw<���~����*�	+~M�&a�@�f�[��2`�>�t0�lm�9e�1��	v�i,ư�U�}��a"JF����
�<V�P��N*Ϻ����B9>0$��U6w��K�W�n�lt����;%l4%��w��ku>v�"�B�N���͎��ê�0�o�B]WZG�5%�1G�$o�W��26ԛ �s(P�N# �������v�1��T�#� ���g�X�B)Â5c�ZZ*"0�/Jh�VPy2�w��@�]V�B�`=��8ni�v��k���)��S�챤v�����N&��+�)�6,�e�"/��$������ �`c�6���}�ش�0�����i��pvpݤ~��t����Yp	\�����,�!@}hÙb١�l��r�U��A@�$�����<d=GߢZ�X�?���S?�|�<���Y����G���;,�lW������_޵����԰�>ueS� 6U����6�s#kI
�8��Gf3o�+�ټ�e��,�As ��.��:z�ł�����J~����MKO�y�7���0�$*�>��B` v������g�Fx "�B/���e��|�����κf�4�[],{_�sO�N�/ ���N_;k�N�'ڶ��
��D��Eq��
m0̓b�Te�Nθ-�U�	�)�ԑ	;�g�����CI$7׶��4Yw�B�֑�g4����+��k,t褹�L���R�4H>�*���5�~ 5�H��1ڲ%ă��bk�RM���vfji1e�V12B�����ӯ��,
�z�gW~�o�Pu��z���7�V�n�?-��T������M)V
.��]��WY��da_��@�v�)	I�3~$s"��M �u�`��O|xk�5Z��K���a>v!����i��ӧ�}!,�E	��ɼ%E��{D�(��@�Y���ѹ%F�U	1���@T*"�X�X�nSH�l��J"�H�7ڳZ��ucLкf	b?��L�"a/��+N�[іǍQ-��r��sb�b6ޱ�,ᦸ̃��?Z�Q�J��y�~��G��A��
3�Q5R�2�$�j�e��T+#�����o�R��Jfm�/j%|���Q�&]���D;!f��K�:Gk=���M��W9^�/��թ�4ym�Ь^F�'e��x9��U�D����5*�܀�(/9��gy�&Z���	�Jվ�ߨCq�o���*x8�1V����2�^���;ɴ�G�f���1z�ǋ��9O=�؜GOj��\��7��7�d���9,7\�̽���U2��$��VP�X҄!��i���nP����	�yK�E%���Aꢱa�KlƇ�~�a�,�dU�i8���_��m��?B�n�p����J�c�҇N�
ȳNb���\��#TI���i7�`���5�4l�K����0%J5p�[���?=�Rg��C�G�R�����s_t��^����N,WM�K�����T"�1�{�%��m�vU�d����0�3����6Kg�ݹ+��^����	�� Y��]�A������������8�A�^w�z����I4&�s��5�,�p;�
�'��k�W��~ZB섕���v�]�)[X���� �Nxf������J�Cp���ȝh�͵�{R�~f��N�d W�wOF��O�O�|b3�,�z���mr�z���X�,�߷���rzS4k��V*�x@u�~����k%�ᶏ粒��^7}1Fĸiw�@��鋡kG�MӀC�����wСm|D�Ɓ����8��Ȩ)ʉZ��Z��Z�?������z�?��:��Z��?�t�M�m*�"א���+�`b=�1�"��D�v��vW�U�2�3
��
��㳭9 Ҫ���	�D��k�9��@�7f�Z�5No��M� �R�oEh��ap��͠QzA�-Q?���j�$N%�N�JR���Gɴ����}�������@�R��PU��1��/�U�͝�R��}׫��Rr����4�l�B�3 ��;Sg�]:�|B!v}7�ƣ���`/ �z�#	�H�JB� �d4��-,�Dлh����+��0!'��5a�'��^�6���7�֏�x^�/\-7��V`�<b;��__#$�x㑺�>,����W�IK��'��dN\�+#_�%U]��������a�9���Ş��jh�vY����h^�x��f�3av��^z��d�?�L�4rv�2����wuBI�a��$x�� N��,�3��U&t%D.����w�[y�HL��WO�j�W9X��ܰ��S�bh�U��}�@d��+zׅ���`���isU��+���M��B�O�Htg���SZnP}<H���f���"�[k��Q!��2��u:kJ��0��G
�(_���5��'MV<,��ON1l<���66�.^::���&�O,C7x���ct��xǝF�,=�"<e�9�>�ʗ顥I�C���>b@� ��:���X�c���M�e�s�E�|Ǯƚz�5t`�z�W���S�A�[�f�T��;5���[9�h"խ5�si�e��r��Z����[�Ɣ�
��=?+��S��f�wpu���"�#�?��uƖ�
⧐�������b1Ju!iJ��0}91�*1Ѹ/�A��$03w�#䎀���H�ls�(a��q�v-t������F�h�5�>�6Ӂi&6���z�c,5�s[����"�,��e�Pc��˘a�ʒuI)a�n:A�;�b�k�X��=̀�_��=�� �r�Z����Q�M�������L�V�Eφ"���/]!A=;������y%��У��C$�?��n�x@����a�$B�yɟ��%t�������K�
��n�?�mەKG~�מ�`�g����<��ңf)@��9������m\=l��* �gT�7���/��E"��QG�)�0�|�KC�
;,��D9�������[��V��*EG�G�zLvl�uC~�lu���v�w�$B	O��
�-�r���ww�xٸ��Cy�A����%e&e��+��P��v6��f~�,�,n'i�2!&���{s�P0����^���)����*|�5{��bR/pO+�rA�hȊ��;o�{Yx��!h�@��Q��Ē(�ZJ�~;��=�]�S'�^Lk�Щq�d3D5h�) 4��� q�T+���5���;9[�Ui ����!ѝď�v�K�V�&٩E���	O!�0u��!��X@�T.?����ij��s�15y�~�(�ms�������\�X�:������M[�(F�hD��qϙ](�ާ�~�{"�:Z\��u̝�|�!y\��~<~������_�`0�?���i=�a�~����q�r�r�:AF��a 4`R��D�p�L��xX��!g.�p��
��ki���L�*�8�}9�;;��#��'���A��\�?�s�PJ7�H%;;����𼣓�$�$���u�w�5Q��~W\�Ϯ���!m�M�K�Ci�⍗ۓ@=�������q��f�����$%������?�~�{>�HS�5��N�@���g&�`{����m�Z���㜹�n�Ѫ��F;�Q;k������Yo\��o�:�&X�X��Q,���fr����K���O�̝��%6�҈d�܈[���L"s�ꠢ���Q2E�������O�F���0p�&�-s;"���b�Y6���u�T0�j��}��ܜ��q2~j	���aP�
�Ưfz�T�~��ڈ�:�S
��N�.;��f��^���M7@Rv��{_Bw��F%�D��mE;?! !H��-�0����.�*�`��Y�?�����#If����9��B����O�l�n�v�=V��AĔZ/��GO�#i��\��'��:��BK�c���yl��8��|P�����/!"Ax��5ܧ}�Pm�d��^���V<��_V��x��[^^��]N?Vw����X�'i<�����]��q��	x�G�֒&����J,22>@Rh-S��G0�:�����=@���o�1�/m�҂mI@�;�4�r��x1���P��ߢ��2;L�����f)�t�į���y`˸���T2�wwvg��I�Thqܕ��.6��XJ����؋�wcʡc~�:�<�oЅ���j^x�<B�-)o��J�,�>�p����w�X�.H1&�{A�6e���_��?�T�����7�%s��_yS���'	���u���i J"���$�o���e P��l�=��]�$�r?�V*�_e&��~�-̸�����C�$3��σ�X���>6�SW�PGf�Q�7��6x���<C����{�����͝/��^�]��eS��y�p�h]�?I�f[$�#Dz����&iM�D;!���+8m )K��I7��$���e��T�	�A�Ua���� �	{e�A_H0��.������]��5F�7Vppy�i�R��+>�.~�BK���2[�H2� &'��\�Z3��mV�����G�*KGK���zD�LHC��JS���>J�&��8G�ى4����)C`����JHC����g�Y�-�rV(�/�=x��4�2��E$d��ڞ.o
�4�([C�U8���_�������!!b�ف� Q�����	�wTwd��hqkw����%������=#;3��e`���'���xg��bG�a�}�l�q%|t�H�'��ݚ�vD!d��{a��[@����W���Sд����5�j-a���:=��m����82l�ˎ�zZ7�n�]|n*�f}ן�M�&�!�)1�W�D#�z�D�@�lgB�H�	��☧�x��2L���ʠ�u�����f����ܭp���L���Ғ�+�����\�@�V|�Zr���}��pģ��W������:Ơ«V��Ⲹ�/�ߞڹ\ń�I5y|�REi��;l��y�8M�y�/�����<Y¥d�jQ�	���p�!y�����:���1�'��=\�T��YDېٔЧ�=�q�� pD�.a��4�/V8���&0�1�z��)��҄+iy�ٻ<�(4�eE�n/D65qtwT4���x��U��
�=��fd�TFD�LX�?m��I�!$�?�~if��ez�{˼��,C>��C�Mlx^bs
ġ~n\�,���o��\��Z��L��r!�� [��Έ1���_���^�m�,��S0.����E�隹ǿre)�����F���h��\��:����$�Տ�����-m;�b�9��6�fw��{Z\���qn��1�\��͔t�>Hs��3�D>�z�]O2���CsT|�A��F����y�fM^���m{�f�J��GB�-��j���J"�%7������\w�x�55ޫc=
Q;�I|*Z���b�S��;������k�8�-�x��oIvA�U��t��4���P��(����T�"�堰N�ABh�j��u.w�����d ���k����Vh���{���4G�f�����~/��3�z�`pB���:O�Iki�=|%w�T�ײG�9O�����7<�7T�4$lS*Iq�+A��^o	p��!�~i �I8L��+�ǌN)��Q:�ع�1�5�`�7TԶ�vM�k��++� D2�*�Gp���
|~��
A? �I>�Rs;w�vgܪކ��e3.m�r�e�����Ip�}����/7�[4{{��t j�ڶ1涬_M�r*�ȉ&��v`M��p�Z��W.�y	.<z�UX�,�Ķ.@��׏nC��˃�W�Pq���X��ױ~+U���¢����p�R`�ˁZ��=up�k����?��hcO�EG�B���lF���Op��\
[��p��ʆA�4Q(��P>z��As�6�.8>���n�$uq�J�N�q)2L��*��D�hf��HN������'rM�j�����4�����ĴC���p�tZ�R�	��1�'�+}��0V���܂�f7��x/j�
~w40E�2ʬ�~�9�:�]����
���]Z'~D�X�}��i�Ù9�+�D��ۦ��T|�q���|�A�_r�[�u��)�Ń�؈�����̓�@�!�mG�*P��ar�Huh����ɿ�h�[��w��!bsqz����A�x�&���!���L�A���!~��#sFd�
����K���R�-�U�3F�����w���l\�/��Ey�pa�1��^��b�ѷ�m#��]k%F��:'��FG�u���Bੲ�+E�l�jG��$h�j��d�@���8d="㼮*	���E@�םu4��v�`v�ل!'��PH5b�����߄�]A-i����N��2�K{դ���4���}@�Ft�z	m��*1ٍ(ps#�ћN�,�cj��yo:[����"=7��������TR@�TVП=>����a��KW�ZI��F�/�u�ES<������<+;�o@��Nt��"��������N1�	���o�Mq���Z��ۮo��2u�d��h'2�_�+F���D���_+k��;n{a���bG_����K��b���/����?g���c��p��zaS������:ꙫ[���Kx���'���L�tve�}��N��Y��#ȭ+�;��b�z�c�J#�ΐ��R*�uoE;��dW���}4�Jрb
��R�cϒ��x\ CR��n|��ĥUݑ�3`'Zd-�>�g���-���$[1���ι��3뙸5�K��dm1VE�*S���6��KfU���.�A���S�ɕ����ÿ��lҬ|�?I����O'�P@I�����@���׼����i��j9�� RIj8Z�yD��dm����F.::Y��n�#D=h�����p9������3C��һ}Nt�Qj|��~)��R�'��_�H�P;����c1�Ъ�	�%K]�5���l��ӈp��5���5����nَH�_��дm���"g�%����;��n�M�?�8g�XZ�`�0��E��R:�,Y:+q�^w��I����z5��x!w�%5Lr���7�x|��Rv�r/���ӯ2&�[P B����$�ǌ��1�k���x���(fE���oY��c�Zl�&�ڮS٘;�K�����KB��ﬅ���%�;��I���C\��֊6�`�֑&.k�~��*�C���Z!��^!����y��5�~�&���>�l�%��h�)�nM��tf��Y����L�N��H0Gz�e��SS=�ܒ������=�zt����;Y�"#����=n?���u��^����D5;Nv��J����<�}����Y�;�8�*�yHŔ+��}����S Gϑ��o��]���kl6�g�bPtf�t\>�nR�Çi`-�؄q�E�_�������tL�&+kmʳ�r9�%������pF_h��ՉV��J�>(��*e�t���|ч�9���d}���ɇ�~�o�~џ�X�W��/�龠J��{�]�K�ޱ����G,'G��V��|l"sU8v�H^�D��Ew��w�p�\�
���v���jAV���Z���gd����ϲs����#�8T�Ǐ���}G-���C�"99��~�(��f��hxy�8�~d	4�x@��`q$Kujփ�=�z���O�z�֔pOЈU2���p�A��#�qr��q	�/{�݇��hSO����:ed��5���{��t�U���H5��c��a�1D.g�%R��_Y"Zt�%k���O�X�ފ)���F���GE%������"�����p����+���ECZ��B?��?v>��}�\E0�[�Z�=�[R3��ki��s�vF.�����C+�����lY�s94D��=��i�um��`��VXa�̋Z�� ����I�]Aa�$���9�U����J�M
}��WH���|���ث.=Y�\���g��aa��,�y8��<�9��D>}2Z_�"�0b$�Kl�d<�մB�Q���Y�z��$�E�:kqd9�	�����2g%T+W�>�Ѷ0E̐�5���N�M�@�ˉ"���/�s�}_�a��ld\R�>��m3�L@x�w-�|F��'�3��:na��Jr�9i�O����!�m�h�t��t�|Q��	"����!���sͽ�k<�WN;�&�T�喬'�ޜ�ۼ��v݈I��hď1O`�Z$Ϋ�}'��T^͎B�� <�ܮ����k���t%#Ӕ�C]{K�V��r���Hu�y}D�@d�?a��y��D�ىP�<F��Y)���ɝ]��ȱ������g�'�M�o9X6�,#7Qy��#-Ego�����Z4�[6�'�F��P����C�W��\޸8�Aq�s���L��qOm�}x��)��SPO�	�_)�khL� H~���$C�������>"r�4��
��y ���>f�~	Wa"�h�4,ѬK	�w+'ɍL	�N��~n�d!���2^v�T7p��8�;^rvtY(�Ў���h����������������� �ְ�A�IGk����븣�;.J	�vv���讻�~�*�`F�Re�a���(߅8H~C�`���(cU����2:�$G��7�'N����.pW��T-�I̙b��u緀BzM:W��31�����qw��������b��LJ�^�RfxI�b�G������bÔt�]�;�bUu[�t�L /�UQ��l�2�2��?��()�q�6N��� �H#�մBα������5�]ݹW�Z���2�~�z�/ڦ۬cEV�bi���'.5�C�!���r���R�5/3?UF�z.(�X�P\RH����9���.���(d��V�a"�	�(k�PE�`r`B�� d2Lҡ�uJ!���J�,~��+�)H�3[��< Oo*.n6�w�OCyT�@um�i�{w���1?NW&��	]%Gt�F�Fผľ�s�u��x6�+ʗ�X�!Gb��ќ��]��+K8�"�,k�vw4+��b��wAY.���z�-3Ʉ]��˵Em��ɸF�����;���,B�(,�� �k$Jj���!˚�f�/68�\������h%�G�LT�(���jc�K�f=ɼ�Â��k���JT\��*!����x�y�5��b���6���=����f�a�(qkމ�D�"�{�F��<���L���;ݲ�G$̘��Ⱥ��y�k��`n��٭���Tr�_�۶�;����uu�������@�z>�m�{���'H#��[��k�֓�X\�J]��ǫ����} ��MF8c2"8z����=szv3R�.�L �dC��iՊ�P�2n�'2���L�r��4���F��Fz�����:9j�Um�u��P�� ȼ	��K]9`ÌB��f~\�nrC��$��7'ӳ���u����{F���T���:����nD���e�ٲ�E�����Ư��t]�'6bma*��<ύ|�Q}W��D�$�:�n�L��c�)����[�x ���,��}-x�ۧs3��u{�X\����F�6W|{-J��S����V��"S�Nϒ�+��� `&9�+|u��`��i-F)�*.ӃP"�� ��8l3@ͮhq�'�;Th�X�[��M׏<&!À�y�\�R�!:�MQ��4G�i���{fp�;���-�D�l_�{7��	5� ��-h���[���I����۝�~�gZ���"�������.�)�?��a=�k��u ��5����U��ȋ��G����<ceë��hv���	�z��_*}ũmL�z>�z�r��w{k����.a��=h���>���+�4�e��UçIb�S6������i5N�K�^���n�x3��l���^��^iW;T��*e����O����88x�5�aXd&�qg�ef�X�Aq �����#��~;�d~n�H�r�� f��V�X$�&��+���)^��?'Ri\��jw0�&L��h�>�7��Gb�a���|�\����v6�;2��X9���1��D�b�.��=��?��F�����Th�y�5g��0a�&��v�3=sz��> �kH6�	�a��� )�>�\)�^�q:��b۫H^y��
��P���^ �ɡ鷛Y�>	\�����@�C������{����T���K�:��p���L� ��V��z�V�i
�I^�i$�l,/�v�Q���;��l=)����h�����_�~�eCT�ӽ�m"�f�R�O���>8� 9F�^��<��Ζ�b�EW�.��0$�ʣ
�FZ��8�<�Z4n��-2��XQ�(�=|�����2��ƺ@�&�'�����9A5��s��Lu���fe0��|<����L��sx��\� {����؟=|��Df˶S��_�Y��R\��,W����L� �~��I���A�3ҐηM�w�#&꘯�]�΂�MV��(>x��f��݀M����Ծq��=j�H��[�C�0Fpj��ܣ˞x�O�y@�s�!��)�ǼX��6����ȟm�Y����E/��U_8;�I�}��sM���]��#��_�^9x�Xb璉�5����j��Wv�j�����t1'ʱ�oR\�#�y�Iˀ�m��j˰bm1㖻����6<�3��G|����F|C�/t��v����_��V�����O�ʃv������$�r� � ���hvvg��]J��#�����l����c���f�g%r����>Ȼ�ì�[~�
�;o\�E+?4!�������25��޳V�*��j�f��K�E9&+Ӈu���h�в,��z�����h�)���NB�@��e؟�#�gK�� C����H,ho}	��Qr2K����<�n4E`��O�Y �|�����	o�І�K�Z�nXU�'Z�_���u�����	<�uG�r\�'�{N�
���� �cS�iP6\[1~�F�����S�)Y3N�]l��QѩX�'�H�!b�ϟ��ΫŢ
��ƕ%yz f��s��� y8�5q16�
�U���¢��$��4���x�i����l�K���`����D5�Qh�taȘ6E��M,��X\q��y(�n���S1�?�b�A�6jrPZ�l+F�C�Q@��E�w��v�ҳ�5����Vn��l]c�=�� �'�q�c(R�i2J���x�m�|�ʞ�a����dLI�h;a�"��آH�Ty��:�,*2R��m�#w�}Jf�zC�����]t^C.��n���>��Tzˮ��NFD��w��;���7���a{˘��n��fc������5��S堆�Z�갺�?ю~���;�;G�1[/��TR��z�ĖXT�zJ��L����m��8V�8sT���1S�u����೔��uy��1�]1r@MXy�5eҤx.��/+���.J�s�I���݅z_��݋�������7�ED��N\ET�T���aU�Ҙ����&���g��'�n�k����O�� ��ۢ�����O�k��>�����Z�U+��4���$x	7
��;�0��C���Bk)��S��Mě�ni������@�('��'�e�&���~����y��M+`H��ɰ�Rx�	Y��o'�q�mX8s�����igy�$���}3�V�c#���& ��.�"�枕��ON�c��q:Jo�uAFI�,םmK��=f;���C�匶@I�d"��v	5� �?�����h�!j�a�R������;���O�@��0��s胴*�O��p�3+�cK��G��.r�AvAcag;��x�zn�� !X�q��2�V}S�qH�S�:4����I����uԉP�p���@�^i��Y�`E2��|����?�F{��u�71��<(�� �g.s62�y}qh�B�^��*�hާc�9�76%�~Pn��7r0CIP3�ZQש� U���D��OfÛ�mW�N���$��+�WN:�*���7����P���L�Ϯ|#��8Ѣ�f=^m�I�&���Y)بw��a
Q���nd��k}dT���c�a�<P��0��������f��W*�N��3P(�V��i|f�y"�#�b|�^�*u���N��q��B|����ik܀E���CMQH���5n���<E^� u\A��菼X�f�D��} ��z�C����e�\�����Pڦo�\�Tyr�f��t1�hQV$ٛ`r�X�9�ȥe��^2[mRO�^�h��d:���D�,{�c�`~s���Y:�^�_�+�!I�QLz?!>�x7��K�W��I�0�e���p ��4%�)DBI)CpM5��ԕ��/�cHi˼|!!�����Fi�����j��gs��z��3�Y��K�F6��>��x�pe*�qVk\c�e�R�f��|�������d�Wj�H���L7a�(�o��F�Ѐ�r�l� �e��}�rS��{�P��c8Ո.sgF d�8����?���5Za�]\��Z��bU�(��꨿�k��2��gx$e3'�P�/7�Դ�Ǆլ��gS	%,^���+LpqIӅjF����z���b#���XY>��&�v�5?tr;��ߔP7k�b�������R>���\V���&�S��yn)�Nn�2+e��/�
\�_'!S�6�s�I�=��(XA�?ڈ���6�ͦ�kSNr�#���ջ�Զ�z�:� Yb=��Ц=�?�:Q��r���V9�Pb��wJ�� 1u��{�#u��繀�!q����h��a�Ć��d����/ �4G��그:��2�~&.d�Zh{���&^��f�g���R��������TWy~^>�A�~���_���bٛ�}�,��wm8�U5��mۼ��C����GPrq=V�뜼ƞ傻�PY�}9�����XQ��2�-؋���	
Y�PCx�b_�hģ�#4����ux�̜K;�/�Q%�jc20R2\3Θ��f� ���,D�Z.8�M�����4�mř�vC�	�&��b?yy{�N�����:��)�sT�n�DD�'��ߍ"��7O�g�	�'��t�;ށ�a� 7�Rb_H�[K�Vy*�T3��(�s;7Y�9G�B�-�8��ٿ��c�le�-P�5%i��3o[��A$������j�z�C��*��p�j�`NUυG�Dv?��C�Q��CV$�,p~�8x~�>��@�gH����4��X�A����G�ߪ՚�����d'�4�Y�Q�����|n0�ddo�@��aO�hE�OM ���?b�?����r��)�!��<�)Q#`� sJmk6��Ţ^~63V~�
@����i��Z"L��!W
�GX�۽���7�ҏD��*�l���J&�U��PU)0�Kה��X�!�3�ؼ���hȫ���s�B���iN<`�zE��?����_Ň��9y��P�[�9�MN.�V��,=��vIZ��ky�ٔ8�U�ij�^cJ�.��R���d$W#���bo�p���	2��ƈP�;s	e7��o�!�|='pe�v���J)B���,��E�oa�\˩x4։t��D�)J|M��<�9f���l}y�lzʼ�)�]�]��؁P�yiߍzs�і�#{�Wx_��#RF_��{�}��Ӷ����@���	��'\%x>�*[9�<2��5730���$~�/hp��@��o���P��^�����o��J��)�$zkbA��E�k[���`L��d�m�$QCB�b�W�:�Nc�o�@���Ri�w�m��Mة���!~@���i�l0��P�̈́����S����i��I�D����+�o@�ѡ�Pn2n�S�]Q�����G͏���` VZ	+26�e Q����?�67���C��3� o�c�����xѝ�kkhy`-��ۓt�{�_Sk�~Q�:��*	��<ʡ�o���F?��8̃)��>sN�K`�,������0Ѡ��d��e&�ï��\5+v�����Lj+�u|ʱ�(!>2�k�b�E	ε�6��7�m�)�o�w����a ���ifb��	��G#|�=g*�&7��tıh�Ho�/�K}Ñ��n�~�*��ϫԻ�L����mth_BF[{=D%h���������-)p�`�u�B�q��s����oX[�7��;!K4K�؈޵T�K�$0�˃'`o%�����B��S1n/(�9Z(���.�7YXb	z�FsC��&�o�f�����d��M��M{�qa9�R,�/e���p��^_3Nܒ}Ғ���_&N����1B�z�b��24�#,|:��&��#�v�~{07��Y����2:?P�/�PR��C�/�p�~��m�F1/�-�h��0SA��۵ݹ� _��ɻ����^�p�~d��a����v�pֆzmuģ4��Q$��%o�T]�O[c^�-jF4�@��V�%�,��D��%".�1$Y�eӷD1G��8�@�2�܏�/��Zp
��4)]�w�V(�`*,�b‛߽�G`�d�l+ hK/��^˧�;Gv嶩>2*��g�����6B~(6d�H��)���
crD� ْ�<���{�׏��d�0~=�|;�4N��a�Kc�Y�oçݐ4�V����=�� ՠMMTJ�(�i�:�ɲ�4YΕ_�.s��j����gŐ����{uLqG��/�6E�^KA��P]��Bj>"m�G��e�9��|�£�M�E[���K^'� �s��|�`��n�0������[�S������rR�d�^���0c#LP�e%��^�J��M�����E2�ެ�H����Z�u�x�(��Dc�g�̇��Hپ�?��Pzxߠ�������{[?��}�� �+k��像@Y.����h%��[�0�ơ+�[C���@�S�8�=-Ȱ�K5A��
g\�Ӌ�l�=/��􆯖���Hr�%�8���q�
K��D���;�Ե�n�Bj�62*3\�^���Ր��Fy���M[�+!6tHl�h@��aI�'���Y�:����3��EĀ(�*���_��y>x9Ӥ�7���pȼ�d�YD~�h���
�e��V}}�J�A`�n���\��K
�{8�I��~�O�7"��~����Q���L�I&����l[�l���Bl��^b�k�pe��M2�d���?�kR�PFy�u�np���q�4SC�Wj|����z���,F_�����p?p��c]�=h��`a���{�"jYϐ<O<KP& /��I*��;���wb�,a�f2��#�7���B�(!\��I"s]�wb�3��$���)9���$�ϊ��`��qG�ϬY�s��0�zd<�Z#4T]���oS<��lk]� ߇l\�Z��>��@;�mm� H�PF��=|���O���G5��H�}p2�6M��Y��}£`7SVT%X��!�+&D�a(�i�H�x�O�8µJ����K�/j.��D9�2V��5���ߚ���@��Gj���W���7H5����~	��sU��\>s�(����b7	x�ڲ�!k�C�կ\G�����a����C5>z�.B�V�w�õ�64���C���a����	�N�ΫR�.�̲�b�Tc>��F$aL�m��	��-U�]��x��V�ؑ��mmLy�ڴ5V��:��7l_�"�3�f�+�d� ��m�h�5W����'"E���Z��{����o����TڻƔ"�����8�ˋ����F��U��έ.�B�:`s���Oo�IJ�B��U�Ù��dj�{e�O�[h��iף��𓲉�65zX)P�5�Ohh�Y�M��4�Qj"���6�?��� �v�����+�\$��"�3Il@��R&uM�lHt�.���ԕ��3Ni\�7���]��K?3���ޙ�kXƾ]"��I�m!�]�*s�Xg���>����8O��-����ϡe�?Di�rH��ˇ�='�#�y�dmŅ^on��H�����sE�n�x�YE��)��-K�*/���.ȩ�B�I�S'�i��d�ْVΥ��\�S����f{ފ�k2e�ñS8��v��WZ�]���+^���p�OױG�x�՗��c$*I���y)���me�.�K���lt�	ڈ�_J5�؟L�;��TP�ܮ_ k��?��sd;���ꥍ��xS�����b��ƹh���&��>���g�k���R�� ^Ҁ��T%�BP�����A[c�5�#��m6_��|���ȭ��7�*�������Y��.濫e���02����^�hǕ�;ы{V!H�L�wӲB�	����@�"��p'�I���:��޳�x���߭R�3��m}[J����s�k.����ĉ�:c����-`�wC�6��*����p���T��A��/x��[���1�ϰ�ѦY"p=�����,���rH���g�w�%�2�Zs
�bb�;T��8�{*�bz�e｝tm=��M���#ezp��G�́m����ڶv�2��˼|�=fh��~u�u�	���0�<�GH�,�R�D�^�j���Zk"w$ ���A�UՅ�l�S۱S��\��- ���z��P��]z�eq_ڥP�)�>��uw�f�8�g���ԊL�w����
�q.���`	׎�N'\#��7r�.�{6���*f���d�~6�ce��������;�f/%����tm.~v�����@�W6 ?��#3�u�"���������~mВ�EP��j�y� /����2�a���A�[��R{ {l�1���n�շї t���j�q�]���p??s�t�}��Y�����5�V�
q��f>�����F������ߣ�q��-މO��#��x�N����`��R�-!�`�ܙfE" ��S ����ޤ"2�/�#�
2)FS.F<m�~�<�"Z}�Jx�-�ѵ�A��䦻���Z��GI6� ��7�U]�b@j����11��q�|h����Y�� QJT�%	e�,)��s����^i�>��2�!�mݦT�7�L���",�4Q�Z}c	�^z��Xj�U�<��o�����}�!�S������I���;�):���Vc;�6��s^������4���z���ũ�xZ�j�Rx׷��K���N��yt`�&�B�n��
$����ӫKUY�W$��×/ą��j��7Ηθ�����Q��{�p�5�� �t���q�3�k>H����^� ���#"�d��v���6V�k&���[�<#��`�z�t��k�;x�s����	S��	Ή3�
�9� ;B��!(�26!-��e#3�T.�R陁|�JK@��6��VBX׫��KK8VWU	J}��Np�>q'A>6��Ě*0���1��D֞=��t �,�ɿ��T�1�Щ�z�o�&W�+�CԠ��<[�Rg߃]�!QC.\Ã�r�7��&0:���O]��(��q6-6���+O��3A)���}�%�}-�3m{/��W�$�u�Jyf�-�"��k��%�C�?�;�D��U
����d�ɳ��F=z����0�j�-&_�^�)���၏e��[��e�������)nK� �8H��f�G��v�
JǶ���pS)�4���2'rL��ep�ǧ�Glqm&7��v�C�}�u�kE�X���j��;�dY�z������^����qō�1�\4���VȤ�0t�L�D��&>�1�)���p�`�b{�m�vL��N��p2o�S#|�%i�U�l�h(�0�q����]n��X��֊�3�a\5��<85V�o_F��,٣T{�'`��t�Sr��dR�%?�#E�cm��m�~�[���2.��������sh|�|��̘���)g��\"�`f�GR��C���Q�6�~Vg-H:ޭ��Tj��,�)P���s���	��!&��ϒ�%O��!��c_J(�&3��3ߣ �6��]��f;t�bI'��Z�쪗 ���*��E��eЙC(�o�u�$���ȻJ
Om�M$g-��n�(@3Eޑ��V]�&��:�Yg�2�nC9�l��S{n�l�D/�����:�)�����.?q�+J��n�|=<��QCe���"y�:��-�¨�a*m��,�fc�Ǻ7;��b���A���C*����P��沆�E"L'��Ox�mS�Zps9�2ኃ��H�1�ی�ޖwO�@s{M�F�h8��<���TS��ހt0�vYC�ňr(����:�P(��m�I�U�_.{���V벖�|V�v�8��a�qid��Ç�l���;zy�ҙ�V��I��*���QYy=66��� buWP˸5g�v�h`����A��o��f�]h�#�,�m�� S}���{3�?Dd��Y�I.Tx|�R�n���ޒJ���1�_fts���x�|���j!H�Ņ���Y��K�c�>�D�<0���3q=y�MN]�΁���ItK(�9�/������=m$����*:��X�6� �^���,m�1=:G3�МOO�\�G!x���sؗ]�������&��)�(��Ô
7gb]#\A"�ﭹ�(w�!�&�n��}��p-G�
�}�:��%RGUs��orc��!C��cŽA�i���"7�َ�\�}�aΉ��}8����`/4����Q��{�[����w�a��Ȓ��D�>�
��T�L\���g�,�����9�#u�`��؇aH�)J�s8!��`]P9G*�	�I�[0Yo�I%�2Gcs���V�h����n�r�4���j�Z&@�~"#AW%�	'qĶ�c���`Ov"mg*#ܾ�����,̨ܫ��5+�vy�̶@��$U���V%���P�ˈ����qOR=�"�Ğ�(�m��NЎ��w�n	�1�.�������.��B��mɦ�{��3�Q�^᪚�
����R�i�g�-d�U@k�lt�mJ�7��)G�u�������X�^8{rG�ab�F[%MB�u�c{�r'��It{�J�,U0\X8M�:Q��`֊2����H:$�����j2�l������R�Wێ����#&�5�:p�o������ۛ�B]���]��Fv�;̗��'Yx�^�z�(�G<"�T��0S��B��+��)�%�h!6����&^k�\�Hz�����\�~�?q�6�-Rx�Q���N��ª�$ho�u������Љ�̐�;M�|�=�;^8y�OJ4I̟�<�)hw�[m���A��* Ve��Y��Q�t����F0:�����?�M���+��V9���dWJ�TN�_{���c=��g�̟�����3NǨH��������\e��5TH�dNamC,����r����w�#W^�\LN
�#�U�μ���Rz>m
��q�j���e��~w�S��._��N�B~�g�XO�ճ��W�6���9�ɸ����y��2��ѡ�l��SNpM��Z"�;L�x�� mݔzzQ�綠u��]��K�b��!�u���H�]k$WI^Gn!.`b�2��]���|$�˝R��H��O-����iLv�"ͯ{-�9�>$,>��1����I���,t7x!2{�6�غA�XGf��/�\�?P�oٜ �0L���م��W�\h[Tk����G ���hZ�D#�sxxŽSHjt�+pW^./�vM����F����9��%4��g�'�`.�ǁ��x��\k�]`����c�0�?̈���b�k=k���j#U�+Ͳ;W��n�	Ve*�`�Kt�^,�pZޅ�E�����e�ޢ�_Wg�8��Ky�� @^�ak����8�=��?���h�=RV+�1�ʐh��z�Ny�H�]�:4�0"�����7����3��I�4w�x:�f05F-�p͔�{ik�q��d[=�V����p��oi	�?m<ȧ�&��̍|���:fu�m�"(l�K
����GS�? �qafӴ&�V���� �ySJG��x�(�P����.�]��DKQuFwVZ9b �%ym��[����9����ш]R��p���$`�OY�^L����៫9��=��K?�XNb�J{�~�4|@��D�jOk� @Tp�T��hb4�ս��N��&L=]��<�)u������E������(ԙ3Z��lTִ����F��siH��Z�>�r6ɂ�%����wP�k��b������=z������
#�����=-�
	���A�7�vS��|g������%��z���i�?�ȕ�n�C����1zC5��4U��L�������]H����Q��K6���ֳdB!5��~�?]�f�=�ub�}x<���~,I's{d�&y��;œ�eb�4����А ��ZO��&u�[ �&y��F�R=]Ƅ�H����DsF�6��|H�]����PIV����븍�YC�@�T��2d��$ܚ&:���C���U:3�:p3e���v �H1d�T��љ
I��tב�o�%�4���z����u��	M+�X2����=��2���dX.�r����m�9e���u7�w]㌟ �%�!�]��r���4QN&�Քm�5?F��ބU�,RX����ZbH(��1U_O�|�e��_�r" HoZ�Z�HF���{,H�\$R*W*��0�ζ��Һy\�pMQ�J�����՚G(-V��E�&�ik�59�)K�H ��n:]nT�͜�9���۲斐4�_ֳ���r��9[k9��1�<>2e԰��)p�;t�ak�u5p�n�me������%۸�O��GC�����To�
M=A.��M�Ǻ�طj	L���ҨFl�;U:����p��x.��͊�)Xl���%�������
��.�sPx1҄�7�,��~��ơE���`�i�jgW�&�v��n| �}�l�t?�e�>�K���zЛ��!ׄ�M�SR�g�����H�q<�����s>��_�4@͔hX��m��A�`QNx&�O"3col$7�E��'v�
���Z`b`���<���JU(!� Z���
�i��Ǭ����>9��-G�%3^x}��DQar�I�~AU�`[�Ɋ��IX��i���>g�Ż�X'�jǊ�'�B���WJ���=࿑M�7���ɻ�^�ޠ����J*�{��4��rA]f}��(V6���*	�5�"ٙ��_$��7Z��|p�"�U|4,���3Y\�U,cY����_m�"��eqB"���º��	��v_��Z(��^]�;�����B]�mM�iL��*I1���j�-x���>~ ��@�y~�fи!��Ӄ@�5ݨ�>k�A�[��	͉ �����.	J�sqh!bÊ�gĖ����W�z�5X���垇�&"GT�Y�e���&)t��q&"^�1��>������q&�!�焕C�o�N�6�!�X2�K�Z�_�/ki�����<�`2�M�����@�a���jǆ6�o%#]t�uܞSr E?�o����2e��q�M�p5�$��Ʈ�/�:'/��Ӫ;ݚЅ�s�#ĖO)��ON����ثc��-�-=R�Pl�JC�Ԏ�aܐ��I��oM�S�?d8hs�9H���jP@��`�B}ַ3��Za$��0R��.�Yf��]��������ל�qFJˈZ����k2vz�z�BѶl� SЉr��Q�O�i�MX^$t��>���ixq�����V����o[R��Ց�ι5�ݳ�����0v�7,�;Y�p�-�`q�������S>�]T�[�n�= ����}&�C�r�lv�\� y���\�:���E��ƅ����?�qF�Ňz��w�vݎ�����*�v��θCA7Ƅ�)�[��ø����yf/k�Hl�o%+��p7�g�����	�.wK�⽦�o ��c� 
�f�!�|,}�[��$GQE%y�c�������i2�6��l�%���;�������3ɴ~��=4C�Z�(,N�9l��1;o�=�Q��Tj9�!��UeC�#���i<�T�jWO*߯�&OM��S|��L���L9�2E�O�c�X��G���b]�:UPX������ώa���t�w,ӌCj�qgS_��{�u�Κ�pC	�k��&�:]�����0��_�(7�CZ�8����_�B�;y��".����9�������-nL���Sp?0�3>�y͔4d��p�<���B,�Rʿ��#Ƕov-�!h'u�r(_�KMS�� u��§����w���!����5I ��Kv��:͐�� b��-|{  �oF�k��]@no�3�vo�D�a/�2���:X�}�v��L[<i�/��(�=tC{:���ɝɚ_�l��"ˆs�]�}�ep�C�vh�Y���d^S�����R�9�'?z�P�IK�d.r�Iу���B����=�|�l�~2q9�B'y)_��¿�T~�?��G�1z��&u^Ɂ;8�Cq8��T����A���)�� }�p3t�����w%�-M�ݑ��/�m%Tp���pa�!�ւS�q,�*�D�����4���j�����ʀ�"?4����7Dk�_�g#�7�<8���Ò[�'�H}D{^0��_c�N�s�[�����R�"�S�Gi��������T^��o�c)P �mZ��u�H�f�u*Z$�QD�Wa�Wk2��� �*�D�yT>fʚk7�6�H*��@B{\��_ �,�m�n�랔 L���,�4D�YG�Z�������J� �V��p��g������Y�j���/Js�1r�m��DEӌ�ԥ����\�r�Ά�0ꜥ}�+�����4d����27�'a��MmUϝ��\v�����R%d̺Bkjb�׭�~�7]�U��B�ܧ�Y#Z0M�}:eJ������~?��X��7C��u�/�e;�~Ioȵ/�Z��\�b��9{�*V�0��\zQ�Y&������u�z�	�/@)��X�MD�2*|�\���-�:�r�&�]�"�0%>����r����[����%=�@M�����I�_�]ʵȐ��ڷZ���΃�b8�B�M��iNr^Aք�Ie�o�ZS��R:Ћ��v��ȵ��͂��#+kU-�d_��SGa�CU���P�8�'e1�j>�`�Fy�y��=?��^����"̺ThbMbɑ��C��U�%<��m��A��˯]G�y�I�g.xK��d��o��CK�����		��9TE-s�
�[�g혈��$��fO�BkG�fx@
�~yg���b�� ̚s؛�i���=Q��N/7�Gpb�C�t�D�6Q��9Ά��dtRXV�Đ���q�9h ��G�<���'��Q����^mM�?Ѯ.�k�F1��o.~=����]�$Ls����}xs��g�����Ka��<�E�9�ݍ�����?�ɽ;P�LZԀ���$ٞ��[੗,��w�e+�㑊�r��d��}t���}~cZ���>�#��t�رG�����_�O���I�|��]ⲧ�ӌ�i/�<��r�v�����c�.�4�������7�s7~��P������X��=�������|'��I߁F_�hC�=?��L2=�2�
1�p� ��&�JO  �J��5��}5[�U� ��M�ˈלJ`\f_;#��rL��3��lX��MƊTm%l��+I�R�e1�����1�7��� ����t����nD�KR�:b�7V5��$�Ψe#8����gh����ԇ�ш�J{�� ���w�FQ��c��g�������̷�/*[�`e��ɲC�F��j%�?���	�N����b
l+�c����=����?��k�ʲ-p�T^w�u�?�7��^�A�Xv��r��.��*/߯�a̿��Iٴ�+D��D<d8Y��j�W��F��%��PFl�W��h�M��/���:�a���/������*���C@��k�W``�X�;k1�䣄�sGY1$��d�����܏�J��W��JӝAo�΁�"���'��ʤ	��?���-]]�v>˚��w����C�c�h�tG�=	t�!���\�j�)�=��W�IbS�ݘ*hU��(��$��������ʭo�[n���n�\�t^�K�tO�Z��'�]��$��7�I`ܐ��F(+�M���9;�n�3�n����r�N���Lp��m���,S�[�psC�:����>5�`��]�ȵ������4��I'g}7R���>�`���%�.�]t���7E��B�-\�'�AAPl`<\�=�-�ƓQ�^���Ӓ&Msx=D��֘|��k�>}ɒ�M>p���E*��Qj�~�UXI
�kh���_^CK�!4)��㴴���}�ȮF�[#R�㗦w'{ol"]�g1y��R��{�#�_�.Tx�������{����.�R�م��}��������%t�mԥGK���]�$Z8���F����̎v&������a̫Jb.�n��!x�yi5��찚��7����w�F��g�L����Ɏ�A���[�zl>�7�k25�ȯ_mIN5z�.p�������Z���6$�X-��������B�2���wM��x�|va֫l(B�V s`9��d_B��W;/�{|�jaD��SW@_��e�Sp��q�Ҧ���W��VA��GQn��r��G���M��/�[{������鵷�4���tm@P`ַ�*ޖ��P2p��䑗�͑n��+PlXq��h�4���[{Ƭ��ߤ|��&A�;K�r�@ť��}�������f��l����f�/�L����>Ry�1���闸�ݴLq���uuv�cP�s��$��c+?>-&�Yǋ����,��|� =�N	jٕ���F`��e�o�}�?ӱ}�K����<<�q3�Z���?������#��\���$�~��w���.���Y��Fw!�h�eNXw��t���ߩ�ⶾ�S�>�S���r�-}w�PX��(l�A�6*��	���{�,��N�`BM�Ǳ�S�}��.q�L�! 5M��Jk|�H�9
��Ϋm������%u�-�Tρ�o9�.l��p��Abh�Ѧ�� ���
��'Y�0�=U���m"*�5Ǖ^��]�\=�f]�c:�B﫟�0'�|�4D"ɒ̂�d<�E�%���(O�,v�/.�4bfz��$�n̚���U�X]*V��NJ]�u#�ܘ�5����IQ�������Pd�$��<�b+*���x����Vz櫪����6{��<���*��[ ێ:C���H��(���P󣥿����Q�k�Օps���h�[,����C�#BN4��mݷ��m�.�P�ݢ�S���F��GX�~$����T1E�������&{�����u�ZHP��G��)�{��!Xc�Y�5��өT�s଎��R��G�H�O��]�ͦ�U�-���5Vi�����ƴ(O��cǃb�>��DNu9�ꉺ��(5y���� ���5��L$��3D�1���+V5ҬU14פ7���d۰�6J�Űʪ��I��Q��DFw]%���ڠ�hR@�=�N����K���)��+���x�vs���r��Û�N+�5su���_Etk��'�hn�6nؠ�g!��d�<��������$��^ő��,��dH�ݧ�[k��jMN%X�]�x�N�/j��W�B[�-ǆ��lo�Ss�[��H� �6a[�G�b��HCcm$ʯ�2�Q猷���_�j�����䴻��!��j���@���$-��{;������]Q�g�d����Н��}��zQZ��ta{�<Tfcë��G�j�Ke;���~��U#��>���)U�b��/gXė�o�V��!pM�CN�H]$P��s3m��x�,4����^~�Qݥ}�x&1\ =d3D+>F`��X�[��?J�5IW2Z���F-��Ůkh�)�1
�3�N��LP8��8Pi"�h�$��
�ԼG��6��aI�_a�g��������Ǖ��d�e?\���_���v�Iz-�X�`��г���c���9�n��o���}��|��s�� .�K@�!9�y6:{dܿ�eQZI��ٲV�`�����?;��&����Hj��؅յ�(h*a��]޷Q�=��vɨDe��l8�;ȶ�4�I;�������졭�vr�E�a3�OѮa�%.�,ڍύ���hH"�j��"\���.m�k�MYf�}W$�����'���pCQ��[������t@�>����3�b#̻+\ڎ|�Z��L١����h���*�@4�zz��J��Q��k����t[t?�!<�W��`E�R��5f~�(ۣ�7b�c�)�c�l�id[[��m}6���󾯌P�>�李��m&��^v��L��o��Og�	��E&k���4�������1����[pNKu����(i�H��'Rh<�{�Q�!9R扦'�S{G2<��KF�>���L&���2�5��� ��Z�F,������g` 5��U�1ה@oJc��' ;���/��L�Vn�a����:b�2&|KRޮ#6��@�A�J�N����i��ߢ�^��F�BI÷RF=�y����9g�|�蒣��W%h�MLA!c2%��6��}ŷLJ������O����]� ��JQ��)~S�/q13^�Z��"� 蕘�i���gHW�QY��eK+'\�U��Qv)v��&�5αG1�X99p�ĵ.�z�d��v܁��-�ahv�\�_6\2����_3D�CV5��k\�	_K���������>u�+�]4�H/�։S��9u��Ou�����~�����ZKo0�6�X�mc��8ި~���/�A��=�1��9.;s׳mJy�$�]XA��*��� ޳� i�a��e!ge&gux���KŉI-��p��hWڮ�[%"8��'���i`^�\�$��:�(���E�z��y���˄g�^*�φ�B�FVG�>b㥎K*��)�N~�N�x�<8f�`����C�D�G��M��#�:�`���3[h���T^y�vv�)S��9�G�K�hڒ�-�q~h�4"7'�`����ϾfZ1dzv�����֗�;��$KdL=�!{;!
>��oNIG&���U�?ĺ߹�Gp�j���cS�ü���_��(5i��f�pqlUuTˣ3�Y]���<jX3�OB�� ��!�)�&zN�btP�����NU����J�E�=�"�w����\e1��1O���_x���Rg_'o��{N����)=�Ff'��'�$���z��Ӑ+�?�SVx	E/�'^@xEex�AEf�?>��/�>�\�!�J/;���!��X�Ф0>P�0jRJB�˕)�i�8�Hh]��M��A����)���4��W�mZ�m�aS[��J NUq�3$uV�a�6�5��a[Y!���漺�o�L⃡�Kș[���1s�!`�n?����!�t9T�r2-;E��}�*H�AWЭᲹ~��Ǝ���?�ltN�?������}�)�OՇ�e[~5T1��^����~|`��K��Ҵz��5���Y��F��5��Ȃ�s��}@�1 �?�+�ч��i_��H�!0�3���C¥U�p�<A���x�Ř�a�K`�0gR�o ��~�V`ظy"��r���I+҆9��ԣ'P�!L�������6�Q2��	I�L�c����`�^�F�b?U��up�;N�JgZn�S�Sw��_cl-��LQ�D�����2"�ņ�F�	���eq�U���x�B��z��"�ɺ,`���x���뮢���9iN/�}7�M�3})�H^�A��dģ0�.U��� ?�Qp4�z�HO�y|�w}:��ǔc��f�<�A��^�(��GiLER����q$�UP/����%^ؑ �S��8�rn��sy!�4��+�֩�R�Lq{52;�Z�T��0-fA�����9Ͼ��GΌ��xq[��4����w4��o�-|l�Y�S+H�����6{�r�xσ}����[C�KL�$� Cp�M���?��li�?Ƅc���ϧm�32Î�B�Yk^:�*0�tS�Z���`)�������-�Ɠ~-��,s���&�rp��eI�x��G&�G���z���t;�Zya)7^��J��h����,���8�T��WJ�X�`H�T�!4W5/V�?�J����D�{�*qq�]9xM�=!VV�-�����z��mx����W��^��!��E������Pu6h��4�H_:�^���RÊ'z���J�IV�c�z�σ���V�aj�Q��+|"�*�c�m��$��`��Yn�	s�� d0z�^T��'��I�-ʠ%;�Ǯ&��4���1<��q��C��`s�%���.ga���)Bݚ���5�R�4l�.x�bg��N�>��3vߋ	�I���<%�^�\�JBC��t�=/;y��`����f���2+��F�f�@�΁���k��O�'��	6A���+&����2��#�����%aS�e�]�7&R�/$�-HO�Y
1ɑu��-�{-�U�qk�p��$�r�S�mz�:gM����ԏ���@4�B�	3$1?C��-�.\D������G��P~��
2r�XA���p���ԫ���N��x0��	��#s�rs�[!`_��%,,(ɁM9�8{��=��Ia�?�������Z*&�����w1E��Y�@��&_FL%!�����ܢY/S)���,9�ФBWo¬�P��D�C���fM�w��O-\w��Z�v���G|ʽ��Z���B���e�SC>鏣z�I��y�)u�R�u�$�,�]�,�Y}
pLt��Z:��)Ǣ�����v�a�.���������� ��ݍ���E�K�u��v=���8�X�7�t��w�-��:0

1(#��[K�1���,�qۖ�8��3 z��O,�T\��^��e��w9ă���My�1�U���
�h����x��ož�W��Xbt���W�^�����`�V�G�K�%9n��ʘ����־�%m8ॲ������sb���L���$��Յ7&���7����h��e��um/��
� -/�eF�,��3��51���Ɨ(�M��z�fX^W�,ɧS�7�Ǽ�� !G�X8���	�LUթ�}-Da���'���C�`����ۊ[�5�UwP�X#E��z�� MrA$���3c4yO<�`�����L�:�?���$̒?~�H.���V� ��N���&"*{7nj���m�e,7_����`ds�[Xv���,���!�% 1O�3�Η/�Sr�[�q��O#F��P!�[�8z�k]����c)��K���l��Ǘ��X��p���c��%�]XO9�[܅�w��ҧa9$�+n�C	��]Ќ��ӤK���'��]zǧ0���MR�1ޣ�����r�D�����SHΫCK-��{0}��J1��=Xn�޿�0R4����
Z�"I��,̔>ό�Zv��-�>M�+�+�1�4왳���S?!X����������v�!�P�
�T���U��"-a�I�ɢޮz���b��n���B�@u� �]�_6��=�Ł%��xG��O(k�="կ�b<֪s����җ��-�c�M��"C�$�)0�WʺK�n�7K�ix���]Z'r�m�JX������r��������輩�:L����>dT�h㯠^E3ǚ]�8�3�3B-��(�3yc�kp����=�����ٝu�6y������Gq���	犾�Ӱ.�4�	�HX��;s��4�;�j��}��٨�:!��"��~D���ۋ&d�I/1>p��0��S���E6~*��^�Ԑ@�y}���0�{���p+5�M�����s&P'LL_�tgy >�愸�4	s�in�0)�T�(k��x��j7��*p�z_�7�P�8�iR[����I9�wP}Q�E���vH�;�����*9�2�I\ӡ��	ƍ �8m��R&���۴XX3�?�Y����r���-��+S�l^ë�"@/�X �v��63�}�)
����P?T���I�X���?�{��ѧ�^�F畂}�XX�qD둗3o��&��~C�d���(ZnMhP�9�d���7�t� �����T���_�&5�ф�N�����������?R��j�+��oz�Xm�uhO�W�zZ�9���U8��ť�n��(��w)�[&����kܶ� ���NnJ r�P�ͬ�>h�l9����g(g��o�+�E�^��o+�D:jK�O�����폖
�${��xd�T��=5�9���V�CG�!�����Z�;�@)�b�:J.9�ć����^���td���r	��d��]�ƅ��|}�dt�ɋ,>���e&�
,�5����:ꨏP��M����W�Ҩ�D�*�՚״��Y��|���J��C2zw
�`�k�H��Z�H6ꜹu�������\���
����9��<��L;�	j���4�@_?6�/�W�M���'��HA<���zm�T�1�ȯ���^YYi��SR�	���Kcn��[�q��/ʆ��ٿ�Ft���	����&l��B} ��~����cN2t�rj��&[���.�.B}i�r��� d���(Qí(�}Ix�}CA���v�\LZ7T^D���;��g��$Mi���s���=ጕ���o8�t��b�p��We�y��
D�q��b-o_.%���2��H������E+�l��a�e�H&��ibޫ1�6|���J�ȱu�P:w�*�DI2���$s#���	3��`}��=���Cڨ��qK>J�#������b��>a�v`e�Y�2]�hfo�z w��[�c[�=X0��ej#���C��$�+ļ�q!	��u��z�=�w��g�	��GLR}¤�t���'v�y�k������^�b\ �g�O�^�1�(��' ��'=%��ޓ�y�w��O-?~�f߲/�C���%9I��N��p<m��,*B��"R���br'i���y@��#�Wk{���Pb�H�8���?@{LL"�N�����s<��q�,u<�e�g$��B�5V�ѻ���Ӓ%$��P�	�����A���B�E$ʕ,u�(��.+��3�$�hd4�pѝ���[fl�$�G[�2/a$V��$UB�p�G�5������<B92E˺��gX���AE���Z�b���=D�E�Df����;źّ�f9�[ؿ3���CX��V�QN;����O�p�?!�O�N���w�[3���3�:"P5X�U7��6���7Jp��M�->�}�f���:�L#�q�.�����@o���)8b�ƺ��ڗ��0��T�5��Uk�e
��J(��f%⊸�٫�	O1F�ꁍ����$v�b[w_=���*E�%+AB��t������3��mؿ�:ܚa�WǍ�tX3p�M_�l��V�L̄/w�B[�CT�Mŀ���CsT��y��3H��O�w��������&89�ߓ��m�ۏDs Y�)����0Zv���������H]6؃��*���E�y��C��ۧ�V��w�'���.��0�VV��E/ǜM)�c�&/t5𐒡�9�a�I�K�KuM��V'+A�R�������.	�3�ݩdߕU[p�������q�/kNb#MKʄ��P��k�PX�6M(A����~T���1��6���@؊h�'�F(��x�b�/���r~ܽ
��v���'��%�*�!û沯m�ܦ��!��]�Fa}M%'��dÅ����CɈ�$���A�?����u���\���y$[Q_��&���&C�����{�_�}_�6�ozƨ���m����Ķ�}�}	,hj���$�,���c��< v�{`���+�J�%A�e�a���^��NLz�Ȝ{�[�1h�]sT��,#m��7:�R }���?3�Ol$=���H��Z�c'Ҝ{��K��餁�(|���4��)�O]v��r$Ȃ��zE��$��c��M���&&$��=AU1��m�jV=��"���>_��%2�7i��Z��"@��,�Mz��'��P\0_�^q=��∉� �Z"ZM�s�2#���&��!ӳ^�D1J��`ꮋ��s]wt��ÂA�b�@g���L߂Ԕ��U��8dS��(;�-�(�/g��.��dL�����:��͞��.z���w����w38��2�X���՜;�i��4�=��8�%'�7��n ��ۣBV���3���8�hFM�>��ygً#��7�<�fW'��R^�!=VH+�-�,I�
��㢑�M�l؝�H?��y9�>slc��VW�����FbG~�vAm��|�:oh�M~��2���p�_��� A�[[�vqr�-�<�3|�4���A�W%�c�m�6@�*�jg/������MT��s�k{�i��'y�-@�KꭆB�1LM���RP��8�b�;�����l��+Ό����m�e)�~52c|��Ũv����W7,ᮟ�mj��*J�{j�_]b���a��,�s/��!R�S��X�����0�STk�l~
pB�|L���x��]9�J�t/>v��f���T�ɪO�5|���� "m>�<6e�]���x��Gń#Hf������V�Os䅥���bԃ	4�u�.��v�*��!�Xr���0?Tv�S���Y\ݚ�K�Z<"���;�������+�r$����Ϣ *�D�m�p��@
�I+~����j��,@��BL>fw���,�5�]���G�馵`���[ñi����٦Q3z.3k.A��-��"�Է�J�S�{!�ʇ5� ~ă��
pU�(~������#i��弟�8�AxI�C������g}���la_����:���?�6?eHy����TM��@Ə��ɖ=�sV`7�<ED�3����n-,�'q�u	��"\j�{�(㿤�@�eQt��Z��6v����4�E������8bʳ���fZ9����(�R�֛uzn9�׏Qq�a	`�nUmM��i�R��J\Z��&�q��e���cK�ή���c7;gk��1&EI�X��oy5	^7AgӺT��h2��I��F��p/�t��� �|��py���)������.�g��#څ���YoZ�&���_��(�7غ��GT����j'���IKJ-�� �*wS����7�IE��5Ve�¸�M��i����Ax�s�*�գ����=󆏮<>a�kO���ֺ*��H���m��/@��{w��Yδ�znH�F�9G<*|��3�����O�c
}з�%�0lR����`CA}L`�Ǣ�(|U�������1`hP<G{6�,$�8�����fdS��p������c��#�:%܋�)>k���M�T��{����J�4+�	�ٶ�
T���
G��}�c�R*�ΐ��;0��e�"�ۙ�r_�Q����#�f��I���6�lW�\ �|0�T+k��_c�M�ZԔӚK���+�z/k�Y	����	�C"륲�k?V��M��ΤKx��=�<�~��!�1hw��4=��������Ӽ�ǚ�q�h��
�n>��m���fO�9L��:N�nDD�O���׉D��y��H�	�ô
��b�J��T:�F<�|*X ����O��xz�5�`9I[�X�5O��3]=[����H�p���e�|RÅ�t%�J�A�����_s�F&2?i{!�S&��?X�D�=N��˚�^�����(�e�OݚP�r�-6Yc�8�U~��َ
L��I�Ռj��I��
Q�;���q3���E�?d�&��6na����5�{���Y=���e\���?*
}��H
$а��(41���D���)�Ͷ�V�O�I�D҉̪]"�e|D{ץ��Lׯ�]��ʦV"~K���;ِ�2ʲ1W�eFk!C�ϝ���m��u��P���VCUbQb�4�ķ�J����\+�f����>�m�Kk��
��i:���ӫ��� 8�9�V��s�JG�]�`G6�����b�$A[G/%q7�W;ϯG��|> �n<.޲ҿ�j|��#9�*�K�AW?g�`q �i5���N���@ؐ+��|ݭ�lͫ`�o�d����@�	n���iU���4�'��>D����a&|h�)7���)�d?F0>X�>$h���aL������"���^u���0�B�vm���$!V1��R�w��+�-�,�Ieײr��L�����r����6#��R���jw�d�\0���j*w�
e��2�+�|���w�^Y�A�3d�&���A簔Y{�kzHu�ص���J�1��Pc5�g�v�Qj_qH�uyI��R!Z(V�,�����F7&��z�K5�O�H�@���3L���9pS���E�i���� _8�=����<R�q��'�O~9��iW��5ʷl�T��g�uE �M�"w�Xʵ�މ;�'2ݰ�@Ԛ�C/�şJC�F6�l�!��J���M��.��o�p��?��)S�/�?��=�tC	4@��6�X{��[��_��uCg17T򊵲�4mJ��L�#�fv�'��=b����:Lp$��ZO��#�W�<������g9TK�
7�j>YI���&�ӲbQI�Z���E��p��r����C�pQ�ȍ��̒��5���\��Ca+��
2���Ye���Qּ�q�{6�5�t\��E�D��ɉ��2�U�)��5�	�Cf/�O��E����E���S��0�$��V�F(����A���+�Vs�<)�E{K��⣩ƴ:��k�΁���믄�<9�,|���������{֩$�<۫X�7�b���Sހ��A�O�!���I
���O�UQ�#�#)@BI�_�H$wW��~�)<�z^���rܽ`�J��y`�b�C�۫)�����8ZB���M������2F�V�h�IϹ�w�@�M��D���s�9"�m8��k���oR�~:O�M��Rr>C�\wݘ��h���~{�F��� ���K���ج���6�/3���c:���/B�l; d��c��nL�؅k�pW|����k�����r���$
��.:ۃ.�]-��z��q���%�Z�g%�Ι7�����K(,�p��R�����?��;�t�i�t���pp%\3��zI�>�<>ֲwj������p(h��V�5�a�_(�]q����ဢ�^�9[3�I�Uey�_{�����%��b���7u�r�����vYT�ӕ'���_j(�oc�[E��ꫠ�����B\���,�sZoL�i8*����P��1<;�x�!�ƽxTJ�.dP�
 G�.���W �u.�#������/и���8�G���NĒ�W ʝ��&�u	C�%~q	k�e��˧=������s��8{JԎ��X��D��r�]� � ��N���P�l?���Mg��:���,��%p�3g��J�)KfL����Cr��z�tbW��.G�.��T�������,|6� tb��1��R�� �%���ʂ0�[h��M�"ЧF������%w�D%�ѲNkV娹bb~���Qmes����I��pdD���͵��x��� ��m�,:a��Mb=�EX|��NN��8Y4��i�[�RW}�Fa_���f� p�:HU�3��`t8#��wF���
���mɡ�wF䒊 x#~���_��Qk1��D���D��z��+�K��D��b�q��	*J0��$}4��i����������0�B�Qߡ�mBV������Yq�D
�莱?���?Z�'�G�X#��K�;�=Ǯx�jg�BT[����lw!�v[{�~w��ϷM��f�"��V+���lYE�8�+pY�2M�ȡ:^����z�{jlZ؀���?f���L�N((�ƕ���/&�b�e�qe1 N�mdlV�v�.�ϴ��+�a��� ���U���<$�c���Ѵ�9���B�FB�c�r^��ŗb^�ND2�/��D����j09��Qy2�O��c͜�C�6�-[蟎*F����a8��2�2�.
U��� ��E?
;�ٿ} �)�dե����~�;\B��X��9��)�FP�C�CY��"��Â,�i�f��?���PN->o��_��1�t���˦G7b�E�`�>P��ɖ �CU�`/�[JQ�����#���h{�?ߩ�#��S�ZԻR@�	@�\���Ѽsj����B��o����x+e�����~�3�@�MEo4�7\����(�ܲe���t�w�dZ,�7��M�m1��m��| ،2Z��*ژJ��'����8��O�� ی0��%�׮���Z	�d��N+�1�m퓦�w�e|ِ��*"41E+��|�t����2/��1�I��1x�e���^�'�Xt=����i�S���y�+�23�0��
twW�FO�1�Q���b�I{hs�p�d�a�����*���G�%�Z�$݇Y3t�n�XB��[&�}V,�E�q}"�D���Xʠ�Nr�-�HgF�����l�)�YבۨC��ס���L�[��8�Cg%P,�����	��c��i�_�O����u�A�%T�Ǟ��0\ #Q��H�zt}6��$\�S���5��|� Fu9G29/��"W�Ǌ��`���܀C��<����_�N��'xX��HUі�M߿� �*�]5��!��x^P�H�����Α��ӭ�������Q�~��3RX��ށc��P�����T��p���������:�_~�r��pO\���[�������<�h��kc��=qA���'��T�pk^X�a�0 j|�D��Y�K>�Oq��Ta�@�5�1]�'�cr3Ǒ\��C�^R�Y|��`N���/ʇ�V�U�Z(�cQ�:٠o������4�Ē=�{��/W`��]�a0r�G��L��k�]f�HN���o�b~;6TZ{ݐ�G--|y���A�*
m�?L[�h[�ߤ>'��xڼK�i�N�Z�lؿ�]r3�U"]<g��Y��v���5{J.C�?��$Ǣ��'m�1���0���-&�tU���J{������Jj���u�� �X(e"��Kfh`E�����a8z���7��ٻ=Jk����~m=�8��o�Ė�(<\%c��l�3�ޖ�©��EyGu�N��������	�ۻ���ư摚���E��{���.�)֢�݈�����Íj�l�G���<v>��;��,J��	_?3[P�Z2͎7%6��q�V`"{5N�dY��6�>��G�A��\C�W��-w�s�k��'�M�kd�;���&��G��q�D��g�E�B�pI����!��ĕ��v+�tw�yv����%�Qe�8��Cs*I��=�)^���b5��,�>���o�k�5��e}�z�����T]ϑj�:�7�e��T�k��Xe{���W�N��Y=����N�D��ZYm��dE��!�6᱖���4�)�It�@�0/�kX	u�jO��j
4)B/�i�t�}��{�b|S4�o�/�%�²p#l����lI�5���T=�M̐w*~�"v�ҳv���g���>�*����ۧ �G�d��ʹJ1w�
^���
�vDn�KZ��D�G�)��
�\��Q�K������s���]�}���oM�c4���Q�����}��GN�|I��ӿ�hwh��2�9?�����|F���}��O�p:�О�z���	�I��qh?7��驌À_t�h=#�\���n��J�ka' K"Z�������E�]7�J�׊�s���`n�B�Ǟ<#�<!G�P��U�V���S���(f��V�o0��]v��*Jw!��w����׌�5��%����o� ����+U*��z�m��,��E2�<�f�F��mw'x�T8�3C���)&��m�N�ﮓ�x=c
�������y�5N�!��
�j�8I ���<����Q�@��V�E��w@���%�Ļ���ogT�Ed��3qR�<z�����cm�t�z�៧8tA�����Wnꙫ�.�Y�p\����	�t	^�k�l�\����-r��i��4&���&�S���^ީ~�J�l�<��1d3мg�^Xs�]ER��0��zD�U�~�88�!o�!�SM�
� d�����!Ϋ�	����v��o�W�q+��j���C��K8�Eh<��W�sm&8	 ��t��=R�O؝��+�22�oh�1ִD�ƌ�Z�Ћl!xЉ�Z�vV۹Q^a�g^��Ht�?�q��9��G��q�`ua4^"ۭaJ@��E�<i+WVYI��N�R�m�X�M%v�5<�cQڂKD����,Ig�J����ΪG�YyA� �����m�sBWe���(��;+��U�V��z�z�n���
`�×C�o�c&$h'��-6��]�,�>�K�t�^-gY�Z��+�<�d�#��;q!^V��cp�@�K�D ��s�3�h��46��?~����0�m���Bt2FƄ�g�gdM��ܫ#�����lk�z-�DE9��$Ӿg�
��^M�%�$;�w7����^~�[3_&��b�#����uѬ*�Rr�����9kX-��t�{igF�	����+����,��,�C\ZpGwc~������������.C��}�vᤥ��oDz"��G����2|R(�)�cTopWk� ��.�܃�@μ*I�����u!��=6�(PS�3�JK�b�-�QFJ=�"
и9:���H��JM�Ծ&�G��O]`�s:<��Cl� ��|�Z"
2gB u�j�J�N�p��5V+JÝ�{���LS�0��R�i��o]�ϖ��a�F~�	Svm�0J������e�9�Jg�!�uB��Q ����&@"�n�K�5�WEI�xJ1��/��jt	�䇋�$�6�4-c��?��I
T�#���Y�J�8�Mg�u>��J�{�Ŭ�P���`w��Y	[����ڿ�0����/�I���R���F��5t�zSr���5>�[&�9rʸ�aB��M2��=b�y���8�HU��s���f{L���A"�%���y���3�ݚ��0�([���;����C]x����q�E��?��
���eXM4����fC6J��\��4����Ri z>�)w�QWP~�6��q�~�U ��5�Y�߾��Ƽ����H�� 6��8ըaB�p�PO�Z�=6'��9�DC���"գ����6K�6������<���$���[�) ��@���+�5F`�C
��MR+��X�[�����Dm��>�d��[�V/�l?��f+ B�ōɹ�����ya�"Xu�7PN��:b1���6�n�/0���6��H�\t������ �z��S��	��%��h��hk/w�؞Ƭ�N�7�!�"��z���U^E�՝��,����RI���!W�����N��.��с���P�!I��,�E�Ԓ���;�(���C؇s�~g���Eҧo[�ׅ1~���(��~�&�/78��có�%�X ��#x��3]�`�2 �X;k&�/�xO|�Ğ$|N�Ig��#�y��U�F.����e��x��jQ��ذ�ͬ�� �q�����m{��ygl�S��R'R��T�V�B��r�֟Z9پp�lP{� �=~���`��]C�����#���Ԛdb��hSn��'��v3�y��T�
	�x�a���y�E%%��/(|!(KL1�q�`��S��b��5��/�\�_u�H�1���$����U�1!h�֤?s��6��LD�|��^�R+8X���(9`��l��4��������[
��}"�ҮՈ�����kP�ɸ�pvza��Hn�,fN���N�[^%܎zH��#�$3S��E>�<�\wW~����k�( e����'�Ζ��3��?���T��M5����F�w�=��4e�t^��qщ�ev��9Ӽ�4fTmreD��R�$���~j�d��+S���x��0�MwR 0��5
[��O����y���9~Z��3���R�a	e��#����%�B�l���h�wp�2��K$pS�[���B:����	h}e4r���ν�))����!��%����@7��sn@���4mg[�J���շ�8��������	~d]nȗ��%�U�����88���o��s�*m@ �(Xd�������r�c^A�%.�t�e�ܭ'Us���Jf;��k�c
UD�у�����C�}�ٮ>�ְj�u�Y�$�~Wu7h��ߥ��&U��kW#�t��mZ5*�uy%�@��X_0���س�e�9�
B���]F��U��vi��D;�0&g��u����;����i��'���f瑞A������Ԧͯ��p��H�����BGg�%�.��a��k�у�Ю� [סT(��vd߸��R[�L�J��?!뺍>��|`���i�hUK*tc� �FM.8A/��k��N�=Os���5�[�J7^���8�(:�����:i����V�bO�0=!�����,����7��'�����"�r*��Ư�QoT�pF��A�2����kh��y�V�T���;G�:��SA[J}��*9�*�C�R���j�O�59U�Y��A�J9!D:�=:��R^��
8�㔯I���wd�o���e�6��;e3xELuA���)�3E�k5dCV��0�'�"�ȕAJ{M�����}	���!������P�5��/qp�� ����<�	֤�
��V��ǥ�m���D'�զ�obPR'BtNW>�;w������/�o�[,����ɼߐg�eC>Mˁg83�'P�)-M�9� ��C;LtlGv�Z�	��3%�vE�`�!��q2�
�kh�ji���;2��C��$����ù՞���K�C�����Ѯ��c:��w�Z�8L�m2w����|���/�d�B:����c�j�T�+��&��OF9P�v�����d\����5�'��U�����ͺ���4��,�#��!�8�N�$�w^p�_���.W[��&�����&�i��Y���:��������'ۋ٬���b7Ђ�����$̣��)>��*A1�.+KR�T]����g�z�JHI�{5q����Q|,�z)e�y(�M���ľ%8Y[ͪ4m����|}5�	0"-k�r����l]��E�p�:@�`��-�Н�Е�����\P��*�؏�\H�|��r�Jށ^oyjj��Opy.�����!�3zW��q{�cty 9niS��/��[� ���K��KN�hǤ枵���i�uJ�F��;�,��TEAW{(%��h����D�t�=>�@5\�׉�C�C/R�
G���� O��Ĵ��8r�ix�tW� ���u3.�s��F2H����Y�b���Q7�ϞR���9@r������J��?��՜1h��r���6t�����u���`oe6.eH�L����l�lj$�g"R�єb.o�9*��4����Dmg$��ﶒ���� �ǟ�a$w��p3�AÂ�Q:����	;8.h#N� ���Ù�W�S�8]*_�Ȕ��'�3�����鐃�͑q�Q��bыg�E3���_��˼#�"��)�R0��:��	������c7.��=��[4�
t��Wh���K�m���?���y��u��l����Mm��K2�3Nb�,��N�.��}�>�^�؛7t�?��8���B����~
�n���rmC�BAc�*���kG���sh����ADÆ��#_�Gi�̫�"�֮λ��5=����|K�${����}�'���^��ƏHl���?�5<�#h&�g�.a"��S9�Z��D��u;�߁;!fvx��xp�j�c9�j���W�=^ϥ�"8dL�l��,|A�
�
]�G�s%��W�^$�iުW�v=qZ���$��*�S�Q��l0�a*�?;0���:���`X3D]_
�5=��hmFA;S�5N��".O~B�i�`胏���D��:��+3;f�?�C�"��X.o踿�&%+׽�M�(�#��x/�-�.�Wk�.�5�oYK
���=n���C�7�'��~N6N�?0�����I�;��s̓��������gН�Q��)�xN�j;2x�{2b9�+�W�u	�/u4z�����'�F����|��ŃU.�Cr��zi�+N�<
��~ ���i���O)���~���'4�T�y�N���`l9�-N�[ʓ'ݼ�Læ�V�5b���ɯ%Ͷ���]8=�(�Y�c�S�^[�{;$�@j-՞!��Iު�nyEpz}o1��f.�5����/Ϙ��٤
_�p�`��e��m�po#���k�L���{N|�z*t�6H�1+�=����P�P���T�"����fmlV.=O\Jo��+ w�j���CV�1��
�gV1R`�A�zc��rMŎ������ݒ�恷P�e������(H��[�=�G팓�Vj�^<^��iJ��O�|���Y��/�������_6���?}��Fg1wW����R� ݃���x3�,��>"�:S��#�O,(���w
��7>�}�lPx�|լI�S�:�ׄa�}����g��B� 1Z�,���) ��'B��^u9�s�{�`�{����#�ޔ-=D��E,Xd#)۽�H� �+e���a�.B���g��ϝ����O�_0���/���	����-\�T��C�$lwn�(+�����x�:UY84�k]X���"�@�غ�0��fF�߿[-`qSᢵ`�	�����7+�N=�3jft�;�,nt��`)���9�A܍מ����܇!D�o�9;0��b��o�{��;hr?����Լ��U��a��Ӎ�-x�D:������^$E�	ѯ�!I��R0��W������l��������[�je����f��{DԹK�����TL�3;Ve,&�^�V�M�N�����JA�����9,��::�	{vF\�C��q�	)�)��Wē^X?D�B�|��LÜ�t�(f(�S8x��2���S�n�6��n�u��N����m�/�<d�����ᄣ�qv���������E�C�2u��Ǒ{����ބP��^��U9x0�]��W�lk�6-l�Lm嵫��߸Y%�>��[�q����m*-���zJ7K�����ᨬ��%
6�����\�{T�
�;P���A��{�9��XO~������R6���g�ᚳ��QO<�S�Ϸ7P����*; 1/�|,<����� �hY+��:���:ٯ+P�5���MzӋ���E�a��ܸZ�>��X��@�:��U�q�=�@lɽ���9�/a���o��U'i*ʚ%�+N��f��3j�`1P.���;��]?`(��L�;RSs�Π�%������R
gI�(�B�V�Ojݘ�Gv��<�0�������[V�;��|J'�Xn�a�?�_��P0�`�!]�y���\�q��ŕia@�y���&�el��<ѣr�p�3��_��$-�+1��Z�Wo�P� �������Q��C��U��Ǩ�`;�~��MP�6��y3㌂F|;�<�C�i9� �.gY\���GA�[��f�"��,�~��4w�������^���,�}��鷮�=�ywT�617�����8<GdD��l��E���$	�!C�����4*g��hBV��`q�H�"T��B�NI.�U� �� �Pb���Bx�z�@�ॊA`v���py�q'X���(�{��I@�,d�i�_�RA�&w�DC��UR��CJKVW�R��b���L6O�	
�U��3&';W-/�g�a�U�ڶ�jr�m�%'d��1�L�)y�����.@�&���YΣ���E�� tH̸�<7�<�u�[-|lmfkE��	�k����[ʻ��B���w�T��|Sc� ����A˥ctiTgN1�u��L1`j9>�@���(�����N�YK��ъ"���r��X����L���.��V�/��,��B�y�5$�E4��bAߩުB��}��]�kK����g�Вb�Vଚ�Oɯ]��B��k���yw1f���(䧤kd��g����D�B�oX���7m6a�)һ0篔����n�l�� �ㅍ��45�-Or)��ѳ��<�Y�~�U{~3����@{�?�d���
��=,�&V��ae{���ZB�F!P]��YD�߱�y�k6���~�&7��u)��z�����E�A�x���8Ѽ�����hK�տ)��,��R~U�I��'�E�i���w�DN��3���vlt��3]���zW�̤w7�yNES��ElG��z���)��lq��bqYp�Hh�W;ٯ)H��պ��]���RR#�]JB�o����������2�^�ҟu����\<�<�;��zJs�쬼Æ����S9�V�F%;�Ф���n�Z ;���q$�6y���l�x��ʥ�x�;��ם���H�6�k�e�x9;��<��I���*�(w�(V�/��x����kc&��-dO:W�N��f�&��!P�JT��)۲����� E���մ���Eg��؋h[�5�4갮sb��L�va�%E����CZ/���6�c��7��A(P�LIa1;m�p6�Z�_����K�!1]Lߠ�p����_�o���{�4j�0Զhϴ�_)6{~$�����`N��t�����#8?G:�n��c�k�7m�1���δ\��|�+�H�Dߺ����C��,���Š�^&�$�NG�ڱk<�u)D�����倢!���b��Sk;����g�V�^��XAZ�>�� |!����Q䣕5��j4�K��'KeW���h�g�kx?�G�N�S̐En$�/ ����rZ2��7N�2q�@�s��[�9GԨĄS �-q���=W�d�,޶J��ة�*�|��Xq2�З��$��_��|�aq����zP�VV��]���� b=�k�1�i5C�.g[�nO�ъpzS�aI�;�P�KWĨ�C<�����L"�8,��eW��#�0"_A��@;��\&�� �3G}A�5�h:�� ��<f��I��Q��f�[����PX����C1���+P+Lˏj {���x4�&	4%�@H02��a�����3p6��&�$R}1�]�A��dw��^���7㸱uh����ǿ�k��#�Wȳ�H钸T
%%$AՖO����2M��#c���1=�@
񂊷}�P	�g.JU_� ���:�;v�ɽ��)>�x�K�M9yM��n���>���d�p^�=�-��[!t�+<u�=��� �M�>��R�t�0�'SR�g��g���&�[@�MP��Ji��`�l� �8U$Wm�=fjk��d��5Ƞ5��F��5pc�:{�"S��7�������@����A��)�XI��"�i[@�>
�kl+M\����lk���et�Z#�|��Ȣ2�`Ad�h����lV���"��D��Er�_q�sL�_ٚ"�K�N�=Ь����f���|��r,��nϑ8���+L��r��5�̟R[�7��LJW�t\���Pu/��%���K`�=�1T/U
>�us��2�l!z�Sh*�|C��Oy��%�݇��ãA (!�L�m qo�D-�b,��Q�*xI� ��=�{CI:��n �1zj�;9b�s�tg��]���bgX���<�Vk�	�V4e���
l�d�n���z&c�M��a��;�C"�b2d�%f?�o��/b�KK�DD�!�[�>��z �|u3}�(��e��C�X���}~��QO�m˜ԿE��]^ߐ~s1���(]i����ڄL%P��*k4��+��Y��q#�����&AL�|��g�c�c;��_H���s�X��l���y�ԃqAK-��^}ؽ�_�xgnĜ�p� \I6zm]�A��4ٰ`k��\�m9��8�r~�G��?������ ��e���䷳�
:��sg�"���[��Ƌ���bD�22g��l+Ehe95o`V"@�V��:�lS�2��G|w��@Fe�`��-!A�J)�P蒑^��S)?�����#Q38�{_��y�c��AP�`�g���HE�Zm��&���A�,�JU�mD	�c���4(�"��T��)���`~�ҫ�ZS�� \l�:����ҋ��R.:�K�@\�e߯0lw���e�M3zL�*W���oFs ALg^�D��z��~�Ȑs���t�Ӹ�-W6�rZ���:����bF,q-�y��-w͋��e�����x�!ٌPt���#n����^����vs����(Y��C�s�3jKE��@�"qk3�~xJc�J-��N>��p��Ŵ�
/�Wj�zh�0Kvŧ�%3�x�1�G�%X'd�r��pէ��Z��j�I��ﲍ=���g����i�Xbut�ʹ6RؾҢuQ$^t���8i~П̀��̼�w,m�0�I�]C����Z �O͵B��mƘ�dC��)gP�z�]����i�Ӓ���iqK�c�m�XP��}����.S-ő|ۦ/C� z�[+idB�;��������;_a�d �J)�'zRů��R&=*p?��{Q�p�*�����G(4fw������.�R�5�������,��A!ԙǾ.���7�?ė��-Gh�RJ;gAF��ǽߦn�h?T����R4S~�^���^T!~Ϙ�"$�.qF��<ۑem [V,�������hq{��6E�t�<ß��r֕:?KA�[�:�A*^�Ϣs����7`�s_v�H�Yi+��7@"y�;���L��(u(b�s��t˻��g���5l��&&i���(3�L�K�h�+
�8m{赼���^�*m�'C�P�1G���M��
�gG���� ����#C#m��Y���r�k��X�'�4n�y�c�G.r/�x:�]L#�gU��[�� ��S��3-��C���6�h�߷������ɵn��T�"����ڐ�@��&���>K--�\�P�-�� Qc�?(y�j9�� �yt<#.��#��`�/�����1�l�p��>{@YĮ=o��=�(�d�a��P���J3~�5Wp�,"�����z1g�#�����J��#j�c�,1��+a�P�,�s�˛�$�7*��Y&���%j�~Y�����b׆X����,�c�=t{�#�_�F������-i ���RxT?��+�9�Aހ�8���|��o�����v����?2HW���k���
�oW2}����*iU��W�s�MݳP�g�]�����Ж�����l�u�3�Ԇ
*6��v��F��ݳ,%�Ƌ��%���������E���:X�a~�~�X���������M�ma2���%�L��`y���Ȁ ��������^���fH�\xѸX�%t����B�'¡����'?�u8>�2n��E��T��cNc��?M?�������BK�I���n�>�p2-��2'3?��C�Z��M8��!�ǝ�V�@�s��z�s��_1r� ڋ��2|�L�Nښ�t����e�*%�~{�b��bә�!�e(��|;��JW}�$ɸ\��,�f/�q�Y�?�q��8H1�V�%�k �X��1D��#Ia9G�k)��7��fY�ͤ\+F�v1lA��lO�ͫ��E� �À:��cȫ������1.F.a(G���QxW�V5�u2h���c��"d���qJ,���k
GR���	H�7��^����t.�q�T&kʝ��V�B�$�������œ�����Џ0,�&d��c����|�ܒx͓���,��0=	x'�%�l��\I�Ó��H���f������-���4c˕,����C�5
��^B���Q� u�\�9	!^\6uj���Z_�������k�����#ȴ_���`�Tc�_�q2뙱�!�t��:b�@xA1�;�	�}N�[Y.���S�s?�'S����>R��z���=E�*�)Q�
R��E������K}8�5�|�hw�X� f��P�%養�@���B+��.��yA`�Gʳw]�q�i��9F'_և�G#_�3źjz[�U3Y��quN
#�$ƌ>�J�#?wVώ�a�� ?Z�/�L@����M��t8��>ǤJ�R�ܒ�Z=�]�#V��R����/z,�ӱ�JCc9FY�a�@^�X{��V��)��*��z.�ӳ�Oc8H5+��ubs��J��(Z
Gb��b�]��cB�`D ��@���?>.��|�E��ڶX�Q�{m���nRh����9� �Ir/��V__K]�q�1-(i�kٺ0�GzbӺWr������2��B�Z�N��D��B��T� �&�]�m�O�y\�'	ڄ��_�F�h~L�(��+ Y���s-)��N
�����L��TC�(�4�����k*z�ڤ��)3f
���� ?��x���0<raHgL���9�s��_�ϡM(d�7�xv���WL��\���߮::P]��&�lh��:�9��8��z2s���"YsԮ2�}�y"Y�,Ij�#T�v�A�[r�<���'��������Z`���xMQ!s직sf�U}��\�E��H�:��l�O����ʈ�̽�!V0�0A_��͸��mN���v���L��)���T�S��<����@]д��7 <�090d�ɢ���B�7��Ju'II��}7�������f3���EwzjΞ��Z��uv����{he
.�A��<:�7�L�s!(f�W���a����QR���s���o4w弶�j�W��O�	HI	���� ���<R�ι(�Vϧ��8������94�W��J��¯�B?��X"����|w���|�< ��.��gǜ	K���$���	hʢJ�=�`�kɿ����i�հ���f�h�f�߻Di~��z2@���ۖ��&����r��f��'r���߇�t��,`�{+5��U.����K!! 2p.���FøAІ����9����?�� �Y�lR�5z	��'E����@kL��Ҷ]�z3إ���T��Z"�O�Ԃ����!2�O��QR��U���N1I
�[δ	z#*�����m7j
�U��c��	D�t�kQ��KO�,gI���_��;���ɳ�'��UJ7����ؽ��[b`�	.D��Ӂ�Gֽv�z�!�= �<E�tf�c�y��V�8�<�b{�8�~�e��Gc/l�MP��߱�u��0
�4?*�p�G�l��������K�.�ݙy'���˘d�ܻz�?�U����$��3��&.!��:Ȏ�ޡu� 4�I�;�ьU�X��b��Y �SF�4�cN�5
�1�*y� ��[җ�3O�b�Wg��V�\�c��M���8���~�!)��tY�!+�xL���[3}Ղ�@�i	C��=s����tqXO���`暞�g��*���RH�GY�:o��ZU�D����V���;U�Jya�8����Y�ԛ����^�>h#��l�ˊ��߻��k/����(�*:Tjndz��]�����?�B�����Q��?���o�i��>�g�O�o�ج�W-qW ��'L"׏�ʅ$f���ͩ�C�� W+�J�+�=J��?�C��g����}���Xܒ)�R��Z�˦�M��ȅ��Bz+��{��Vvjr%*�}�$k�\� ��,�ڮ��ݿ_�������]p��!O���ِ�E��I�4���z��F��6>�z���U��ހ�5i]�1�ɍxuJ�e.���X���.&��?p$-��Ŭ��R
�E��w��9a� �3���q]~Ӂ��L���9�@)�68���`f�|1���J�?�W�)����8���3�{~<YSZ#Ɉ�2R�m����n�ܤ�N�8�R��q�BJ���Rץό!oQ>
y�3QV���[�o- �T"�f�
%e���9��y�㒟Z�ځ&�����K���|�wz���^a���fmH��ۃl�f����3i[�nI_�
G�U����re~������X6Eу�W��qP>�����ƢeUC*f+�L9���J�9
��*����ޥ3�ou�Ne6[�@_=�� �� `	���4��Ç�iMS����k����`�ў~(O#8�_[�3_�s��B��Z".�O`l>$iT�^C�H��C�#��X��ch��0��s��7`��Ń��|����twgǟ�am��a+㜄��s��lp&��;�&�l>��B�������J.t���Y�$P	�rܳ�@&�*���yᔔ67p�C�!h�Q-�x�����}.�5a��5�ɶ	, ����up�w;#=�������b��Z ��;�g�{7%q*�Obr~F�h�X��N��?�!�e�^����B��1�<����;)!��q(���:8S��l�J���m`�t'�8��D+H'P�AL�� xI,5y��N��ϧ9�>�5n[_�,-�m�p�y1h+��� ����)�^�cYכ���Ts'��Ė@��T稇����M~���9��g������mi��:����6Jr+�W��l����',���c�=Ik�����`M'ܙF�=�pb�\9�G ��Ƒ�f�^xj+�چ�(��F�v�E�J��x�XY�2�]dB��'���H�F?���Z3"�b��#(�P��},LWU7�*����{�����4�/R�͟�Ϋ�N�?� #?g� �e�Y
��WEׯ3Iu#��x~Q�̜R}�Ru�@��B�5=�$�:����b�dd���7�������bSOf8���
�8>>�V�Z�'̆S�Q��ggJ#�$�18Z��#��tz!�2��3�S�ZM���N�����SKdڶGAڹ��nR���\����<>=�k۞i�i��T>'��D㋽��NG�|��H�: ��!�]� ��9��9I���`�n�Dv x��Nj�t M��%~ ����XS��/�{@3��Y��^��!��&U�������6���o�����r�|+B��!#����G�rh�bfaC:�����w�Y@��	}4�I#Њfk���z�7��U�'v�����mv>��"c �W��=�bC���^̒�ǝ��%�[.;_֖��lhHڱ葃(����0cŮ⊪����yA��%E �봗��c6|�'������	3`�+O.lf��0����+mPc	֚�֒I�X���>�l����u9�j�⿻����Ē��f}��9A�= 0g_&���4FX>��c�+�\���XT�׃sjѶ4���;�3,��0b.~��̮q�`e�C<<�R���v�s�~țз($����:\��⎇{�#��@��t�B�?��I�Zo$�mI0K��i(�(}���s���m.�Ԓ���������@�z��k���/8��}�HP��Bxj��Ec�v�4suZ�<ԝ'�!�p̕����"�	Z(�6e���a̝}�1'8/<�I��' �pE�$˺_&h7J�NX�����9kQ�P@�{�`n��RK��,���j�������2�\QM����8W���/C
Wg�IUS��ç�hفo�7Cy���0=|�_R�Xp��5����9e =��w��=�aD�L�@��h�޾���=��Q.0����T�4�E�r�$��6�J0�*��Հ��Qq/ٻ�Ѝ䛮3/y���S�/�6mRH��;������S�1ٙ�mv��r��"��8��q!�R�� ���c6_ӓ��,�߇�����o,��	�v�#�8]�r��'%D 8�5p��U��.eI`�5Zwr	.������YVl���!c��"�U~�Z���8�T��s���s��	�8� 6	w�%H6�t��VT�Mw�$:� �yh���;�5���v�#�V��jr mc_k�U��V���W�Ө���t�|�譮-�=37~����k�>�_�"��>�?N�(�:R�t�'[4ri���b�w���牊���%3U���s�/��f���;��rդT�]ؙ+E�c��J@w�f�O�_W�yf�M���`6r~�WC�!r��{���`�m*��ӄ�B���+�:�ge�f�`vuSk���Y.t"S��B��>�H��ә��K��/�S�%�ҩ*����i%Y�0(֏�=�j��C��+F�%���R���j3�Z�p�r�s7�I��u�h�7���[������
+��Ɣ Ҟ�/=i͠Mp���I��Id�vne�{Ӎ.�_�
�?�!M�ߠO�����.��|}�۞����Ϯa7:��<�WG-L\9o�Ig_�O�g��=��k��4���$���On: 1���,B��=E���-�E�����@�4��fl�	�^s��ۛp��C��y��E5$���)3|\��ʧ�i��)	뼐z�ѯŧ�QIL0<�"�y}�����E8���[���#)ET2�+���b��@�t7�S�M��	;H�<|v����dy/"��7#�v&�������v�Iuf�wU&�Kc&�d5����Ve$�5j�$H��~C���1�sR�z�����1�l�V*����_M�^h/�9>F�;�f��&�JVX�m|v���H3��#V�H
����	��q�f����f�q�~έ����P�<?���긨"�N�'_�b�r���~j��ҏV�����haEX:�O�گ�zu�*����ol�4�OZ4"K�o�$~����������R�f��&H*s���)��B�Ӭ��j���٧��g|�:�7o��ߟ�r�S�$������lM��Pv�(E�A5��U���P�x��2���*��߲�wb��	<<�\6 �����_�RS�\!	r1;��R�(Օ(��s7ڲ�a�	�զ� )������.��2$�t��v,w��Ԫ#|vW�TwebU4un��j�7�9-{�I�ȏWU��㌱�	��,cӟi��ֱ����&���Z2x� kB�����҂�p�T��E�,m��J)wk�2�-[In^��� ���ʛ�q�k��/)�\��\��������"@��yT��JZǎ��u:C?�)j:��9�3=g�1�_���S8P � �9n�kENK��L�!�����n����/9�`\'�)ٱ%���'*��r
o� ��P�Ԧ}����h�G/���Q�TԂ׍� M��-�e
|��WY�tɁ���YКxwǾ~��w����ӏ�vĖ��+����k�Z��f�ɹ�`.��=K��h�d场�-�Zp��PW���<����~�j̥ߖg<Gi|��C���7 ��n�9(����N�;�Zd���I�qcyfɣ,�����g�\�����%�'��h�dCT*+��$���Rmt�V�����H=}cc�o'�q�g��l{&��7��Wo$C�k"��_����M�$$_��h��AN|ր�.��9�wn�^��2��-a�r�M�'�n�vx��8������^9^�4wε��d��<�ک�g~�������?HK�0'u�Nbw-��0ڊ�ҠhP5}m����O�럖e.�gm�jX��G�1���)HI+l����	M8�	a> O!J�D"av0�2�7�be�!E��BP�%�'�&�]/y������y��~[�+��>���'X<h�JkaW�}kt��F�U��̉TQ��OĻ�ȈA+C�p�����;^��pt������1* Rk�?=�h���יXl��D*���&�!��W����r�Cf�M♟Y��9Á\l��y�η�ܗɺ��##������ N���`�e5\�V-�zC�_Q4-��;r$�(�Ǔ����>�{��%����AiU=��Q8틕ɴB�I��ɝ�� �L�o������S����]�(� �F>�IO�y�Z�'k~�^��x�駮���q=�'�:�N��$��q����xs�A2���`sJk�n�~�iw�핂橅c�Oh��$BP ��@�q�{m���E�'i�L��a~����t0���[M���V��a�@��8�����bT�b}��;�^�(c���W�&w*�
X�7@ag8"�%�ǲ4��fA�<D��\�ې��ݢ���8&�"h��D�n���&$ ]-FP4!���<�������!��\��yW:U��-f����K�i�%#�n�YMw��.�^C�T >\�!�쟠�)@66��ҫ;GQ�x�[��8a�k~fmΣ�%��� e̻<µ��[�>��s�����s�(���D��g�G:�dp7���l^n�E1n�#��b��`/���s�_�J��ߪ�c]a��F@=s��
}9���z��vg�V5�����U����W8oFA"�7 �Ǉnw�F��=w���&����$V�]��`) �g�n�,�N{���k#^��VD��k-A��5��Dݪ�}^���\bH����վ��hO5�
1i� <k�7��a.,�@��U�uZ��,�$��os�!�*[�e<�8n�0�HH�F�pͭgdX?�*�f<"X�MV+��RIͽ�P�rB+F�8�G;В���̋������u��۬����M�c�j�xi����u�N��^�V$�*��LQ�I����}�F�J����ѧ����{4Y+Q��H��b�QlL-��a8�Ϛ�6,�[��:q�W�u����g7�u�e��I��k/&���f�h'c3lIϟ���w��vh���w4���X��QG�Ͳb�߶P��Z�cD���×��4�8�)��O����!F��Uh;�>4�1 JJ �Ә��CyV^� �}[��s�o6��V�3���8#䁃t��p��S��O�L߿�����9fYs¹�����և��u�GAL�����{B_�;�b}��%s�1~�Q�,f��a�n��4� ��u �;�
t?@+H'kW��}K� <*]4������Yv���ٲ�g_Us��MkXITڍ��GW���K����-j����/�!#׸~��j�� �ET4�>	B���L�'��~R��px�� �S��ȋ�蘚��\i��A���l�=B��W"?�~ �f�n��)�Y:�e�v"۹���xX'M(r�Xq�=�J�t�o�H[�qx�R�G!��Cɯ&kY?vC�z#w�����L�?G;*�G�+���~/���l��	l�A�׳CB�e���olsX\�G3C����ơ3�|d�V�.���'�5�z/~�]�� {��\�aOY��P@F�ً��{�!��yؤ�ᾖ�|�K����M���[���MB���G���!�د�W�@�詔k��f�.��Ւ�M�12xe������=��@.����9���0m�{�c;LT������=�G��rA'��m�4^;gL���Uc��'*�@kd[�.{�5�7HJw!����(�Q�M��!�[�L)���E/Wvk0�6c��/A���<y��Em�:��B|}��p1�SB?E|?k��:�-ȏ�n���\��P����z?("�K��{���a��@P�C�8�y�l�
 ��J�8�lj]�e�u?���'�#�^~�wy��=TZx&#�����(��9�)�����O�fk+4�e���?��}��� �K����[�)
q�
�bv(���+��kw�:���n���5&��q~�T2-��(�4eц�}��I��|��*��rΠ��S�y�w`��2���'���^7�A]UG�_5�|KT���A�א�����Gt7��=�mމ�t�|
����y_^��:[�<gٯ��G;nn@���T/�L���R�n�)��)G8���u~>�&�Ҫ�B�$pȊ�y�<S�֣5��z�r_B|)/ꈏq��pT��&pj0�#d��)X�L.�h|굹4]�vW�1����B8���<Dm��O�<9�DqRR�'��k��!$߁dTl$켺E�����k;�D90+	��>�p�p@��<H��ʠ�b���ym݄s�hB�"
e�;�/T�0CE�K!�@h8�>�Q��Z6!�cFl�����>1�PԾ�:�AV�9w���$�}�g�Ȭ�z��B��R�N�����K�~��Kq�KE;�u@��"�:9�Y���I9�4������+�����	�U
{�\Y��Bn>��ҙ�ģ��2DO?�R�0e�N��ճnP��K��� ]�_�	}Z�B����ˬ���YL��Xm/�ٳ��b�VT4�C/Fpm��5�L,f31-�F]N�"@R����p�4������8HM���m�gH�z�(BG�$��H-��S���$��!��]n���34�72� Q��k�Tw�gtԠ���[�3��	J�Ѷ$�2��B0�?u�+���!�7�k�ݣ�< e�(>�ҏ���u����MX`���'�p�z'�=�s��P?*z/x�o'����v����H6f.$�և^�Э� ����=����Q=k��^��B���1	��Q��M�5/��w호�y�]�Ǯ���w�C�{�|>��t��Y�|Qh͚".5�"Lo|h[�K`�7u<�1m+�1T�b3U���2������B����\p!������A�ZDjkwu}�fZ����/�#q|��G�o��g�а�	��n`�}�0�q:E+��D�{$j�Ҁ�D�y�%̃5"]�	w�^��M�_�a�]��P�:�ը���ڵ}��ޣkx�Y>�
������V�h�l�{DnZA�g�`��`�i�.�o��kD�Kڰ>.��b����	ͷ���,�c$!>�<�8J�az��'��Ҡ*�$D��萮�ɀ.'$#Qz���� "Yo]W�;��8#r�}{��!���+��4)������@B�;�D~���F|���h��u�A�	Z?/�z�����fGJ�8�����W�=��&t����]K�V�w6E���+J�@�.=�qT�u�~*��=񲶌��C;I�v%ݟ�O�fq�X��3q��=��NN��\	L��b!���6$Y2��\j�����S������"H���$1�4l=D�na�|��H���b�#���y�)E�R��f�$Sm�.��Q�,�inP.��Qgд;�}��݌w�oIά��/�n���n� �e�C��2�3�]e� \6]���8�L�$��V�0�).��_�ͮ��m!h$5o�I���Ƶɓ<�AQ�O���A1F���������(yi�~�gm1��j�.@\���n����u�GZ�M���r�K��l��u� ������dv��n����mgD�|R�`�	×�
ٜd�p�^�4��b��l�A��O�a�������Qz�*�h�����#����J�pW������0���LM����WY�x��#/�d�j����=����V����v���j�9�W9�\��>��&���q���(X/rd׿�{�xؓ���h2h`�k��@HI�w���s�Ce>8;�~1��<��c�������K�0I���zk��4P�����ũ�0�6�7���ߨ�8N���������ۡ5����K46=���� ���HV���¦��B2p�'�>���fkf�(�\)Y$vk�������^��C.;t��7�<j�6@#�i&p{1=V��%����9�`T�&х���q�(��1�8�nk��R�4T�}=SWF�3"H_��z�d�$�1��2+�B�zP�2���e4�:��ٕu�F�'���z��;��|��N��A ��W�\�7��}ZK���)8��kuD�s��y&��?�ɶ����<��%F֣�dp��)�?�Z�f}� �H���MN�Кmb��O2��J��0���TN���+L�?�H_�WwU+�[Q+��_P�F1�݉DH����,��K�4O�e�J.�C���������_��X�
XZ���[�|�qI���9"+�
�_ުJ�Ev�h籄>���	����k�_������4�A���[U������qM�!?H_2n�&�����8�j�t�p�>(��F�M6(]d�ݙ�/1�T�d�z"��k]3�%K	Q�>��%���.٣j���u�]���\o�$ݵSTp����Y�/��D�J_�)S�,��O���M�2����-�U�!Is�NLʒ>�I* Z��خʿ��x� �l,m3���ͨ�T#�a��r�����3}�܇�L;^4��e�~�i,�|���F��B�L�~��T��M�������暍�Ŝ��Z�����I�����\G�~�+/����]	b�.kS�s�U{}�2	~�k�Ϝ���U�n%��= ��6̡�Ghw�΢D�ጿ|p�U`*x ��Z}w� �"��d{���Y�G���3���B �.j�7 ()��˱πW������[��Cb�����Uqʘk�JO�dRqt6��FL?����A�?K��ߝ��T��B|�-k��2�:����h�ޭ���J*�{��?RŽQa��N *���D`�K5�_k3����L2��������Pn���@M��Ny	�z@W�7ï�4;~ϕ�̍���	��K)n�O8����d.��S0��Z�����"69�)�Z�5��.kk~�^7�����)V��~��p�j'�I���S3Ԭ�j�z)Ol���w2�gYG�:�d�ʤ���Z�7|� ���] \~��WnĿ�+-������p]]=���M���-`êL�xb��W�g�����dHm�|ʾ
�Sx���z������lԼT%�ˤ�
7��~�#����>���<q%��1�p�7�M���gF��Gm 7T�~�G�|�h�?6�ۦ%��L�ta�P����lo���c�T���!��
"�O�#��wDfΥ|�~�J�^p�J$y|���n���q*��ڂ���TY����N��v�*��k�E��?b�J��&�}��"M��9��m��O{.4�gv�������@x���:ط˄���q�_��1f����lF��5aa*>��o9�r�pꍫ�y��'�6\�w��C�j�p3�[9[��sYaD����V��V��ӏh
�T��z5��22�?1(&`���S�0kn�矇g������MQB����,�]���L7ޥ?�ã~y��`�\t7L����C��v��T#>*Ls9K��}��D�5+�C��őy���5��u-(��n�_�Ʒ?�"︴'�eTDL��a�O3��ȭa�^!��`:״sb�� F��W=��|��/�o�l�`f<y?��eZ�v(���]>/�#���Q�:��3���g�5M*b� @���q/���}}����k�oP���E��?��>�}׳�:X�Z{Jq�C�+�9ٴ@�L]��B��m�xB�_ѓ���5��-�Ҵ��,nT��Tz��tcX;-B��g�2^�[ul��5\{!x7�)X2*AN#	L)�U	�5z6n��1$a|T)t�#y��16) ��Kɋ�3kn�3^�d�{.�1]�M*С����+�FT�9�r���(�L�k��j�V�6@@��f�{�$W&<��-�s/����١!X�,e	W*���;O�$�-��+���c����Ԭ�.c�$d�Ȏ�#\��d_���m�AQ�gL���v�P�z��eB�*k"��H]b>�cv/X<*�w]�仠^&�3>�]K4;T��TgfV�S�G�� �דR��������}w�2�e�Q��X�~a��%L�����)%��S^��H��"�FH���E�a#$�s?��X�N��Q=S��*��~c�ą�� ��VT�`(m�M�2�@��҂�Dq�?S4�
Qŵ1V��O��n&]�p`�n�|����~G�����^P(j9]0��8����mW=�q�ŋ��,�;��p	aP)_?a�=C,R�ϵ���<�����1�/����&�XRJ��o|�4oW���7�u��0����_���9ը���]� `�RRLX>ټ_�ڸ���#�h�~�(��5�~-Q��ަ+{[�F�4�J����n��줦:�>*o���������������
r���
40���`�u�O�h��(�>{�ՎGs���]¬�p�f�o�4�ݴIE�,��B}0�B:ꤦ�β�'�&atKju���`������~ߤ�w�ܹ��1��8'1���P�����a���/�̇�����Ǹ�**�Y�ob�+��=���J�:�Y��3M�N�����&^��Bw�r3���i�	С�r���r+F�����d����=]�{�R|e��u�~ ��0���ō=y"�~�#F��Y�k������f�W�wOr)���`S>j>�2�8��i\��������Do%��� ���E����eB��gp$��E�*�r��d��w�miǼ��ín���S�<Ԑ%T��&ߑ�W��������9�k�&k�fV�4���
��9��3|ck��{����P6�WD+�)}=��83��O���<F��޽,��д#_�$E�P����'�!j�\mD�!f�q����-A.]����H��Ŏ��2i�Y	�!ǲ�&���Dr_ɠ��*�
^_>��s�Qi�,�I�X�Z�{�h�eo���st�]��6'lGB���ɳ�Q2
�w�޿��"�lb���[7�`����f�}8]�m���M��<TP��E���zzu�,!u2{&,�{�ԶU8������Z�R`���G�.��R�M�ҭ�!pA��'�/�kH�~�v�$j��߫��V6���ʂiF�R�O.6�?�j�����c�b-������2�����������i����R�,�	�Ί��'Z$I�ᮗ>�O髛4���ϰ��Q&�
��&�'j��t:�1ֵ�Ҙ�A�[=,I~=���W�<I~�#�ǲx;���xM����&���������S�����
1�T�9Ȗ��̨��f�%�w?˕$�_����$�o�ߟ"�*�]�/�L\�S�:S.�fH~�4`�6ߜkZ`�6�w�:�K���~b�+�Op�oE����ՠY[{��u�eB^?JV0����r�gv���b�3�����fy[�����`�2n�N���o�|}�1�u|0T^/n��qu��76`�w���2!�;)��۠�4��κ-�3�����4a��ga��mx��:�O�fT��8���&���%�R��yb,�=�&>Uު_�|�wu�^�����p�i"��60z��|F���^)���B��z&�}���! �j��v�F��N�j�L��"�Lk�%P}��9T�r�6`��f�yu�w`'��(��Z�dT1����gT�W��f����Uڭ�GG������1I����
����u�.�!Ւ�^(|	��Y1}b>C�!Op������'Mbv��2�طϲ�=�p�Y	����� C�é�D�TG `�(�\���%x�U&�"�D@ȵ+����7��	�#L�t6�B"e~�g��- ��ԣ �fA"�\����K�m4G���,���M�������M#��zT�8�׈�z�T�q`�R֫#���j�Ҝ�,�O���Ü4�*Ql�sRU2����%l��y3��х�Z{�[R
��X��o���v� �[r7h�)�&&��}$l���2��+�� �rv�3��s�]�2�K�2�����6�RR?7Z���B�v�e�
]F��.�5� ��ֵ�q�%��T�V�����0���"�g��"ʐJg?7>X󝉥xAܜ�`��@y�.�z�7�T��]W��M�$�݋����O!MȘ�L�cf��q[�[e�s�# ���K6�F��v<�33z�7u�ƅoJ�4D1b�j�m΀�iE�41�E����W�BHLԜZ�"�B���w���bH� ��hێ.�k���hX�DC���s/+�����������>�9W'���S&R��<�o�BK��E��52��	�1K����E��H� ��8��;��9ǔE�k>6��q�	'�����NS%g�(V�q3������'�V�c�x_V~�6�@�u�vWE��Z���3|p�^��`K���=��r|+Ve���Ŵ���㩢>:�A~;�J]��J#��X+!�[ �Ⱥ���CH��|fл��}�ع4I�g��4���F�.�Z�&�v���/�_�<w������t�g�� wSh�bY��w��'v���2Ȼ��?i��h���J��Az����V(�Ρ�����Ȩ�>��,ŪOM��1?p��A�ʂ��E�F�
b��@L���<W��Y
d�$�\�/J��qy>�,�(���V�p��ո�J�3=�:������:贵�+P�򅞂���&�\:"�
ؾ��%|�g��e|w�9m���ɶ�����?������*)�rZ�&���|�~�/5_��仸!s�������,pv��g���^�=~�^�+��׍rw�W*�_� A,�+��~2�D�U ���=��iګÑ,S~��i�ΪTm�zW���'K���Z���CW��&�d��g�j������f^K���,tۉTw�tq��3/+?B��?0�bi!{��T�����5!l�,q� ��ڒ��b8yomr}�a�N.���Z�>^-�g0V�uDV�i�
�ǗսR��[�0�S��~Q�,�5Q8˕���C��K

�g��o�h�����1u�Z�	`��/�N~C���M��Nk��A��g�4M��'K�5x��S��_����y�Ϻ�=쓊�J�B��*Y&��̽� ;jg�R��_Yː%8�7�t��æ�B�iC��2n��ڒu���ԛ��;�jڱ����W�(1��c�L���?��c�~��>my����8ֳN��j�d�cM�E��R�r��!޷M=��_�3V<��6ԣ���ڊ%ƦH�>o�ٽ��?�jtmLۡ�B%1�;�}F@��<rK�>g5V�lµ�<�5Z���� �\<e)�K~E�`L�ǆ��!����Γ����?�<��\����\`d��4D��)��*�n�-���3'z�J�Q�p����$���1@��-p�[&�)D��s�ʃ�@��Y���� �R��W2r[&�G~�F���ju��˞����cy�g�@��n���p��
�ݭ�xI���`��_Tǟ,��g�:�D��DEo�ֻ�Z��l��]�Z����
����K�=�N�o*Zi�=<� �����C0o0��O��35DcQ(*|IgUDټ�'���Kx~��ҵ�CHo��Y����˰8��l����`�kk 6)��D�z�3�m��D���w> к��&����_����,�-�<���m��ɵ�q�K
��/��] ��17�dEv�It�5�7���5.��Fo4�#��}=���7�wT.�1�Ws?�V$<c������. ��9��9�v:�{q���ٞQ��Bip�$�/�X�y�<C�h�X{���c��2����B��I2�6T���A��K����ܳ�	}��3pB��*�rXnc����
�?u]��n3��D�.m������>�m+z��&ԉڍ�nu9U�����趱t$t��V��4��L�.Q��8�k�g񵼱�G�K�|(<|m��/ђ ,��PIު�/¢����{��T/gC�]a|ӗr�����&��Vv��E�1oT�ۻυ�6��n�)�9����U���|�͜�3u�!��}���ĥ@-A�C#���$�^�����*�M}�\V¢���9��E�d���)��v�Ͻ3F���\�a�~�X�څ-���V�a�E7d�?y�<<];4��E;B/9_"��m��'���� �w�s�7�d�����4��:'1w�����f�X�)�.p�fV��2��a`h
F�̈KP���&���I7!e<�(��. �(愥Y�w��b�ՙ#:�D.	؈��!!�fr�^|��N<M���Dm���6����#RA�K9G�Ȏ�6�/��sz����Cm;:|���䊱�U ��Yia�!n�OD��$��NvG���DU<ˬ��A������߆�jL�UB�����ާ�+]V���U싯�^j�/��W`��r�t�$��U�j��	R�z��H�l}����G�X��k�P��pl־Q�5!�3�V���tN*E�~
@���#�%`SP�)�"�	g�R>�^{Ė0�q9j�=�C�Cw�}8uq����*�{=6ˬ`ĳ2O�!�6,�y�P�r����ƯD���Z�ih@h;�cl.~��+�-�M�цc�"�1�f%j)
�K�%*{���
Hy��z�QT�ɧ�^)pT�>�����3+� ��2\�S`�RE�sbk���X��`�Y�{�B�^������x�.�b��o|����Xٿ�"�7^V�"[-i�X�����>�k"���`G"^؄��b�6��o�ڧ��}�����^Kύ�ᇁT�8!+$�?�3.��ڮ�w��)� �y��GN�O:R5B��?���0����:�]E�c!�;�^fȠ�|����rƝ��{������ǺӽI�D�#�������y~��`r]�����C��o>@RI��a��ت�C�F2d����f"���F�n<k��g�&X����#=���c[J))K ��~�jҋ�!Mh}�4��nP�Ji�5�ڵ����hU�R����Fb�u4���<q�+��?9�� ����NҚ�C<�9�d����:R��凃;Ή/�fa,�۔�C���:�i��[���:�t
iB ���6@�E?u��v>:�_W�vد�Ai'��G,���a����/^�L�WD�z�۱�[�8�gSV�:I:̬M�&. �w7RO����B�(���M;O9��#��9�����nd_�͂����6�� �2V9&���1��x�<����iBƃ��!��%����8A�"�?�,�|��:�T�R6�CqAi<��I<���A�Z)nL	[��fü���Y��O�E���[��R|��̛w���l����rf
��Q{tj�Ϸhs}ȥ�d������5�b���@�5Ӄcg��٢��x�Q�1Oȹi����Ė��i����(�B|Cz�z�P	k�����J5���ko��� ����z>ژ��ڧ���4}!3R�ѹ\`LBỂqܥ����(�i�u�\���$#G	FJ�l�q�������9y�"�����M�vN���<v�����zͅ�n�1���֬�j,Z+����o8�aZ����i|���m���L{z��0#��t��çS���w�Շ.EsKi���:C��0P@҆�Ͷ��!
VjGZF��6��4}�4� ��l�`�\��'MNnh:\\\/DG(U�5m��X���j����{y"����������&��PԞBA�˄��.�R��T��k��������P��a�3g�.��:�J<�\���2o�c�W�D���<�]��Rodz���~(j�J�`�e�L�N#�MbV��.�S	(Ƕ�����n�A�Bi���ȩ�*�S���|9���X���nf`�HߏfIQ6Ă J4;��[�P�N؊����������!˦L1���.�rI7�~�o]��0?����p(�5��˼���2�:;*,����MNp�-�9'�wȕD>v�ڞGKSڴݛ���X�������d�7o�)JU�Â 8(D�E�i�%�=7%�Upe��t�L(�;(�����r����R~R��:��*�i�����cP�L�b������UvQE����Vթ61 ��'�=/]�5
'��	��hG��:�J�����ME�.Sg���
	�9�""�װ��5���B��[���h�e�X�ٚ�/�~�mMY~K�[JE���lH�g�>$���V�� bH	��A��p���պiؔkݎ����\�w9�a���T����V��E9
f�y�e����̐�+�j��Е9���W���Wk����10yT��ܻ��yX�$�N��s���������0t>1��K�#g��*�T�/��}�^9���R�4�;ɔsb��" Jk��;z����x;壶�o�GA�C�����,�HSE���l �77h Ԧ���9��0�P�0� x�&���͍_RV�E͌����b�,e�yt�]�&�W��fa{:���Q��k�E�^J#ߎ}ޖ)[Lw6�}�;�E8�}�9c�Հ��|tݍ߫� *�!���+�74,o��Yc�n��5��_��>e��]�W�}�ѫ������R�ȣե*J�F1��Yn�4��iV�\�-sy�������>�I��Ӊ���C���#/�|�i�d�j�	�����q�o%���RW�>u`c�;�:��\�i=R)�X��HB|����=��*��֑$��5M^j�sp�Ϥ�FXaO�o��O��W���"�0� ���K~8M�RR2��'�#Q�*
�ȩ=̐њ~fѭ�K\X{!�S�.ȃ;=�{���~�}3.~iTW̼7l���Qwjc ���G?�2��X���\�Ds�q�3����n��a�O_��D�j2�x)�~B<�!��Ee��G��L]3bZ��W��<��HV�2S��
b������-�[趉ef���U]%�@3��ܫ>d&I g�s�h�(�� �@NN���_ؖ# ��������R�����Ae���?�c {\N2�A.JʵT�$��moa�|����<<]Çi���#���m����z5�u�-� �QC��	E�:�B���F�	=��L���Ht��;M%ϗ�P�rw�#�R[���@��}�Ē�,���:���Z�8TV+�FGe�sR�Ø�hQ�)qd�m*�{��V������<�o�����**C���h��nk��˙����մ:�a(�J�򾚈oɣ�fp����v�����*��}Gs|���/��>%v�89��X.iI&X��0H.N"u~�����`|E��7-ܰ����[�2tOA��A�b.�I}ق�T�k%���s��6;� �"K��J�GK���5F�x��i}�<��r��\g}�8��3�r)A|���2����т*��Gy!'	Ռ����%��]é���,�a���հ5"�)��A�Ng�d�Z�4�`��B�B���M���$�4!WX��`pq�M"��-�N�tʆLPp��9�Ք��*Д(���)�Vw��um�K�˩~��m�Dp��n��J�5p��$a�Wo�2�R7o��d�;[0/N��:`�� �ҷ9 E��o���~�
B�����z:�SƩ&��K�|��)��󑗁���9#1����t�k䳙�P��w:�SjC=N��9��!��$w�g�Y�}N�k�4���J�-�0N�;@��m�q�ea� ��� {b�sEHqݢ�P�^��F$?@HP%Ј��r������ߦ������w�2= ��sACZ@�n����F ��o�y��'�ƹ.�}��:�+�����͑�.��(���}�5��C��P5٫)�d���gV���!�P�4P$�\�"K�^����N�R��}���s�N�����O�j�I�=p54J�d�����p�Nˑs��a�AN�LK��+^�PG��
�S���R��54SϹl|��4����PA�����ê��Q�|�-ss�捬zV���1�p|U5B�qT(0[^��4�+�����x��������<�\�S�<��4;����$c��m�N"�w2�E���f4k?�?�vڂ˴���2�ȥ��P�$�q�-����C�)3q�/5�wN�F�e	>�����/��"����jE��x
���-q x�+e{�8$����R���)�:�w~�+{b3���>ʪ;�����\�*�]��׌��೨�3�(d&h�{
0u�U�xw�E�B��tU�f9�����*���Yj+t�ȥ*��#gK�w�A�̻b�A�#gE*EI��D���3TǑ$B�??/g���_:��=w�5��}mvqv��\V�=�G�˓�һ��8
tn����TsT�&o��Q��� X@FJ��z�I�&JV�U1�d�C� P�i�[�}�:����O²�Ŧl�����ЀMi�t;��$9̰�����k7Q��^�Q���XϞ�z���E��J��ٝ���Y�D����ҍ�\�k��_�,�Es���8tbn#�>qa����炭$�.1������?#<�½����8�(^�E5��U;�$��d��8�[W��^�cS��>��3�U\��\тa`��9��Xy�=P�^#@�'eo��YJtC�_�.��¹֯�+^ ?Y�n�s���.��/��K
�֞�s�z5�V<{Ʈ��+��,�sq]��`%tq-��'��?�s��W�@�%���4�"�$Ln�5���wq��r�QD�Ę�7V�q�r�DL ����c�d2v�t�"�a_��o>e�
� $D���͑8Y��4�f&}.l�X��wy*e�{8����5Y���p�3-�&�n��p��(�0�W�e�^i2��!PNCi�C�WB�aLRJÔ�ؿ�����\aG�w�L,}�\^���2p5�<DQ�-�}�g�S.�'ci+)���C㢪Ԥ/(_I�ȍ���a4fNA��-�/A���� 	�7 �
�7ב,�&��O��0~AWW��w�AMu1�����T^mҙ�m�������A'K�Kl�T
m�T4�_	U�ӯ,������Af��.yٽ��A�0�T(c�����T�&�F���jY� �c���T,��|@��#���\+ �E�nM�S�l�Ӏ���n�9wQ�6�s#�Ń�O�B����I�.p�X� I2W�5� ������+���[l`<��)���;U5J����:��� �V�ckr�������aY*���	G�j��Ax3���ꅻ���|��5Qۋ;I�n\1��\Vb!x CL��B⚋���#��0�,|P{�Q� �L}��� ��L7��p�!"�]����������ٜ`�l��4�%�%G���yJv0*L�c'2�6'OX6���_�L�2u�.� !��.���������
���<Z�$\ׯ���spl���t�q6��p��4���f���,�qpnj� �z�E����t�F�\8�Ӑ�F�!�n��(AS\��	��јX.J��?���@�a
˄moP���DҜz��e���@�T)��q\�@10藐��a�,�P�@�'�D+�iAl]�p2��Ϩ�!��9�k&��bf�|���ۼ��v�ƶV���'f�&%�6��	+? �q�ROU2��b!�v����������!�6CMG�qǨA[���L4sŧ�!=�9�c�X�`��� �ȼ�+��9�a������I=�m�qT~�>w����aS�[���	�8;�I_6�_ �;JkP�1d�p]�RUSYM�(`&i">�'����̋�z��)6F�����eK�'
����yG�_3�D*�5i�3:^�L�mk�(T��ͭ�e4+���m���-�>k�ڂ҂T����|NU+�g�ybӊh�m����`;T�u.�N�Y՜�]{j�#X��ύ�)�R��H�A&��>�xC�b�T�9J������TA|�V�h���(���:q$�����P�-�ԁ�,r�w��N����	�s�E��M����>��Ŧ���Ʌ��l곭���	�f���~ә���(�#��S�����S7�Nm,JR��JbI�C��z��K;�6j�^H*Q�����fA����,$�ȣ�KNoe5��W���7�̟S��$�����>�GC��_ك��Z��� L�}&�3z��l�8�K�B������㉄���՗�N � ��됣�S�q�D��m���G�^J��͵�<�8M̀0�6�q9��F����5�}mk��E�������UbBn5��y����ǒ�q�R*l��F�
�.kE6����!�k�]�~PPxzEY��qP�8Sp3s�\)+��.H��T�~�tF]-E�����/����"'q|j��2�I	�.gN���R��ƃ"J�0s�t0M�sHqϠ�7��S��̚��uF�����0;vN� �Gm7?�"r�D����	����n�:�����ƀ��Y�Ik&�
d%_�:�� ֒N��|M�Z
8z��R��6b�����1P�獦���.�Z��eCIς�
eτe-b��S��^��@\ν��<���nj2z�,�$��s����h`ai�:��Z�� ?#�M5