��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ���������������$j5�3I�uc[oH1sa?�uRG��D�#ź
��,+c˶��F�J3I�ֺ�f6Zؒ@Md�o��?¦Q��Z�^�\��l��z��K�g1�KM���y�%ǗD!��̛{s�1�A7��S
�($Cpy�㜧(������ޟ�[m�P�00;�! �,��� j}�����:��*� iɊ�w�7Z��k;x��-1�@�@aO�\& � 2��޳,��$��}����ӒMX�p�"Fj'@��depK��;k5t���\i5�0�Q�{��7Ԍ��v���(bY�{�o�#�0��2����/�zz��Ե�FB uz0)%8�&��8N����U��z�ġI��!���@�ߋ�k����n��߳-�@T��1La$)X�޹�eP[@z6���nQ2�:Z��梍 �g^j���XS��e���q��A��eh�h�;=���b��x�k�l|3P�/y�w�wᕗ.k��,��C����\du	�|w%q/�o����J�ܤ��t+H�x��gw��I��T�$hhS2��6&̦ y�q��h~��\@��,?��gD�	��������K��@�;Ů&q-Ʀf�o���H~1���q�Bo�hh��t��ӽ�� �i�������]�e_�&�dyW���Iѝj�������;8��%�NstD�L<�p �8N"s�����S�������1j{i+��q�v�O��P	5�- I:���2�
����1�-���i�5!�����v�1�G1���b� ��0�S��5t��4N~��ElB��H52�\KQ0lg2AI��g��Ԍ��2�Ik,Q��O$��7&���y07fa�QaH��Ɠ7�e�oI���3]Q��o���o��tv/��ä��Y	K�p��%�	m8�vz⩿�}�o6�ee��3g����Y��6��#'Glk�7¶������Ã�������!,�t��S��) ЧQ��/?-�)ލ��<Y�[�vF�N�~��8͇T��:���f�@��ǘL�XbNNº�,X��錩�ꑅ��w(�J1+UPv�j��^�x3�8���wȎ�j�7� ������;��^����N��F
:��ۊ�է���?3�u��5"g)�N6V�H^���`����� }gz�	�U�5�[UD���V�ɡ341����#vi�&�G�(j�RZ!���T��.�U�ċ6�������
� ��K����f-��ߴ���V��M���$�Ҕ݄lmZO<���L�:�-S>�U_2C �w���h�� +��ؚ��Pe}��V�G&��-�bl�
T��i�����vN(:V�Y��Q���F�j��[������b �?nA�1+MY"i[����}ej�ƣ3�i]ʽ�*4��Z1rjh_�i]��G�;9 ���A3tqjT/_�`��p'�dEf,�ǯc�7׸��Xאz�,*�:�30}���{��+k'�Jp}�����ꢬ6cL,_�m[-PLκ��HJegg���d<����Ѥ����f�1o(�0<#f3�9;��nD>�8�+��I>6���Ţ�������Ѫ����E�F�����e����� ��_M�=j�d�nC��G�K��c�/؜���ׯ@���S.��b���ء�R��O���2��-�1�z�5��XI#�)얊�9���Z�r��#�kaVM����ݖ;uP��i��{�1���o��P�q��+q�ѬJ��+/I��¢� �c�cx�s���;����6��W�1�KW;CT�i���M_�ֿ�O���s��Hʡ�(��=�0ـ�����I�����H@ᡲ=`�6�<�|TY�����hB^���L�>�b��HF����ٙ?��V�x6~�ũZ�s�j��0#m���}4v������c�G339*t� la���L�zQY��Gޭ[0��.s�ך�)����y8�*�VB�S���hs޸���b�.̠Ҿ�wv/����7Ӆnh�u?����yx4�e���Ye�
&� �	/�^M����]ԕ�|��kF�1��`�6��@��d�s�I]6W��53��9RS~�\uu�61��}<Iߦ�	Q��j����1g�T����O�],��	�Q'�"�s��h��.2�|l�J�U����Z��M:��zGk��@���T^v�Ro�qV=��cp�������Q��焗�Ke�T�	�����Hr�bH��k�?%�r�<D�X
�p�[�P���J{��?�R�� �*���l��y���>�́���3�)=Ki-ɨm҃�3)�&���(���k��Gu��Ɣ��ٍi��q�ΏßI�y��l���9x3X�?W�Kg�f�ṫx�N�7ܧtx��YLk�����r|a;H�m�@&�~U��\ѣ����9�g�V�*-��eD�7�)	�'����G��Eŏ�0`Hfdhx ���)��#P�E�G��N_x��a6��hm{W�A$ٌL����. �����n���Z�M⿩qܪ)�X�#�'tBZYK�q�g*׌�o |q%Υ+�Ӈ�f�AR.2����R���S�ve�T�dO�itM۞w�X�)��T���*YN�k�J�gH�/jh��Z!���J��62��g������{�{S�Y�F̭+e��K�MO��J۞.��U���\������U�G�[D�d3�~���c���A"��133d�C�<����F/�ׁRE����X�p����qc	��EH�[��T�-����ߥ'}��,�y��]J�+�n�� z#���>2�xX*i<^ހM�=]kLW�]���v����AQ'GȔP���9
��8��$�^v���<��a�,!��t:��>�v�"�aiD,d��;p(�0�{�d�"?���P�0r��D��P�F�� ��!�n���]�T ���Kntv5-��I���u"b|zl��7�5@p��N����(d� �Ixa��
E�Xr����mb�V������<%
t��n ��[+��8'�g��7�C�����F�OR���Lz��Y�����a��*�ߢ�y�D5%�����G����P%r7�iNU���
�_�~��eq��-P�Rh2���.�U�|�[���
Oc{��Q�9��|���)m`ڧ���*�JE���X�i� 0�~���0��H<�dFP�-l�v�����+m�\��n�F�{�5X�+,��ѓY}������<zA�猜��Z�ܷ�J�*k�{�$�Կ(�~^r�]��f��Y��#��#��?Tm�yG+�jP�2��S
�"1��Lxc� 3J_b�AB��'.�>�	�I9��!��@q9�&6;<D���i?Y�z�������o���������!$���=��o9Z��"���f�5̻5r�*0G���0�g�\H�&ME�~�_�����Bx*?��bY�d.m`�+ǁ�*�.����9-/�eu�"f[���%��z^����)�-����C!+�^�P�P.l��C(�� �7�]Q�)�%F���T��sC�ԥU��?��uJ�Gdoʻ�vK�r�攖%��L�I|t�F��������=�J�(�584����՗���k1"�R����h]%�h##(��,��&|�xTW�
��qYj<w��Y$ �p�3>�z���~�֮�Z���1`+P���v��s��xX��q�,�>��j���e� XA�6���]2X�Ȥҙ�3�O�8����C2��7;\%��_��k�`!�2Ī�!݇{����~�I� ��麦>�q(�rl�׻�����Y���oo���xo��GG:�֕
	�B4O̦�Z�L�?�I�e59�k���}kU��ɪ~�ڪ��P[@����
�}��T1P���M��Fr����c���΅�!Ԡ�{�[e�}&��~��U�ճ6�[�$��S�$��Tr�_�?��ա�������]��G�����K.��0���ǋ(�@6+F:1N����I@oԢ�H�����k`f+3��6��w�d���f�`y�>���n�[��?9up�ׅ�����e��n�"�z�t��2!U8�̌��O�y��g�e�8y**�3�E�.me�ɯj��SD���|�Z�k1 )L�		��a`IɅCs�"2�W��`>���a]�Z�z�غ)}=Z>���+��gB#z�C:���OE8��ܑ3���
�/ۖ���������
>vD��['�.d��C��6O6�ƫ�W��Z�pYw����\��(���O�]�z�y$���M�����qlИ� �\�G�����-�KԳYs�>x������x�a��,�������1R���Ʌ�������K���Lܭr� ��Wz1o|�!i T���V�� F�14P�_s�:9ME_�rAX��!��Sn:H;��`ɲuЫ2r���Y��mҘ���_+�����ǡg>���^�R`(�b���N�	ݡ�X���[���Ռg�������JE%	��c)��{�T����ޙ	�y�V�]өB�xh"�I���5^L�.��ZG�=`����+��fނ�}���鬋^;�BU��������l��MA�]-��)�Q�_A!,�ݜjA�j4|��X���U70~NU�G���ǻp�tO��8�D��v��	8���}$��x-��o��(=�@���[���蒑5�~͜�l���ܙH���Y0l�;˛�0P*MA8� �o�<��)��3�9�ePp��}a��G�G�O-pnZȮM�Pc�ڠ3,Э��<,%z�O�V:x *ﯶ�R���aL`w�ǯ_�־e��W@���M��w|8�6��Ml���V��z�X�I���XԐJ4��G�}��`�M�q�g�ab�3��
���=<h�K'� �7�]'��1�V��D=�q��$�� 65���N��3�3��Iu�5�zǜuݡ�tԳП��_�2p�7]<�T��8�