��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�#&��#�<������::A���� �\�7�ݡ�y׵��G^.R��C\K�xef1�SDs����G2�km�����I��
�[��-��3�oX�by[���_K,�����J.ċS-���Q`�oS��{�������2���A���J`@��[��Io
��e����CQ��I����;*��%u�l�j|���x�����3I}���}ÿi)�+����#�̙�4O���<*{d�kfz����P�Š���z��t�Z�}z-�Sj�넺i�:���n�|a	�ZgҖ�GQ~U�F����s��)�����.rR�,$�+l����㲰j�6�oǑV�sjNѽ������.�0��8 sHZڲ�;�?b*��w�U\u;�z�V�q���!�ρcx����&����� v�@���;m�F�����U�����;aC�E!-n����b�F�l. �cA$��ncg�n	@��f��A�R��ּ��5��"N)O2�.�NX��U�ljzi,�
����'�Ғ���U��]9�5_˽ V���(�%YppzC�lS� @����e��9�s��'�ړ�Tx��JP�Ib���~����P�|��6��cI���aa�G�@D�J����32��&�!GA?a�,)�;��w��u����"X7���B�F`->�����p&ay=U�+�W�]qw0hJ�']���ub��ޕ�[��Ɯ-u���&��a^���tc�  ]�)���85����� b�"]d�S�2͗_@��,���@Of����(R����m�Vr׾;�c?`߳��ٷ):ѡ`�0��Q/����z�SR��q�.�ԉ���l0��s��a�Ӽ;���yZ3<� �0q��wx��G���Ju��#wY���M�2&�OA��ou��F'�U����E���I��-8&l�oz��X�G�ȓ�4ւfՉHs���Gܯ֣H�}�~'�e�B	���⅘�ܐ�b����.�^��۪��G��5��h*�����g�_و�<F^6?#1}�S��|�0;�_�N����|�,@�VuQ��:e���/Y�1X�D�Mm��7�<AZ]����*�A7���|Y<�:e���sD1���a���$)�+}̒�f.��&�j<*EbvGZp��n�E�tZ��4���T�.#�R#
¢��<׆���� l�mՠêr��@�i$[e 5̚(��c���uļ��m�60J�[�n��߷�'���keL����l�痉�Y�#-7Q�k���Vy�G�W�«v����(�,�OWQIe��N��Q�fa�r�O��
��b�Ÿ�QL�Hc���42hS�X�Q��"�~����RN��G�����f^O ��"��'�����{�;�RNN��)<.2�d���0���v���v�W��m�ޖ{�/�3�%S蕚ͫK��C�h�M���L$�w�1¨0��R$kK;��u�e��P���� �Kn`qHS���4��b,�O�v�ɱ<�&��H�����h���lw�ז%L.�G8"�]8����IR�=������f���K^�d����Bp�N6\i� ´���.� �)x7!����Rc���S�Lx�4G��E�hy��򥙼b$���*�5������ �����-��a�6�P�<`��h6��Л�g�	xC�A�jS��"���~4b/��d�/�j��_��\6�l��O�rJ�P�q�(���K�%4����-���_����/,z�����r��=­y8�Z�Q�&.B�o����X
�����ax��Gp�����>�ػ��jL�v<��q��$�<�U��S	~P��M���5�y0�r�u�b��J�?s��c���>���zՙ�V'����W�	�:,��$L��&)g��f�}ע{p�a�^2g�����.�O�HU��}�\g��JZx�Ke7���(ٖ����)&�*�@��Q�ˏ$�=���Q�)Ix���=�z����I$� �r��C���4Tgq,���OS�-!Բ�u�Ϭ����0���0�p[Ʌ��H��*��*�ȭd�(�N����3�@�)]>$�v�|�c5JS����^��Q�k4���>��T�'�m�9$1��I��h
�Y���X��X~�A��z�wZ��t���X^���Ғq��+"G�x)ڡ�j�\��`Ό��;�S=���$�o�����zs�o<�Um�mt�P��h�d68ݮ8���G����j��,�& �}�o�1�|7x�E����)aό=�"��:��F��d5�Ɩ��^	f]��v0�(VK�Y��WÅ�;�-M����(7$)T�E��1<��Z���U��A��x+S�Z���z��Bv����º�	�'�w���[�o#����JfF�9:)=,��ō=���v&�a����b�-���V[�M�������� ��u)C���;�όN���9����Rd������$/��*�ŵ�l�܏l�]L�f�O@Kv9{�����R�w��x�;��]�c^<h���Q
��nm!�!l��^A d�G���lRG�J4�l�lcn{3��8��\[\b��E�x�^V���Ń� �#�?��;\��,"�`}����M���Ș.^�`��V��|�����es��������ĵP� 0�d�f���o����5;����=.9"�l�
�"E�%���I��#ٌ0��������,X?]�㕠T�QxOf����0�x�P]�s��7��2U���G.BJP)�c��@Z~�8{/PR��8��t��J���ꙟz���9,1T�K��Ѿ�_�(��f��Ć�y���b�aL,����7�Z�ly�Gá�����?�"�v�8�la�71h��iZM*�����7����#C�S��ߵ5�6�W��E�Q��3@�.��NŪ�oL��n��_%�|���}`�5m���X�z�.�W���-�{�0g�֦I�
�W��h{6zWdD$k��Hr�k��Jѡ�-���4͍��
��`I/�|���M){-RĽl����k)���s�il��q��9M�ґ:|�.|4s�*]f�g�~���B�� ��0�VЁE���'�W�'���Vg4���ޞkʜ��M�D�Eʏ�)�O�:�咫BO�{�-qy��~�2tBJ/Hv���&(�	M��C>)����]	mwn:
�3q���Фh,T�7i��r3�5�m��=���&���Q�˾�X�EE���{Rε�
C�� z ��µv�bg�/'���^���R2gUm��Y}V{姭2�/V�9)��ݼ�qQ���֪��qs�ҠLs���Z��5 �x�oZ]��j��{͔��'�YN㩄�K�(���@eƾ�1s8��9HW�^Sp��\���p)x*d,KR��qzzP���`Cִ�Ǧ�I�3!���-�.��4��V2W���ڔ��nR���Sƾ��){>�0.�����nͲ���s�"�J�Zjf�8+��,.ҡ�ҩSY�Bx}&ܫ�8�䮦���g��T��]�7l��\)����]�(����ʐYD�UN �`"���7��Κ�+�`�m@OoQM�w�uE�nNr�M��g����Vp��{�A=2"<y���`�]��s�0�3��J�Dd2]^H !�� .ond�A^h�S˦� @��VD�,��;u�y�e�_-ty=w�b':�����>������`.�'���ܡ���.i�D���O�����/-w]d���t�bH$��y��.��k�t���Q�ʀ|
�ӯ>Q|��3���W��*f��7�kd�f��8�Z���r�m�� ���%�Q��Wo��o�ml��m�mM�1G��&��)G
Ƥx�����=*::vrt#Ļ�}	�ɯ��1��W󝥣���ؕ��0�G��"gn��2��b�����x'DH>f-�bi���w��U*X��AA����,�����#�����a��E�4E �	�J#�0Q=$Vl9j:��	�Z۰_m'
h-]Z�Ն@x����������zz���ء��}���^8���d�v�	����� ��yQ���BI(�k�AT-�ٻ�y�xt�I�J���F#�K˭1v�f����F1�ݜVP4�".^6v�F������Z��I�h���JP"	��`Տ�g�0�:ʐW��Gͩ�z����ф��w�W�Ӵ��ԃ�W�5�mM�j�̎����W�AO/9y{�����X� 2C�u`���a`y�hL�\���S��R�P�VW��Y&�)V��d3;Z�1�`���]���C�x"���-��é�����\ZK�-RA��y��?�z�lE��8�	L9��mA��c���s1	g�5W�����˒H? Ӎʤvÿ���S��>vzQy:$�AeY���9�Bԭ`�^Y����[mF�����B�%��K1k-��K�>��S��~ۨ��rD^������N�H��Vn���;�Ԥ�ӭ�72�R���-���G�p�;���#�#�bF�)E���!�V[|�W�����e�e,K�B}n)pZҗ돪�r,���!�$��Rʦ�o�t[�j��]|?p~1�Q$Ѣ��E%3��v� -�,�楐�*�r����7	���1��x�$,Oy'����"A��RB��C�������oGk�5R#�[�<wI��#�
�c0��V�P�+3�Z�_*�T*}�'����@K �'ڦ]�cn��Bˉ�*�4�C�z�=Ŋ<)���8�� ��$z����E8Sz�v!Gg�vh�ɖu
�.I�a�=I�����g�f�+Y��+7���MC}����ݧ)q��(Ǜ1�6C��T��F�u�S�;�a+����" ���c����p�&�u��B�T �,Y�'�?ѳ{ѩ���	��b��P�·��;w=�����9�<����~ӳ�%mq���.�-��L�@�<Q�"T�?��j���7v1�т���b����0фw�D��~8���3��8������@��4c���������}i�n��J/�)D�$����u&�u��6�d"�B3��4S$OF0XV\YC�״'�/w�>l��9�1�q����`�'���w���F���i�@����Zk�<�K)�&�>�D<a�w�k�����p�k�F�a��|D�DA���l�� �񪥐��4�dv䜇N�\A�?+�Q[oZ ,X1jM��E�[�ܯ���o�4����,��_���Ԟ:�Iǟdշ��[A��ku �:���z���傔U�����.�rI�F��L�
�����Q���Υ��N�]l'*ޖXlG��In�t�����Myv�鶰���)k��Ϭ��;}���F��-�Yc�u��S����=�:̿5�Ԟ����t���E[Ki��c�ލ�[�'���;t/�LQ���-B\��c-��� �����O�ن�qeۑ-� HT�����Ӝt�d}��f�EC[�R�g'�9?���tP>�X׺][Ƴ܀G�TYV��ոΝ�&����{�&V�7RW�i۹�P��M%O@��"��*'�:�J�d�TWu��'��w�M����p����f5;�7�3;����#�&V+�|\��l��0��s��ى1�+@MSkI���b�(ǟ_{3��>���ְ/��j_��%cNW?E}�Q�R���3�(؀�������U�J;�xG�->��LDR�r���r�QT��N d廭D)AYq2KW�5��/�U��F�x�7�b�w�nE�E��b�[��!d�0ص@Lu�7���gq>ڞ�sD�Opߋg���Ꮡ�����~�(ƱՍ
C'~��LA3�KMsd���
�w���u5�Z�Y)�+�4,T�F7:km%v����Po$�;]�Yz��Y:��yS�	9�4�l{'+A��\[���S���ٔ,��p1t0un���WК�����b���B��T�o��NT�ףy�.��� j���,����L�1&T�ٺ$�I���<ɾ��w����$Z��"�9�2����|<��Mf�Ofp��0]S�\"9�ME�����I`~]�s��k{��ir��RY��� �=N�Н�0.��bn����駏��\�&h��m�A���#>�@q�P��P|7��P�����?R��1J8Zr\��h}�v����;@J����WY�7K��@u>T3o�/h��ap���j�����3�R#֒i*�y�����G�����T�+'5h��NZ��z8�ٍ3{�/V��W[�{���ߴ�������w�X�QرM��Lͅ��gg�*�ə<�;r����mLr�|�U^�R�(��n��1�=*��p�|�8�y�E��;UO��\�)��O
���.~�l�����g;���5/�_xLBҺR�Z��,��Y����*��J�s����t����{G�/����ֈᨁ6���i�S!h��~g�fo��L&Vi����Ѷ�ڸ^��^���Ԉ!*"P(��̾Al��b�.�c���3�e����&O�۸WJ���7
���C���<�,!�[�A}އ/���/4DH��X���_�UK�X:ԺX@q9��\ꈢrJl����x�M̬T��׷��Ց���Uȃ}"�Ѻ5�A��z��T���b�|��89@�c@MamX�R}�G\�[�BAߥ��b��W֗4T�y^3�M��f͉�����]�?A�����5m��a'�iT*�+�eҚՓ��ULq�b���"���p�e��`h�۩���Y�y�0
ULlPp�{�5��=	�Oc�>��ӫ/�Ǖe���&w?Q��sgז��<�����{�ϙq�E��ew˕�Zk�!����(Ơ���4OI�n�ٳ��<����N�fe[
�s��q�2 ��w<�d��������}*����	�����Z!�LH&�e��c�>�0.?Вe*�b�u��h[��k�Q�$F4��L��"��C����z>@Y9�E���p�W���'��s���힐.�\$�~|�*3DP�U���"�I��`���w�0�лG��-!{`���~����J���Ȗ��.��&��x�"��
;����B�X�TɁ�$E�����Y��D�C�{��I��h^�ۏ�(��˹�ˬn�E��L#s�]�M�D ����N��MZ�9R��Z�5�ā�u�׏w&�q��-z�?�Y�����!��Wl�|��AFd�q@=6�O��'�Q*y.�h��%�����<�����třafZ��ck����2-$��h����<L.�e��skύ
��T��`k��_�,�xY�>Mm$�v�:	�p�5����W�x���sD�z\��L�����/[���)�Ga���P�87�)y�����Ck��n5�⫼)�v�놐�����g�D��9���e>'<����eef��:)��QV�.����+��2eE5�Zd�0%���&!MJ6�c��is�6����{f��?R��U/g��ɿ�KAf�p�	����e�?$����q���%�q�T�TYmY�a���ԏJ����v�'r@ԁ�{Yo�
��w_����,����]5R�@;�x��k*��p25�g���T~��'A{.O�z��tt�'�y��+�@�ہ8%R�oQ�&'���XT���߇�Q��V��a�c�_<�e(Iq�O	���1��:�0[�w����\��G�0�hN�u�)�`��b%�������?g$T?�v��(��7U:��ⱗ�$�4|�u�s���́�K(��
�nK�?�>^�FUK�y�0�0�;-�A)�}�s���%ߥ�R��8�����Oa�m�C����HA����ϧJ �c,�<��A�+��DJ���*��Q胻�+]t
��|p��
L��$ӌf��/��*8��%��A�8�eW�yWz��ɭ�i�Cu��C�VG�!&�;~�}�%ޘ�Z���r��ː���N�w��jr:6V�fY*�#_?�������-���}�K�O&��d�d(�;e��QR��ԏ0�Ÿ��x��}���Ey�I{�������Gq�V�=Ou�ҥX��v�ee�W��q}��Jy�=��dP]�W��:����;T��Y��hט�
�7�8>��C�EHї1P��mZ�(6_ϣ�ǈh8�X�J��V��`�Ξ L���R���ȭ�����V �H��ܟ�a�|��竈E49�{1`�������z�"��l���1�ڤ卦`�5���iE�>�!ᒉ~��R���^I�B�2	n򻦟_t�����/�D�v��@��l� r�H�r��x�l'�Jz���|<�yNo��M�OTj�f{#k���5�-rQ�7�}RK�˵ɀø��$bLMڐ�~���7�'���ңב�@��aT��΀S	 �X�֗���aU/�U��H�B`��؅V$bq�+
��{�%��r+���`����_�[K���<o���99-���]�[<�g�w6�ܩ����r �����,�'&C�q�P��=��e�5�ޤ�C�a��G�-��WCg�̍���FP����i�wD��{��XmM����7��l�;@�ֶ3`s.Y�O��ls�|��jm��p;�f ��S�?+'�?��gls���o�j��b�qls�6>�s��<�N�����~�
�#�:��̖U�=Ka����B$.++��r�?	�
�WVT��*#�n�a�^z���ρ�`�Ht���z����$ً������f
�S�Uo
�Ԃ�u}�N�����K[��'��9� X_��{:�Ap'��vf�/��I_d�]�m�/���35�&��Ԍp��G0����\eTti���/ϯ->��_��+�w�0�@�0U���\��[��
ޯ�󆣭ڜ�}�ĤE�7/VӲ�8 ��x�m�E<�\a�j����S!3��W4�?�=t�((�E6�F8�ȴ� ��X�2��s�뾏9�x�Zo_�Ö�e�lD~Q%���	��A	����=kf�T��om
q�X�b���p�:;�5%��|Kc_�ѫs�3B�H��L��:������;����}n�]�$���t�ӝ�� :��b��ey:pd�k_��cj���)]~�j�>..��Z	�2�C�>I��
�QOs[��a��" `8XQ{�T-)>�2-�h�Qm(c��Kgj5�Y԰�=d� ��e~���< Y?7��38GC������J.)߭s�%�lO.�lyڊ��|O2]$њQ��$����n��y𠽲��}��DCƏq3xI�RH֔�J̫�����q�U�rZ�]�p��v9`�������i!��XD˙XR��7m/#���}օ��ba�{�g���o%(m>����%�a�瑊��2ƙ���룕X�u��0_w���>�p�|k��ְc{Wޠ�b[y
����G��W}=��)YfL���D����3�.���	���}ӛd%��D ��y��f�{���%���G�Z���E8�D�<��%�N����5׆Yo�mL��������^z��v�*G��	�N+�m'�E\�C���)�t#	 ��,�/+ؗ��%�5�{L]�0�����rIyw��#;jRե�<ƞZ.�\�8���b$5P ��N�`�����L�<�Tw#X��U��Rt��~��=L�$��0_vLTb�jW��{�K�s&��	�@q����7=�v�M�?�&���K{�O�.��=�<�\�QVwU 撅�u#'���Ψ��LY�7�P�&�I�SI��vT��lE������ֶVJ^;Rs�Uq`���)��-��9�����Y��.wm�4��k���O�Bذp�IB�zl����d��4h��#�w��l��	r� �:e2��̪l�G�fg�ү��i�g
�+����$�S�|���eʪ�|h�|P�2~��y@�~��C���#�??�v�MK@�e�(� �/��/'���*�
�;%�Mq
=�`(ȐL���(r:�3>�m��3\�N
�))!�|�s��d�m���Ą_�+2l<�
 �g 4�n8%����,�r�[�غMP��M�6�R���P�g�1�L�whp��[ס]~�����%��D�o�99V� ?��͂�N����"1��CNK����`����P/��s�sy~�̆���S
�<�S��MO�ڝ3uF��N�̬�%��9��4���ZF�kw�x.Cn�4S��"���s���e�� ��=���(G�OPO�\���S��7xn� �oϲlV$WL�����2��$�Ta���}Kߌ��s���ܘx)v��+j��,-}�4�"�L��$R���qvsM�~���1��fT�Â�v�h�}�`��������hHD��l��r7H��"o��t�mX��9�X�p��c�h4��Y2�F�[A:�nz���J����ѝ0���������V繚Ç�8�������Au���y(���9�u��Lv������΁a �0*���P�rA��)��9b��L!Y��>��/�ǍrMD��)ȗ�iCcG�Z�c� ����'?a������@2��/�?���)�#�Bڷ*��� 6�u���]����-E��&"�T�,�,���
�P�i�,:���Ȫ��A"RV)e�T,�?��­����+^AK�?�����m�ø� �+(�I%Z�I�;��qZ��Υ��:�NUE̝mȡ�D��/�&�)P��Y��@��qό�]�F��4��_V�׈@D��b��%�F��Z�(Ր�
�>
.����k���=�0>i�^� MS��|�^@9��U�s�?��b�b����G
~]�P"�)�-����N�X��6oN^;ț�[�V�?��B����}��fX����/��XN��וw��h1���ķ�S���d�a��-�|1���T�unQP9<q�$W0�j���1�jI7�nƲ���8�(��� ��(F���I9�lٳj..8[0�@[p�/4��?]�����e����"#� VlK�7�������+T���P�W5��FY�M߃*At��%<7u��<�q�aG�ا�D$��x7��O�HVi���ǭ��5�J$�_�!��������o�#5������u##��DS��S��"�������3��ˀI�#�<&	N[��nN�V�*���u:�e�x�q��z�y��2����.1(�Dro�n�p?VN�8"^}�
�?t��eLK=�g�j���� U{�Դ�!Yn,y"gX�4ƄK�`��~s��a�B��H��VǴxB����kD<�gd���7�\���.�+�vrw�|P���;�`���}�GwGc���KQ�!3_j��}�����1q������ �����z�V��N*���p�ͳbA� �Y�Sx3$��1�~脣 ���8�&�&r���>��ʐ��t��O:�[������|����AF�������?��e
�f�E'�gCӠ#�/����e��Acʡ��smO\�ҥ��<�'G	�����a}@o�� 9����O%����-ַlɋ���������!�M�4+e��$V����U��\���}��^ ֏$�L�'��U2!�,�2e�2꺪
��V�Nwl�󒳫��3��Y�}�\��GC���u���k���a����4gl�?�D�u���d~�!J�F	�O{�:�8A���ჳ���n�ݑx��fVZ�@��9�Et��������( ʉG��_�Dy��2!,>nϰ�kBc���n���7V�;��-�L�X��������F��(1����S�8�&E��MeT����Ez�(�>���e2��
��
J�zA��a�!��c�<�n����M'4���3;f,B#5Su��=h6��reD����ޚ���Fj53� ��	]��_{^� K\��A(�D&�VZ�����8. d�xq�Z*���Шbe`�vE��m0�0��L=FՅ�Ìh��@t?�I�O���G@�%���m|���N����7�_Io���`��UD������R�+*�p�X%]"{rPd��"E��"&�	��%E�'Nc�*��>�e����!k����Zd��W��O_�돻�ZO4�ɻ��[(��ߚο�r����<� �^��r����ȡ���؇��������Q;��*Q�x��Вr�*��\(75F�X(��.��%\@|�lo��l����{���Yc�(O�$��1�E9 |B8�%>0C�pЂ�du���5�����i��ʮ̈́i�M��]����o�ZX!Q�Fݡ` �{|ǡ_�7c�Z�����#8R�o���<̄c������V\�@��1�-,��~R��X(��t�t�(C�~N�&Tbs|>���Cйq2�>+Q�����f���\�e9�i%���/�ݗg�̛�?��.�IR�J��v�D��>�J�/���*P�r��0�;}>V��S>�� /��LJ�Z&��6��S�h��G8�3B5��Ϧh���(e�e��TpS=�	Kg:�:x>[�2��+�E�xeҤ��-���Esk
�xE�|O�;P�=а6-�.(�����^�a�>�I���3��x����D�?�x���2��j��2����pqrª�/�g�C ��,�C�쑩iؘ�&`>��Bz��pt40�3��rb�x��pU��1��B%.Cg���_������n�yvu�sR�p_;v��lq#��#}�MC����i�Uͭ˵�"!����/N+|��8��=�m��R�״�������=������tV�ԑ0-�ý �g�ps�Sڙ|��dTxL����q�y|�����k�����v��J�K,X�,2/!͏*��Yπp�ߡ�J�7`�tu�"4[��va�"��ܶ�a��q�UL�!h���v ���d���c�WL����DZ� ���G��jy�VR�ݟ�5��S�'3�ۧEt�Е�����*0���� e�}��Gl��@&It�(��E�.��p�?g�4�
=Up�#ꢯ��c@N|��λ��~����.�1H�@��h�YJ���j��d:ݭ}j��(��P[����s������\���U�#���r�v�M�U�p`4"2�>y�j��9�9�������u��$U�,<ױzuUI�J>xpҋ%;�ee�h�H}ޕ�X���ukL����ޔ#}�c��^�ҩJ"����p(�շ�i ��#tϑ����ἦ5�TlFr2���3Y�Y�LWfQ�ʆsVat�`�U�!K��	�(�+��[��D���O�$�h��`�,��MR��c�E��|z�"��Ľ��{���z�x���g�� �zlk���c���Ϣ��W�y���8� 0���_>�T`�e+��d��-p�[�n$u����kEf)W�^������9a��0�#���f�P�H�'��a���$��h���:�v�=1�f�^��B�Q�:&�WZ ì�Q9���>x�_@�ZI�EdB/>�������C��bg\i��y��J�;���e�A�Y��-�2;H�`�őV�=g䌪�lyh 4Z��h(@�/�v,ų�@�5)�qt�%#��eb���8�յZ )� w�e*K�	����w�f���n�|Oغ����% �g�A�w]�b�p�L�Y�s>oy�!Kc�*\L��TJX�eMJ�~�#�R�����?���{��q\Ѵ�a� Ր!F�q����ёc�Sh��
x���@i�FDхK+��dw�"$��5j[�DI�=�Uv��D�#�R�����RY���b�y��᧎�[�v/�lO��4�����zAG��f�qm����z ��`�T�|1����%4��z^k��*G�O�fb��)��J�"���~�..���`�@��l��,�Xi
#�bz��.��u|��)ٽ��U��:@�|М��i)-�Z��)�$eee��:1w;z�vz[Q�ț�Hr�w��,J�-&���8M.oA�Zǂ��õދ�%���t4�&�=���g�������]&�KK4�{*v���-�i?È�}��h
����$H�^�&��[� ��p�5T���a�|�tҨ�'�i+_ݺ?f4��/���H�:$?�S_0P)L! �:�|ҜH�,�6��7_�8TuR���"��kN���, �r(�e4Qh�O`���Α��T�ȼզWF<�?Mj5uE;����b�����ɣ̺5(k`O���u4�)�=3	��_?S`wbh���â�I�_�Z8�f��u��MՉ�kD�Ng��R;�ْ�[�Z�3��7�J�3<ݗ�NWIn7-%�2c����r�������mzd�����b7\�<R�CN�h��}.�#5v0����K���y�G{��i1I�.�*��F� ��q[&�x�[�:�ClY�/ϒ.81ܿ^lؓ��!�X��QCiu�]�eCᛋ���n���5q�4�y��J^k��weKq�՘ڼ?�)𝻫�f��`�:)���ٸ(��ohV �/�}��Ǽ�ހ ��|�8*T3�u�8����G�֜��;��|����`��Ƒ�l���n��P�i�f�/İ� �LI��i������\������	F!��q��N�������9Ueʯ� Ҽ�鎑�(�ݻ>��&DW�U��B}�IE���}n�R{� ����F��)�<�紙{-�� �$/5����؞������9�p��Zs��ǫN��
�Dl���ꠌ7a5��9P�2��r�B�BF=1r�\>s��KuJl����x@Qo�kFG-�c�m����$n%V\��J#0�/(�?���C���"�(kfD���u�)���~�����B��yH��yX��I&!���X�!�:$۔w�-rv���;veS�f���RK�F	�T���S�n�d�H�}1h[p���n�����NB'@��l�I�\�{�I�%1=�v�xܨșy2�*�y�$u@y]�Xm-Z)wQ���< ��;�h z�a�@�GŔ���3+�&'�F%��wX$P�;K僓@�DA���< ����T�&i΄s�����n�KfX��K�-a�P������Z�^�;��#�)DFSP����e`�Wn��2�p��\��%MY�2��	K��J��9G?�= y��"T�7җ��O�|R�R��~���]|~@Z����QbBϋ��ܘ�g�%f�ɑ��e(\��4/>�/jÞNI�+��Buw�K��l��2sZ4)'�7i${�ɪ��;�
$,��t����球#��Hǩ��Ƶ�>kO L0�L��&�K�p�E%��lX�
 *Q��8H0m6�T.|4��"��R��PrKvh��������Ë��1�{;:���f&�I��P��OQ���8V�еm�Q�7�{^��5��-�}�\ �Y�P`�F���
E<����#K>�0ݙ��M�N�s�j�w����ks�"�XvMn���"GLu�D- {}	pN��?�@Y.:'vP��i>�V L�̪$�V�UQ��s����&���~֗SwӜ�,�Y�R���j��[�R�Jnf���H4c���1�>{3�Q���.xd�W��B(�%�X{���Q�:/͊���c��U�Ͷ[B��n�)%����WN�����2��!I�T�r�����:�{�*��Hh�C���7�
dk��K�Ip����/�H$�im�x��MO8���~�h#UT��x�<��w�����)����T������
k�G��=�6KD���z�R��������gw�ݽg�
�!Eq�j�D2���j¼7P����|/x h[�Igxk}/1��V��F����3w^c�w{^R�B������QD��;��4����F��o��� ��9$�l����;�ArtR�<����Z-H����w���)X��]�;6u�Fl@���0���P\	V���B5���:�sZ��x��:�4_��2��C�د���v�{*\�X���~��EZ��@����Ώe�h�טj��ІvU�)y�_��㩿-�����G^7�����R$��A
��*��^��*����m�m���فjwh%�_�+F���l��o�������4��V�k;��9|i;R��ca��U4S#�֌N���l�b�I��(�{&�jI��綾����ܔ |��A)^nM��M f�a#4t�u=���� �-�Z_��ë��}q�eʩ��D����$r��+�
ti�e���$�P�F+WC�*Ɨ�&8��P�b�.��%Xh��G�7��$�z�sW�,�e_	,e����6̛[������g\�G�d�B�V�u[�}��"(S�8끼��Ɏ}���E$���7?��H
e���5�B\Ƴ9��P'��^ju{�z[��>[W�3"z@������t"|~� ���U0�9Sm�<I�\q"��6���ֆ�s�?�D�ذ�4S�b��2�EE��[vxǦ����-i��t_�AT�;"e��Er�������yW~��#�U}�9��Ed�ܵ>�_��A+���HV����uV:S�
q��l)1(�	|
	a���;������ާ�M�D�=R��I�5����
�\�F/�7�^�^ͬذ��߀�m�;yɟ�?����>.� ��lß��t#�VB �����xϡ>w�B�B�=��SR�i���@V(���6���N-|a7���y�<�{5U[�WF�;�H]���3@}�i>���c�=�A����c`G� "B�"�ކ���Y|���Řr9XŪ��2�E��>m��{���)�죜���^	�빰�$r93,T�\W�[��K��i�[a:/eы�źǺN�D���6@���%K���A��F=��
������_E��dxBT�����q}�M����5Q��'Y��>�����4�l��l�����'��M
�>/t@��i���C��ZE��:��e~��9�s�����J��V"3}Ў��"Yfŋ�+w_4���V�ֹ��]�Lm����h�'��\H���U�}�.峔'�9��1�1��4ĩQ\f�#Å)3��j�R���>�L�S�c5�G��$y3��Z]�7�m,q���`BZ�,�b��'� qaN[��6M!�£�����h���!��=i]�ڼ�,�(���okji����Ԡ��<gPf�V�x����(T�Z�?e�-����k�H�(�Ȇ�Y�z�'<�orǾR.�����ra�x����Ӗ�q�L�Cyt�r�HʴB�͏���S���-�J��ma�`��K��	� eU�L���b}ZJa�6J�#�ɗ$�-�M�[���e�r~�NQg���ɱmCt���+��Y���_Cx\�����Q� �<�?<G��E=v�:��W�b�i���}-�B=}�/i��4F���U)��`���dS�5�O]w�U�6�MJ��1�P{1�=&�h!-v�j?�!)[1��3r�1��\i(~��%�9[=7���P�p�>��,�^�fV��(B���Y�������p����p�p삗�~�.b����.P��$�A�V�(�<m�C1��ۿ�{"���Q+����W��4�E1��G ��I�4av��Ig/,:��Q�9���ӫw����gҖJ�Q���C��c��MT��k�=�����&�@�thL(;u�*����o��r��z���~^4�%7��i�jrS�z!y�=$�H�<�/����c�M�G����}��x]n�1�3�ʽ$��g�� ��W�(u��,�9Fҕ)�Ei�ͺ�3��Ҏ��U��a�t�I)�sk�αQ2SG���,�EB�+�6~���Oi8$kc�%�i��/Kp���0>	Ѵ���a���Н���P�1�2�&��'X�����<x���B�H�	���n��?�ni����~��Cڬt��PZ�����p<��A��;�X�2�@W�<]p�^��9����&z� c�A�O�D����5��ׅ{p}�Bsp�I��n�Ց��N��8��4RO(˸��렟p�>�1����7�Ȩ��IhaԱ�|��&��/���*�Tm8����-[� <a�?�L���*�"1�[������}+����c�	��8��H�h�W��D&'ţ:�y��]0E'�?J������ԯ$�j٤� ?�;ci�q��V)�v4nЀ�!�:q�S�NG"�9����^K,���{�8�@�H���Q�+r�l1�c�l�7�H���3,�N	��8o��G>o����9}χ^i^�D�sl�g��{�?ޯ��������sb�^�*��ޟ�~���0ΫT��Y�����	P*�ƌ�/P�b8�����k��my_4`d�:��B�q�M9��&�%@;���3-W��?�x��s��Q�y��[]+S݋�/,�n�G
��B_�f7���J��э;���.��zLN�P ����
:?!{]�����'Z6�/�_����k�.�%�MQ`��p�-F���$n����f K!Y�gsW2�����{/�H~�=mAL�D��в����9�k��S���s:�T;��"�9K����(��1&13^&hh.���:�H��D�΅s��<�N<X�f�7�I{j�Yl6`6�h��x��۱��.rU4��uY��f��x��@[���>��U�nB�}g*����-����HA��V��X�+&D#1�`�^��R$�B��Q��́�7h�m�8X2z��[G��˃��1�!�2m��������%�BN��ŖҘ������c|[�
'f��!��FМK���MĢ��.߃U]��y��u����k���	3P� ���g;�z���oط��º�t�oՏ���3ģ�o����vn��q��z�@Y����43�����DE�^����?��O���V��#`_g�Q�7�+x*�(�����7��i�����f�<Y*Q�GXH �c�(�(�1�d�$�I,>���'ֿ~�]�Ȳ�p)�� �v���po��$(� z�CV���*\ADRe?Q7�d��;����k���m����)s��0͎�l��Q"V^B�?y��R�%�=	�\Q�K��f
_~B����RQ;c��x���+�O:P�n� j�Y�y ����}e�8��h��p������Y�Cq9Y�Gn�%SU�|M�h�ƹ��x���J[)��X�֠#�}�0	7l�ٖl���<8�c�)���")<�[1��n��܆��&�e��<�CM����nD�<Y�͓�7$jZA��J߇0/���!����@NF��9Hy�}l>Q�d���Zm�% ������G���������PD9�k謷��9��y�q��W��T�T6�V���M���3����%+��!��A��D��	1:�nc�NcW9�e�4f�T��/���2���l�^a���?FDZ$0����K�G��'}�ЅTb`�_�if-�K�^�P����K����g��\�B}bs;��F���B��ѩV�]�6�/�w2��ZamTy��%|���0��2�?]E?N��:-$Z�%́�!���u��yΎ�@����JG��@#�(�_?�"��/�i������-$�h��O�.�G���7dm��1\ߨ|ʻ�5� �/�R"��#�z�e9څ�!�6��2��P;�X���x��&�s�m���CCeto�֮�(��:m��u�f��پ�܄�n�b۸� ҳ�c�5q�w��*�/s�L��bQ�W�c�%�h:�� ��	|��˴@ra�4�h�CX9�[�(M�a��P8�<�H�c�$y��o�+���Ⱦ��˝�R�HEx��j_7�k�1�)� ��L�L�g1dAa=qx�?ZB����~S/�Lߢ硡�����NF�gb�=�g6��Q+[���o|ոkJ��Լ�{,��]���H1�O���:nB6g�!zG����
�4��~@��҅.���� �G�L�����d::U�߹(U����'I�6�7Iࠖ"�F)Y�xL=%#c�ٵ����X`u�I�eP���2Q2#�&�E�R���f��B��b��� tHIA�_���td���w�+-O�Ѻw�G�����e�c�9X��M@}���hhcl����y���OB$'i�>�	��� �������'�`=��L����.g]��U��Ӯ0�o�S�@�'XR��1��t��}Ϙ-O�J��)��KI��d���#����g^M�d���y_3g�M+I�ȳ����?[���}����� {}#�������0��~sUV\+�1�0�\oj�W3�)1_#g@��~�lJ"�7b�+|1�R&�K��<���4��
.abRG:�7�ݸ�~�Nʉ�ѐ�+�v�y�,eЧ�M h,J^/��1��]��������O�5�*(�+��j�� -W�43]��%�y�|h'�s��8��4b��~o�����1�}���Gu���E �^Wu���p�2q4lX�MO�8�w�J�����G�gzY�ќ5T]���	������|���8#;�L���v��
����6�O�sx�=��U��և�4�9(3�p�6BHm֡(�����줿w�h�$� ���{���e�dwo5C�pr@���F�Z����M(�9�Xvg�֍��O���.��"ͳ�K�	��Z��Y�����O�qD�w�)��)����:�(�$?E+K�����q���])��;�1��'[�ns�/oL�6.��(��x��j2�����ϙ�tv�k�|������w#R�Ҽ��,2�2o���A4�K����ܻ��JK�
X	�U���~A��E��j�܌��@d���&O8�:�e��iǁڟ@���͚�/����jX�.Nzp^�Y�����u�5l%��	�ׅk��D��k����]]Z�{���7]hmb���Q���t���x"A܌S�QD��ֵx��� LK�Àpf�%w��XlM�88��嚐�Z�O�Ye���T�m�P���/�M�^!�V������t� ���2L��bO_�(
��(�|>�2[��:[�/(��ɹnvt���"P��BA�����_�J���l�c�r������l�0aFm#h�|O���'�-��z��t^�˱OT��&ȅ��|�����G�$��@D�?�������K��rcP'<3<.MC�
8�Ya��$�|Pp0��N
!'�hڇ�j��9��)��rj�C���0�����'��R�Չ*��7y'6Vӊ�!����|i��bѴ޺�?)5x>�g=�0V����(əG�U[a��|�����&a4�%ہ�{�Yy|�s�}��w�C�^�$%�Rl9�rC�$o��E٭��pEݵj/.:�U�ۭcӀ��|K��&��0%B��SjI�}`�@��J�Tym���J�-�E�P%蘪��L:�ـ�2�n�|�R��q4��ϯ��P�%�����lN����b����k���ڢ���c1ǟ8�Al��|4.�K�;1�B���&rW�2��@�j$�uW����F��l;dޕW�LQ��pYh�(jgXƩ�7�1�����?�����8<�/�����x�ХYߞ�=�����i���NK[�^��0Y��?^�v��R}��x�"�&T�FMIU�Z���t�F��5�k#$~��w�j�O�F�>Ψ�,��t���蛟�69��$`7v���5�j��\�9ΫG�W*�΢{�	1h/ �I7u2K�)5�5Js�����r�ƹ����=��H�i�J'IW�ěP3�r��NO�n,�K�)a7tzt�H��`u�>1!]M�4}�/�L�dt�I��� �D�J�E�zp��i�)��R��� �V؅ɤ!ާT[��Uȸ�ᬹq�i
��H˱5ŋ�<���l=%3:�����Kl~x��P�_ԙ��P+�-�`&� [5R���i�f)D�r�Ǹj��
���͇�v������\F\��:ܔ�rz
�1��bO�Yy������Ն��"�"*�-ճ�$�E1p���^�K���(_�ą��F�$(&���"n�E��R��\�F��=٬$"mb���*so�xo�-�[��Q�k���<�v�[.|��l�N>����Ba>j�M~����B)�В(g���?+��M({%�4Jb9��wO��Ș��m{w���c4�gQ�_[w���"	i��!Ryl��&TO��NT�~���7��-
8I��J�#Q��}�Y�kـ2����f."�^����QxS^�Y���z�����D��)�Q�e$�=�z�o�˧�k?���Za�w�h<�Ў/�!����!W�!w^�S34�m��H�_kP�^���٥�Ǯ���yA�$��<+�Uj�C�~&ݶ��!�ł�?�"���&�y�r�����.�z&e���5��+������z�4�X�,ӓ���A�g�ʿ��P��6՝}�בO���S |�����3�C�讁���b 	�א����ڪ��r����?aNHk��f���5X���5�x'>�40��[N��ac�����@z��\o��\�ʐ���+��i1zT&3p� ̦8�����ɬ��_��uVX���a�n�O���[c���V'��~�%��q
g@
5������i2n��(%�A,u+��B� a�#���(��pQ��ўuP��>����oN*�c��x�Cw�\JB&zz����)S@���x#���ԍ� (���OL�ѰL����d��:�c�k{'Ѡ�#� �ßE�~�b8s����ݟ�� XR��:�$�Xuh�I�|_�5��>�b��0K��)����
ܪ��"G5А��f��.Cd��������A�����k��k��b��?/��upM�ܧ�vBѡ�R|����"(9�/��k���p!�2���U�qSW��H.U��PO����ԥ!�f�s�34�1�Ơ�5~$[Ϛ�"i<���q���7�Io�^ZE��8b*,&p���\Vt_�3�凓>��~r�
#�4�Amǐ+1��;��E�ॣ:C��2ОSf��uÞʄ��)��5JP����8�r�*�#�<������Y�+����ի��~M��2��P� �3oH��n���f�	�ʠi��q��hD���PpX�B�c���mV��sp��q��s�� �R��`�ȕc�)�:ͭኋ��T0|C�u�΃�qE�9⠧�r��� �z�Y��g��V�1ԛ�Nv(Nd�C:q�Mv�%O�y���=�nl�*G�Ǣ��^T� D��[�}�����EPo��|�z/��.�覌iШh��e�%d�'�=���������U�e�'̣���3C��9Y���ռ���E���2<�]��R�z����X񌋡v&��\]@�Tt]-��B�Ky/;BL�s�e���h
����k)B��?r(I2���-J����q�@�ł�(4���ڼlg�ů�P���ᰢI�"�)�z�g�*�첺��o��֨�{/��>lw���Z�����EA�A���W��4Jε�6�K�S�4�(z�:SF��������gmTigP׶��߮���
�M^���i �� YT�O �6r~S�����P��)��Ƭ�Q��P���Ns���s\|���v~�����La����6�d�YU�T�?M�=���Y@Br���?J��R�i?
���C��z�>���I_E���c�Q%9��}��\>�4X�R�^o��o��*I��P3!#�F?�?�ȡ;)�z�q%�v5�"LyΫ�XQ�/(|?^��5b���,�Tu�V�8�Ol���-#IS��<hu:?��68z[�p�C�������1��*L�R���ݟ9W�ɩ(��U��"�c%�U����R'R˽ɱ�b�돐aA$-�y�|��ua^��*�YK��~�z�I'��B���nߙ�q��;��*�$kߖp�����>v������fd�)����-�����iQ�ǔ8��|�2}:Av��ٱA%ڷ��wD��+��U���]��j�u���s����{U?(-�;6�2�p���
�����qz�v��(�gH,V�E��D9-��/�.��&	ȇfјc|E����� �h�L�U����m��m����Ӈ �=Y���L�����Q��!�j��@+Sj^\�!���
b�J�	�,c|s���^[�bh������ˣaۍ�)����%t��8���1r�(��e�(ΪO�ysJ��I[g�Q� 0r�7�"�LR-|�#{����r&�.S&�mD/e�X�� ����ĥw�m�F	s�����N��EiQg{}�����>�i��d;�I>F�FYM�R W�0�p0�N�/�y�ktM�����6��k,|�Qmq�ӂ�;f�`=u�B�'' ���y�h}�gJ �z̓a��7(��b�c��@/#9�0�dh�p��j��d�����]+t���; Y�>�|�S�Y�ڝk.��m8�ޅ�U�&�LA�)�U�[��x���[:_�T�՝PJK�mm�|Y�P���@�Td=�C���-~�R݊��v�#7>A��p�^$����� D�^�s�Uu�6?f+�~Ɗ~��C�[X�㋈!x��A�Fz��,��p1`�.B��y��*�
��gt��)����uMD��8<�;����H��U}���j:h�(�̉�5Ͼ.�w�`���]_�UC���O����e鵼b��I��U ��ٚ��c�y�Nr6����C�3�d�r�0�.��}�ӽ��y�Y���5�M��{_Ij��l���n7��b/yΡ���v�֊���X��0�m�V��񏯒zt/F��:��˻�����]YK![�^Ǹ
\`�i~�+�9�������9̈́�S?����N��*ئ�W
�8��l�@`�F��7�����^ʘ v��q ہ_���R;�bx�%c!����%�P�abV�������r���ɀ�ه.
���슏���y<�(u��V�B�������P��_4u���S�q�L����9�9��[����y�5�+(k�O^R��^d8��5����G
r��\�tJ何���,�1��K��M���z,q�_΂#���&��a����0���e\��?�q�=��� �{fp_S�.�"�E��j�F���SF�������!|�l���d/����)glH�N��T*��P0;�4�+
s�-��<�2�/�I����Ԡ�,X�w$v��"�T��o}��\Cy)?��ɂ����
s�t�\9'��2���p)ãvr"N�����~�y�Z.I˦tj��[�')w����=�K�+�� 3{�|�����}������2���Y��i�L��h������s(�"==�
g(V���ԙ?��b�n�|L��W.����?�Khr,�PzZ�^7�J&��7\)�8�4ke�����~�nҢ��^���C	%�)z!��b�?�䌅t'�ZuB5ʾ-�J(+х��r�)��A��ҽ?>Sc>�3���N7�a��KU�6� �n�J䶎>�F�$�1�W5NX��w��Ϛ�C�>����$��R�?�"�����u��Z_(#Z�:�E���\�=�M��Hb�qk��Y�=  ��x����p����)#��o>1o�%B�n랝��K��"���Tt��"�',��ѹC#.\
���f�k�9���I�Cz�����A35ﲋ�>��8Y,)J�!a�ޏf�M3�O=�6��&d�\Kt=~Hc��P�~qʿ�ʞ�B�E����	ϐ�c�| �G��S��~����E���k���'�����X���bq@��?N`g�a ?�D�7bLU��]�����z������)нް]��t���?��\
�+�]`�Ƈ��2
�Bp��x~�(�$���d�;=���߸����T���̦^�/&���d���
Ef��Q#�xSId��R7�?"ȃCW3�~�v����E�-ARu2IRvҼ�a�����m/�3�O��7�\���~�Ko"Ó̫����=8��,.2K���� bJM�X��x��!z_z0�7*�+�ɨ�ǅ�Z��<��F-2S#��@9�@O��fB�+A�
XH?��EG�Ny׋j'�8�\೬`-�	>ǫ ��Z�
�.��EI���A�.�F�O4�ג��$��w�,�Tw�҅~���Ӻ���'��z<����`ʆ�9�ywp[��o�)����D��p4�חH��Z4� Y?|*�d�ٸ5��V,��<����.}ȟ��1N�w�m�
յ�Q�͆�7~���>P(��?�yP% A��������qP���Zr�!t�}k�5%�Q̺y��w[7Z��:��.ُ[~Qp);㶎Z����Zs���Pi �`�X���b4�6X:��c�1-d�(��f�f�E�nim�����βә�ڧZ��61�q��E����O�j癷8��6T5
�0�D�w����XP�`��<ZW�H�������y~�Qy����@	�Z�zt_l���F@�&v�@���sD�S?�)�e�R�]R[�=��ddvJ����F^���^��/���N��_�pi+
`�s:�9M"]�ʔWJV��)x��FYLġ�Q'Y�8$D���o�J��>�	��W����]�M �?yg)1&�r}&��j�7X:�Z7�3��g5b��pQ�Y��_}��Kݪ����3�6�ґ��W��;w��n�0�b	)ʦJ��=���(po�aJUc:���VÞr�ƥr	_>�����p׋U�k�_�s���S�Om����q�}��zKl.�W����ũ����W�9_0V�
t�u�Nؔ1_�>U��`yN�S�'ե��P-F�.�:S˻�N��e�ོ�Ʀ��������U�_�JY���M
�*(X�cX �Y�B�	�+	#7���/������	Z�' Y����L0&�{����%���^�gG��M9Q���tк!�\��oZ�dl�z���zK.q*�c�7��S��2@dԸ���X�����I�r�<!�c�5��,U7����vS�Nu̪�<	Ũp��{�E5֟�V���d\C�p�d�οtۨN��8��[l��R������r�X�!{��aoQ��m��İ���=6�����}:��6��,��-�1g���q�4ץú-u3��r��-�Z(��C|pQ�:':͞��4�a�?Nh?��צڣB�o��M5O
�cW^ǧH����Mc�X���Aj�kvD_��T!�Sq�㑹����RM�i���f��ڼ�ߜX�͞`�|��ħq0�pK� d�J�����9��۶G���n����� C<����y3����x(. 6�bH�����g�3&ޯ{nk���`�6oKW�m
M,���:�<����~�`��@�=�o1����ٵ�`��L5�����	Iy`����G����6��|�oT�I�	�P��S�����a��X�N?���3��;x�H)�Y�� 2�w�/B�����Aq؞����|L�0:I���h�1Q���w�����6󔌂H߶�#?�������.��g���-�>o{�m;:\|U�m�K�e�K�y�:�$���F>��)R����	;��3 N(���8B�2���8�-=�zQPH�C�M��0C@��`�A��Q���G��!`���������\��L���.l�D�I��Ȕ��3�+F������Vq���S��zᎾVy�E���[A�4������p�\���\%_Y��Llnvg�����0 m������(:vf7�IoXƔ�E�������$t7%-�7H,H$P7��b�)��D��#���ˣEe9�Ҍ1�ַ%��\cB��{m���Pj�>�kd��]����6U$Y�R��7�%��(j�S��y�C�(0��]H��0����N����j����!��~Y��u;�\z����w��D���B���]P70+����2�K�d#�v�l�!�c tT�9U��N������� ��X��?ʒ�b�s������_S�Ի>a�t���?�kfS�j���X�C�A-dM&�͑�7�#z4�$vѨH����zls>T�x]����&��|G�nfn�>�D�f�w�,p/��,��"���������X?���6i>�Ĉ���b/��՟�)��5:0F�a��*ynn]]d�D��(��`E{���;�N�H�7@V�Y��y�d�V��禣`�5�[Ę,��:-��&W�.�9 ].B��6	��n۬�~�j��K�7뗥��Q�'�W���owք����=�������ӉJ�'�W���}�~w��\�3n%ﳀv���k�>�CS�@\)/M}��%<W�8��Ԯ� ��eQ����S�J��#��9�bv��CW��������u�<�ƅ6g����q5�ۋ�K?�߇�X.��GܤTx�
����,��Ԗ�'��
�A�G���;Z�H:еD�SAPH�j������RP����"�_S|��R�t����v�MR�u�cT�x-�Qsw��<v�-�yu)q�8|&%SX	N����=B�-�ƇJ���ww]%�P�2�gq�%-|@^�}5�8�ug��2��v��k�A�|��j|.���+����?�EuQ�;�miIQ���*�c��"����j��?[z0�{���ڍ�ł{G���r:Ţ��J�:��/�,��\b̑@��ȶ�����*1��P$���W���j�?{&(^ރ��zy����+����'�>mȧ�V��U`�|�q>Ȇ��D�ah&�(�PH����`��~|�9>���N�Xx�NT�]���^0S�p)��;Ha������B)���}��+�s�Y�,|}-<O�B�����kY5������rD���B���.�x�%7�J�:��)wi�B�B,��{���gNj#����τ���ۦI}���F����n�&�q�8�iCG��ŻW�l���,*+�75���Uq�;0�D*�nװa�x�P�N�ږ��G1�����d-T]
��·�y�\�_��_%�s>0��i��%A'.���B'�ř&՗+�i>h����\�1²M{�o�y� ^����t@������R4��p�D���v��r�gJW��'��9GssN\d"�M��~,lmڸEA$��n���.��0(ס��}�x'�����G#2�^���S��/��i��:�KN�/C�������bb!z伉�-����;ֽ_�J�J�lխi�}`�"O� ��W��Ep��{�\!����iCI`v��z̮Y��&4��nn���#jP��Z�1j���� `�m*)��U�ٻ�K^�+Щ�6�R�a���i��@ II?n4*�Y2mTpXz&ɑ�w8��,�=�vz����Q��0+�q����R��:�[:
���	�a��	�92��~t����J�