��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ���������K5��5�PɁ�� 4y�	����@/���NR�
�z�=�^����j@����0��0�ZR�W|SLK��UG|���G����
.���68=��C�eH��FmG^�%f��ϘIr𽯇=�'���J��r+����7Y�(�snS��u<l�/W�B���+���^!8�GK��Օ}�?[v����lF��$�4�w3�BD��ˋ��9��ʯc��QS6݆�E�M��#W�iIL�y�^9�,�#��^���	�0w������ ��.ׂ8������`��΅Q��s��[�[o֢�K�{�&u
�^1$�Q0G)��\�ȧ4��+�>�C�*d\�qU-�y)�e?���O�\�k�����B�Q�##UCG�;D�9}y[^��#��R,�t7SGj��xO���^�b�+W����i�P�׌ROʛV��
|��ϕ}�D����i�Э"V���޴���smvİ �ڔ?x*��H����X	i��)�h��4��1��1����L�8<[��i���O0�q<���1嘞Ǉ��/@o��lq6CE�8����H�%��}&g���
(�w��ЂV��cJ�p?�)�=;���������t�S��mQ0�m�wN�K�������?:x�#����A�ݸT`Z>����?�x�杰lIr	-�� �*:׈@$OT�R۴������	���D��Kg��N��3���d\�/(|Y��:�����9���Wmh���Qpy
��"Ɛ:/8��p�K�ɕ�l��ڃM�;�
2�&��SK��x[=��N�N��{Xy��:ݷ������йp�M2qg�ώ	rT�M=��	6��$=��U�6(�(��\;敡{860[F�	���㳹�GV
t3);[ղ���:�n��f����Z�}R���u��}�H�Y\��|j��i���Y��Y��8 �Z[鐰�����pi\G2D�"���0
I��,ˡ�?7x���-����RR�.���r�ʜγ߈u�(��L߫W�䤳���󵀝��l!z=�	�uLJ��V��ǀ�	�p���K��f�y�]68�(���ͅ�>ffϾ�^��OUp":�'/�ď˸��XJR�]h�}]9�
����4�`!�]��:'H���U��(��M��U!��&�NV�T�激��	C�k!m	)���U_�ٰ1q�}�D��'
Q&qA@����k��_��E�����o���*e14��H� (��V��i��d �� 	_���0W�� Y6;�J��52]�*:"V���O���j�W|�U����}�Ԝ���~��Az�*Y��ǧJ�U����:����*N�<��2�vƉ`�B�FW���"#6��c�� �K�~�%��E��97:HF&jo}]�[�j�6��5�Z�$,/���ٮl7%����f`���&v&Y���tb0@U�Zt�.��Bd� �Вl�$�����DD�B+j�FYX�:2�� g�e2�}w[�/�G����ŗ���=>�����V:,�ե�T.��p����\�N��a\n>d�2�Ƿ������&�_��_�<
P�Fa���T��S8��!��SO�(�y?��	��,���L�x�O�/�!����h�j�BKs��1�v�J_���Q��mg�+��0�89�����N@A~�(����������KS�)���k:i�y&l����72�S~���#�@�ꊄ�k9��a�d,��}�&��o��I5���a�:R�Ѕ�{�+�!���ɪ�dhZ�t�4���_���ֵ�4���K�s��⿖:�V#���8�q�^���+Ydݣ���Ī7���E��'����Nz�w����3+��/��`�pu,�W��/�f3{H����-N�J� \�y܅տU��Q>�3@��:@��:�'����V��s�\y�C���^-�ܼ"@���I4�4ޢM@)�l���~i�_��f�`\'�]�oh��5};\0��^i�%���Q�;'�xo�GU�U��@X
���@��L~�q.6�����U�FX1��t�l{���l���Qg�5�$i��A��W��l.Ҕ%*�)dB@5Z��l�g"|c���Zڲ��e.`�T F��~F�DERA��� "�zn�6?`�֩S&�`,[���Cl5x IE��Fr�h��u��=Y��C6]�KqӬv]��x�.�M\�JC@Y��6�����_�=�=$�a_�F��S���q��h�pQ�{]X�5>&l\��Q\u�F=�_����QhS�^%�QuLq�Z�ŰS��)��p ��,�1L�B?P�����E�����l�U������(V���Ur@Ӓ��E�������Oč��$�LԲ�hkE�C��u"J��\K�3	� ~@���{Yv���i�ˤ��C�!�YnT�D
|�x�Zh�A�(���e+-�6�u��=Jn�ujY�4�[� q8����v�r���8 b�6ebq+`4u�9��y��h� � #|6��2��q� R�Y6�"?��R���:�xRס��Ȗ���4	[�Ԉ��:���T�o0��ԕ=RZ ���\.,�L��ң�U��Ai�ӷ����:���)�Z�z�|4y~�=:8�\,O�ɯ�9H���[���i�v�X���Jf愝��_�>�+S����F��� ���z��h�e�lq�|׵��}K��ӅR��_�I�8��O9�2�(Yu��s"Q�x�o{,����Iý;��~�ii*��m�G<*~��o��Ww$���_�Q����<�C���5�pkIkfwʘ�,*���<9
���k�O�e]���3Ȕ�	�W�������h���G�*ۙ������������D�r���[�R1I�y��9��B�Jn��Y��$<�*Us���3ؒU-�:�ڗ�g](����*��S��qR.Æm�5�y�9�[T��O�6��4�_�rb����_����,&f��w���)������t>R8�J�}������Bf����sE��sf
7 ]-�v�%2�(�A�d� ��%��>5Ό����t͓9ĩ��yH�W;[Bm�ܷ*�4Q��AàE0�#=�)���u!���d��� ��G$
�9IO}��kdO�:�����ҏ�a�n�Q���1��vC �ΑHY��F�b�z�"�Y��A�Ĥ4�K�A�L3A��wz���T� �J6�֬�� ��&Idz܌W���8�"�#�;^��}�pvc�� v=��{w�b��?����{�I���|<�� y:v1ħ��˜N1K�3���s��PQȢ�ڬ�'P�$������=��d�"#_Z���W��3ro|�:~��\<kMk�%;̇�'�o�j��-i����}���v�i��ݟ��O޵�9����y6X��оk�ɖ�2���c<���R 5
�l-�$�pV��4d�ܫ�H;tM�~О`�y��*�z��Mm�.���[���8w�C��I�P+x��V�$�����z��_qu;�7�a{�+1���ٝ6� ��=n�<�5��K�3�D�!�N�lK�Pܾ����;ĺ��˷U�
�V3�sy�ql���e���j�L$̀9�+�b�D�Tg)�w���·�}.�M>��+e�"����Y_�ծiG�w��}3������N��N�5���~6���"�����m�ǣ�z �,��$�\O�Ⱦ�%Sʣ`�`�D+�O�b���w.�2�3�է9ՙ����
EI�b$'HH;��*F\�i�<!%+��C��|���A׈�E���1uO`!��\����L�rp5)����^� ����r�`ظ� ��r��S����x�@:N?g����X�HrG�IVW?�s�[�������٠)�H��z��;A�W+����Ia�K�P_Vh�	=��}9}����*al-9\^��9��{&);F"?�֣wwMx�v�]B����;^��Uo'{X+�cǫ�1w����Z� �*��3�\�?"�ފ�/[�?����72�'�lo�'{�m�<�\�������|� ��O�>��f�g�:�XE�Ρ�{BfD2�i�sx�����,6У�λ� �#��������i�r�?�517�,\u�ۗ�eNT�Y�eP�!C��5����&���e�X8Yz�ր.K2�Z�����)�P++�:�=�P��v��"�Y$9�n� )_P�#�����pў` ��o}U
Lې(/GX���r�v$j��X9��-�?�oq'��%�@�%ISZ����Ĥ��Q�LiP-�8��/3��h�T��z���o�sO�=����1g���9���n�o��iK�,�6��ٓ���/:B\8^ ���P�]�0����7&�/vB��q4 ��NO���¡��kC 3�JWxE�X�<�zz�Ξ�@�̄����&����&�ˑ��ϼB>�:Y@�b�Q޽RtĶ��L)�"�~���W����$�m��ĝ��Ì�)'�`�G��`��*���Գ��3���o�ra�#;{�lsl_��y�#�|94����m.M����&��}�Q��[�m�냸��H�t�Q.��Y��wp٭,)�`����ɨ�s�"