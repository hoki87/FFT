��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#���������l��U�~�׏O����j9�PY���`T���x���s����uí������P��"��b%>�1eτy�<�gܰ�N�Y�	� {��I�ɍL�ݫ�G�R�k��Q�!E	�5E��.��:�͂2��y�m�-�.E��i�����YS�
��@�H�ۼ��nD��Y�l"BU�.TԊ�=�-�����q���Ǹ��j��ԋ����tr�a�ٵ�]�b	��%�ɔe�)rYOjX5;V��R�������M\�	D��ҏ����9c=�Vͼu��Ro�P�Jf�tRvsY��c�"n�XO��	3g���Q���^�Bʹ�7gQ+Г���$�-��t�8�����A���<����l-��*�|d�B
��"XCQ)D���1����qQ��b/�?���q�ЃyE2RE��9�v�4��ɕ?�d�O)��G9��h���}�X�!Q7d
����dEM�3�o'��#���Q���ce�&y�i��@��1/NH�W��"ʄe�������[���R%�}kha�vv�3N�{x��ɏ������,�����abpj�����q��ޮ�V�D�͏�<ǻ��%)�	b�^��-����/�n�Jc���Q�D}���9�4�)�y}X�7��Ѳk�A#NZ6qI���X�|Lz��3�;o-�}}�X��+HTه�?�ko����UfH`���
��r�&v���{��^?,���z�`�|<K��C�QZ�r7;yX���X^��J �kgv��'�G��[�51�#�ʽ��c�{c��<,���b�����hm������魘�G���lu���SM�ĭ�5ly���R��u���G�!�m��Cؤ�� ͰZ>��p�M����~@4e\��M�T��'���8ϖ�s��(0��`�!���rԭ�h�h�==(�1�_"y�i�G��կ��,7�M��K9���jYQ~�O���3�_CV(!nuf�U�";9��Yc<c�g2�,�z0�1z/]!#�����4�r��������{��mN=�<Iճ�	��	�;[�R���x�e��UVd�ѵ��Q3:n�ܩ�3>^�Z*��,�f���K�%���ޝ�u���v\�p����]�}IH�L�(���;'�V�ľ�P6_s;��m�W���>+�D�,v��g�>�R���%,%b,���r��|��pv�Y�H�u�����ʤjo�����I��R%@�X� l-_˜"b�(�q�I[Zpa�8�ݙ*���36�m�Xۺj�U��o�
��=Q�Zr���ٝѯ��|!� Ȫ9��&�c�+��nb�9�/A<l MZ��)��������Yt�4��3��M�{�-��O�l����;=69�>�q=�z�s�"��i��5#�s︝�zץҎUѤq	�<e�&p��m���%PK��c3m�6�_83m�u�G�_��Y)*3-�ҷ���R�����o�i��7t?J�+�7$5��7�Ȏ�k�>�
W���!΅��3�e��� %<��@����M�N�e\=�5k���=�V�V�0�j=}�8SGؾ�Ȫe��J�AD��u����_I�r����&=�oT����$�y��Y�q�&�����KRu��=9"d+Y`�|����b���7��͏�?9ݕ���]�p�)Bg6��C��ND��~Ruc�LR���QB�M��I|�sڣ���R���(�(��<u2�s@9��>�0]d�����=�#�6��Z	(|�����HJW����'ah���+�li�BP~B:�<��ލpÇ��[
џ��Lօ� V��!�Ǭ���s�'�l���`k%�",0�ҥ�z�s$SX���Q[�n�e��F�rI�_Fs�Ho��T�I��H裲���C��amm�_A"�CK��Ԍ�C���m2��n|$���E_jcdZ(�YҤ��2��N�:��t�Lc⅚;sn;��³H�S�������mD�%�dy���x�]#t ��4$ �l0>��<�T�����)ҪLѸeq�(�1v��7�o���d/�d�t����2Kp��� (�H��Ϸ���a�lQ�~�k��#c�H#/*~Z�PCd2��IK���*�����;�I����g?G����^����������$�`�q9�t�C[����x�y�ds;ϐD$� ��A��sQfW�9�x�9�F��!a�?-�| �ĸ��$لA��d7޶w��'�P2J�Rh��80H�*g�n�$
@c�u6�iT�.@���J�����0���in��0��-�ܝ�����r���l[�T�Q<h�lG���&~o��� ��?�����-Ţ�Ώ�P-��]��w��7l�� ݴG���Ǟr�j.���(t�T�vϏ�!]��By��SM�+	�,Z�˺oRI��uiB��'�@wp����d�o&@�(9�/�����y�|�JP�_����S$'+�#B4����7m�J�����Ec����p��n܉�15������?�j1� ���P�yKL�y�e��,��u��$5'M=7_]�!6�fؠ~���NXb�k�"��yl,s���D���/-�@fϸe�_�c|ͱ4�rpۚB�������춭�?�w�AcT'@�������*��7�hϾN ����~h]��+=H̗D�~�v���ئ����	)p�c�`�=��#�)ۋ���6�c�`�ۍ��<�Q@�^,ᮿ�6�|��P	���;k�:�P}Z�$�D �M+Qűq1��؊��(��&�����H:�m*A���"X��2�ϼ�M�#KU��Ĩ$T��6~�1��6l9(S��G����h��P>FO4��ڼ��0���_�F�\tq9�XPC'h#��.�_Ԯ2����u����������ǲ���F�R���kS�`�cү����%JS1�!���u�t�[��p����)�����\TF�� #;3�`�T5�� W����}:F9�z� �3�;�o��y|
d���?���n�~5��٬Q�·��������;Sh�}{4��3;OE����|N�+��R1��޽$�8��*ar�"D�Fu,X�9싖B�0Ҵ����h�QUu��#��+� _�c���_�zK���x��ş�'�� ��<��p8����P��m}�s�C0��J  �cbI�𻣂�3�dSν�b��d�r�٘X�A�GWp�������A_���Fz�e���������M�3�W�_ܹ'|M�!��O����-�����<�zE���%�Z�Ԅ:j�S�T2��Mc���p=�\#IŰ�Q�r�� ����7�%�Z��VOT�z#^Ѡ��1�=I8���X�Z����??����,9��� @���hi]�#^
L��N���H��i����?T��?�y�7}�Ŏ���:c2���[�#G�-Wf!L�x����,f�Y�0�Oi����h0.��y���P�ڸ�LNt7[ [%����@���G�/��譫l����!�}*n�������� �xs��n�v)(K�r��3���s?����{ո׽"y"�rR�%��25t��]1�-��)Ң�(%B�{Jlm�d�S39)D��fԒ]�x��� vm��|����tS{�Z�A��E�l�9�w���.�*R�T:��.(.��m����y(W�nK�f_��k�q_n�H�7�����2���S�M�I-\W��:��ϣ+ΐ�f)�@q�]Y\�ˮuSD�t����-9� ��]���D�p�b܏�]���!Oz�哸un��5|�1]eC]��ʚ�w3�n��բ�N�U��E{z���͕�d6��ěVop��Zn�Q\�Į-�]V��$��:�n�*���.���`�01W���+z�!vF�������b��@�������z�g��y���fxQ�N�3����:DeI(�c�ֶ���E�/�*55Y���=�:.:[����p���ڻU<�N|�����
2^�&��>��+hЋ�l�TЍ�"���-�"���&F<ib��-I,��v�kǅ�l\�g4x�im�xH~ �7L/`��d�V}iу�R51�VFD�Q/Bx<�4�:'�]�[3~�k��tŦ��@�����/���3�r�J�_���:?3�YU���{��>�鰾���R�ld��fM�o%9d��ڟ��	��\.�I'�y���d-J%�u�)H�ɯ��^�3�(ش/sW���N�����7h`�Y����������j���b���U"SA4I���yv#۟)Џ*W��B��#�m���z~t~0���S���sMl�,Cm[��
	m��m�U}�N!R4����\g���stk�&2�
Q�	�U���A�<Hx�.��<�,�4E�*��4�s���yG�~��U��k�����Jϸ�C:Ee�9��T}/c6��!	�����4!`�V�eeD�2���# �fE��#�.]��O��l�o�A���=���ܻ��|#
3 �/j��i��ߜ�Z�:M�-�����<(������W���~qO��$rtN�x��q*�����d�J2xK�C�C�vj��qV�0ЭH�k��|�-T�f��Vt���>�~�Ѳ?��NK�(?�o�Ӻ{?8$�Afx��'b���c���1�-�%�=��P���Cx�I���ZN?OZ��NB{��M$!�ط�<���S����q����O�'�Y3ؗ��y#�����9jO�Uv��|j�>��a�����sLW�x�y���UC�H�Xا�y�Y9��Zlٺ�M�G�'B`2�w�����-EIϩD_ĉdٕy`����z&	�ת���ֹ� eg@q5ʬ�3��o�4��ܶ�W�3�U��#H�iR���LQ�|0?N���H��nu,��]$z�ľ�%B�[y��p9�+,�egB\��7r�V<�7����_ٞ5nQ��T�2X_~NF����gz�&W�b�m�6�p��9����[Z:�r������hrB��>�>*@7�
ھɆ<�(�����@h�!�:*N<[.ړp�֏Bd��U��EXyj��YXr�z2�WΥ�2�(�7:?�C]�!.� �t�fLa���U�F�Qy۬G]V�����ԋ���6O�K��HЋG����b�P,yS��9��-C;*�
�A�Kصi�o��]�C�NB\��2�E��H�K��dN�<x�ٌ攐��av#��=�0��ݕ���dr��rw;K:FtL`m��9h��R -uR���_E�z��O�K�XxI���g��4Y畕{-B/�nv�ڹs�:@�ꤶg���'��=<��T���۩i��o8BHcht�#�w��?����j�Q��W_x�gwU�N��3�Kͫ� \�����$��֯4z-ۢ���NFl�*xW@�*�A!|�ᑧ��K�VsY顋�9�ɶ��ν_�5X膄kN��N#�5�3��@��<Q|UY!�WO�l��������%k�������/πѕ�9#i_�;7�|�zqD!��D��9!����1زI=�(�-�cp�AC���}������t��_��������Y+0�M��t9Ӵ�����i����qh�Ly/):+��X��W�ԙEL	=�����'=���/��e`�õ���F��,�/I��j��O�MKl��>�O���sGV>�ERf+����Ցwp$�Z�b�x�y���xw�@&�N��+qA4�6���"h^{{]�,��v�� ����
!=���A)X,��R/,@�}"�-E��d��AP�9���J�	a��Ǆ쌆�;��)pG6T�C��ţ_����Ѧ�n7���U���v@t�a9��S�*�бh#ҏ��.|\�0��������7lneݸ��4���<�C���gG���J ��&��U�H4^���+&n2hy�01&b���@�k����7od9A�a�y�;)�q8����~�B�ӆL-�U����;϶)�����<�I��}��䄜)�v������R�td�?�+4Q����z�=3���>m>%�i�<{̂5�F�m��x�2S�����5��R֨������#�"�.(7� �(D�
����0'�ʜ�W�ϲ��P���[�/��.�R5q��ht�*��B�3Q�}
xb���U¡�ś?�`��P��|_��"~�Xod $6Hlb�x��87|n���&�_^bh�uXo�ܐ��=�ٜ|m��d�
c ^�*^6&BD��f2�f�a�j�U�n�\Eݺ©�j ]3u�Ҩց)	���T~P����y�h9*t� ��Q7���3fu��Ю����T�h8��V�_�6�돰�T�g�����/���4���%��Zd��qU�g��q�޵8�(�F�ڑ����Aڹ�o�~��wDy��"�ذ� ^9��v�t�H{�?�nʮ
k�z���e3���rU_�HW�^?�u�\��B��NGb�Y�d�Q���|ˏ�N�k0B�I�xZ�Φ�9MC�I��}&}��}s�hϙ 5z}�|cMVy�Q��z|RD`Q:�6�/\�arH�m���~�JX�aRqz�Ɉٴ�%���d����+��:��x��=��/g��]f{a]S��i���V~���@;�0�)	�־�Q���I0'6Z�����~0
<��I?)�ĝf��j�9x6��t�Bou��3��V<�~}%�*�gN	J1Ƶz��<D.����+��|�e�\�	���e
Dԫ-t�d�_W�Ͱ@���D�͵4����Ч���WS������yG�g��$�_4���ڴ�);v�o<�>�˞�>�W�|3m|s^���E����_��LyN�2�a��O�}{G��:1,�^��.� ����r�}9<�zd�{�3�or����w����j�
j���w=��!9k�2a9+�O?>)tq�w_PT	��L��8w��S"$3RÍ���O�<�+��'�3�D�)އ ��Ґʍ��.�fiG��RR*��nC8���:j(����b����_��1I���3��<3�����6�3��:�A�.���fJ]7�����Q��d�ؽ�Q��%�Ty�@d�m��q��in揕k��DW�ԊaI>�����Ӆ��V�_�6k��eŽ�0o���Gm���+�<<&2���F���z�ǧ��35�'�${���~�|���	ux��Z0i�m\�0Z�VGlY��=T�k�bs��j?�������m�I|�|��\�:d�e�v;��ƴCs#94����:A�3Ǫ���G��r_Ɇ��(+�5���A���Y68rl&�F�y�Q�󬠘��W"��O�bX���i�$Y2p�̦~33)�Y��9z���r �������F5cF�yn�_��ם�C�4�CՂ��qL�@��
�˳n3�B8��y�խ��^����y��O;09(�h�]�� f����Y!�~���Ќ`Q��'�~7U�@���׊]���vG�q��~�-GNޫ3[������x��P�;�^'�Y��׍܉���RI^�D~Ǌ���{��XLVx�n�_�+�LZ��A��ǔ?,D��! ��RJ��	w�p�H�o\����C���<u_��I9���'�u�.����K�����a%��'��H����&�v���ɠ�ܲ�S���n-ѭ�ʦR����k�0	j����� �[R��\�2�qka}�8R��N�1��F_XH�uU�͡��ܜe�b��2�vT�t���Z��x�]F��I�t������..1\6?x�P�ߕ �P!)e���'��,[8�U�QN�J_�Zh�y&&B5|�/V��o8�c�6�D�.?�S1���w-���߈9Y���r�e�zY���vs|�M/>�������^�X���Y\ $�;6��'��cp�^\3z�|)�^����)D�E9�iܤ��G*�!��W�MI�i`$J?L�Y Ʋ�C�Gr�
��P$X r_ebn�ڙsA��Z���Po��7#D����f,!�����O�e� ֩6�1�����)�H;���ͺ�Z�`��&���- h-�*��N����u�%s5%3Jp������u3�	[�&�h8A	�+`�q��{ڵ<�������&��x�-�e�U>��^�v_	��?��x��EX;:�&,��($�OML�����&������PI���* �Ȥ�^���&�K=n��E�^�����A,z��v!�y�e\��~��N���w*=N]���m��H��cK������,�)��aۻ����� �e}%���Sf���`��!1��3��7Ѥ7�ݙ��:�L�Xf� �}�(�?�#�Xb/|jq��q���FwÙ���;)��#`�(�x7mUH��ҭB�
���_�I!|K�h�����Kܵ����>�*���	j1�ͯ�E�b�8�3��S�_/�?����:�J�;�Hcv��<h��L�]JF��@��r���)��fI���/2�^a:��p��� w���+xZ�7���#Z�w"�N�H�U;��ad����;���y� ���ڡ�d�m�YR��~t�h�k�s�����p��Rw��\@��;�<�>V�_�;E��ȹ�����-��e�x�����ycH�Yo�dBCS"��U������#" ��3��n�_��w�(.�2�mm�+.Y����U<P�$ݝS����E��i\F�!`u���L��u�W���Gl׸�,�;�ł�=�����)�C]���-�W���[WV��A�@[� ��"A���3�=�@�L(�D��s�vU������n=W
�u��*,�8"�m�������V��ܬGP���m����D`�8�`��0(�����z�>j��M����N�b)|"��GQ1��Q=��$w>sC��ݱ��������+���Y޾S�l������` p����(�z�M]l}{�|{�������F��Z���Pe�O@N��oΫ7B���ȶ�<E�E���Y���Mv��!�M�7q�Bu
!��m#"U32k#��#�:�0�����k$���qhN	�c����"m��!V�B	��r$�$Td.`m�@.��=�����Ll��ߘc��@y[�aB��~�U�E2E%�0�w(�eJ"��n`���i�uK�E�<�o�v5`PcC�����C�� Ӓ�j��J�����T�3LF�Q�xl����K��l�/���'g�I�Ԕd`$�!`u��R7A���C]�$��>H"|%�<%jM�-Y+%�[�#��J�e�W`Q�UT@�I����2�����	vX�Sb���Ut*o߫����u�oo��T7�|r[�)n��Ae��؎CV��#n�9�1����L�ֵ��sd2��('Ҕ%��Z����+�1�axV�;���l��IvK�Re{O2�s7����ޢ�@�b��{ۮ|�D6�6b��Ql��K��%�xrW#��s=5X���y��g;S�CVS�R��bV]$�wȶ�,�z����H~nŤ��'�"s�F�a��L�)U��!��$�#|+e5)�űnF�����P۝Uu�-ɷV8��c���w����hG#�
�3+[Hv��	%�Qk���`K:�����*P�X˹5��s�`9��t{�W�ԡ��^D�`pTQJ�ҧ� ���;GT.�#"Y7�=���N"zZ�{�Ϻ$��&�����w�:9��3����gJ+`�����	m�f��if~�K|�7宒�������MBtd�xT�TvL�F�2���;;��U��hC��}����!�b�=w����>�Ap�F�R$۽PMف��_��X�<D�{d8�g�d�z�"��A�QkB�B�$���D�'R���3%|m��uI�~�oD�J��b����m!�E�)=bFK�mӵO�
���H�1�h��6_��<y�������1��Z��髋���%I�|m�&�F@`+���kJ���Jb"���N���ǰ�06P�� �T��҆Mx�K�N]V�+�p\�f�� ���P�bߏ9��T/=Nt1G:����I����b��$�f��aP���	5�o�gAŏRm��Ԭ߼�b��{�d�w��%�vL7kN�m"�؈���+:)i��J_��4a��-�X���]��|5��Ռ�R��������L{�&Hp���ᘃL������0�u��d\ќ�w^��V���$�\�`�z�k�ᵟ0>RDh�E#����S�<��)��6��^�:W�g�(�H�E�m�;d���Գ��s��ݥ�>�&j�46�:3G��>�
i��'Y���~m��.�[�3OJx���搬K���A �ֽXA؍��3.BH\#[��i�@�.�:c�o
'�Ke �/l`/�&Xp ����{׬]P��(H�<�/��ȥs�Pa���)�ڿo�;̰��fqZ~��@F"߁<����R2�-B�3	�����^�к�:'��%S����d�[O�g���$7��1%�º���k?����-DD��$������q��ݠK��6�`P����9��U�D^��z8�Qo���GU��}Zy���t��d�No8'�Z�74�k���n��,��sH���ti�[¹�����F|j�����D�4��vg�o��9  �\%Hy��7���@�i��R��G=���h��C�`�g��Y���|+}�X~#�^��:�����|�0���3*A!���9P��D�H�=&�����te�D��"譖� +�u�V�3����S�nϱ��ۈ�p��R$ňrgG��h����4���W��)�����H��u���'q����א�LibLP1���C���0@�RK���ɔ[�Z"�LȩL�0���V?�^�iONE�,6cM`j�`UPQ#$tKO�S쩷���>�W7��1�`T�#��c��1M*�ybz�z]���������T���#SJ�M�����d����LZ��qK|�ɸ��v��cФ��^�ֲ�3��8�$�B��真��>��g�d_q�y�`v�SXeE&���ʎ�@���]w�bEǛ#�%���z�tVok�B�'��p���SMJS%����!ml_ˆ��6[+k�^����X�;
�)C�Og9yb�����q���L*zp �A+�&E��"�K��<��z�tO:�1��c� �6d=�I2y
y��?Ƹ�������Y��������JSm*X��_��uGTHA}����~��F0�Dz�f���<�N���Fنv�ы������Z�vi��M��Q�hֻ����18�焉�S_�ĝ�cǔ́<.K����T"=m���8l%p���A�k�Ҝ�~����ߐ4�d�*_$T\������3Q65��5iji�)L�R���09
z����~�ԬM���D��,�kwxo���2�!R'/DAC���\k�j���#���,���,Q}ɇ�8E!S�Jx��!@j�c�
�\�%��g��Dd��m�ۯX>���ooK]�t8�7v`���]\����a�����ww�Z8��^�d �0���]�O>$�+[<��<d�>9�!��|̹j\����h���D�,c�9+6K�Oz��Ae���!��P�>l�˛\K)�"��_J�N]����"1���'�F~J�2�w~@yH,�wS=Y ���b|&VT���A��8�<�va)D�J�B2
7ix��OX�s��V��x��dT9$�����v�*��ii�I�SՀ��H���a	�q-�Wl�W����C�+��0�'�5��JkB������O�Bes��WJۣ�Q�� ˚���\ߺ�e>�0Z�dt[�2�[�/	�[����E=�S�Uz�cԾ�ON���`�mW�o���w��,�����D��߹w�k��>��'Q)��0��o��s�$��c�ug�ʻ�a�:m#�b��{�#'��a0��R�p�{ �O�*�̛ i����1�IuřA�1,Q���6�{���V���q]��g�]����o��~/�L���`_̦/\�Ѷ Ou�ώ��0Q�~�B�C�ʼ<��2i����E0��ൿE̺�勺�$�\�CJ��,�~�k�zd��
g��4IÞ3R�=�b���;��b�!6�9��M'�����mg:>��ݤX��;�}��N�B h�(5D�=�g����U���@������>&�1(!4��v ?a��a�3��B�q�#�Ǖ�|���Efƹ��|�^)N(�+朵���R�kF+65�R��=����;���i0k��J.,w��?(����ԓ-Z���At���_����/n��;����@6�T�	bi@�S	��$b� ��o�f��J#`J���^�R
��7�	�q'N4̆�i��UZN�G�ܱ�x�Xk��m,kݼ}*_����3nY���GHi�ּ֭��
�BZ����La��Np����C]H��ݸ��	|���hm��;C|� -� 7oOȔ�)��5�POEX�3
Puk�{��Y<|gEgnS�j��Bz��X���"�F�o��\P�)�X����&��S+�@r��|��U zX�ۏ�r��-"o�if%l@�}�dZ��9[qU���.��ǉ*

��//�@r{@=�d����k�����g�p'�iL<�k��0B���n�L�;���eR��FQ.��Yf��mY�������ϾpK$Ųy��i}U��:��r��/V{�����5YG�����捑�%A�C�ꞇ�Ȃ��6jS;��{w�����6���p�~)��ޖF,������yM��!�e�1�9�G��Fg�uH{7���/\�jg
7L��I*$kU���a�����lA�'������9���yP)�U���uf�m�؃�7Ou��qd��}x��EJTKL�f�i~�qc8�07��r��c���^6Wf �<+XQ,y)����������@"8�spQ�qL1�uj�I	M��l=m"="��W�K����k�lX���u���>#y�>�?�#ތO��:G��i�W��4d�\�*ʙ	+�	�,�˪�p��F���~J亁�Z�]�	T�֎8FsX���zka��@���$�H䄵�I_�J1J�yla�Ǚ�l*A��s8�t�#�-��|�P�~$��V�U���?o�Z#�.�%$͕M��4��f���Tڂ/�{b��O��0
8m*8��`3tb�H"V�����)LWq4~�ե7�H�!��x‿���5�eȇQ Y�(Mw���(J�/L�G�Ε�L��4Oc��-���u��p;�����`9��ǴO����<f7�S�Vk.��w�{�[�Xڮ�2Z�N�2�>��?2���ѫ#Dr��٬kTV��U���=�#�Nw:�!!�;F�}e	J��8�u�=�L��1?���1�V�b�2o�����d�tG���6�ll~%��#���k�����!�6�v8$r;��������Sr���P������{� 6s���۰�[���;�X��1ӱ=���o�毯.|�� �K)�!�	�ֿ`��)��8��Zo�*�_�hp��y�δ���D����!��ӝ�yR���U�[�7dZ6��ӭ�D� �5��s�0�ΐ0�u��7��^��ӿ�a�����922Z���k�Ī�Oް$���?80k�����q��8��_��� �&���/ZQ��R��ќ��M��g���#�5$��R�.�W@��?p�cޣf��6��pnU�Չ�\��|���w*�J;I'�Na��߽nþ�X(L�c�j|>��y;�!}R4�ż*48\z|�����m/���x�����y�U�ldC�����َM��<;m�#�W�
��G ]�nNV��1��ȡǮ�����*x�pVt8M�Ń�8�/6#<�<oz(^��I)�������7�!tΰ��-�Y��
F-i�:H4���$R��l����� m��Sf'�R�����w+����(��W�;�u��h�>_;��=Uպ{kc����}�,�H�S[�w6婬�<��}�:J��9�=z���4v���m��@�P��[Y���Q�sJ��'�y�.��z���SӇ�����rM̰��\?�eM�T�QE�$ё������Գ@�'ĉ�?��A��R��Gv�=�p����E��JD��M*�=��;��)ao_ZE�rF�����?V�	���Ʃ7k����IPd���ܟA����e�d
efo�a�bE���Q$��C}���.����/�.~��°�:Ϫ`4s[&;<�-�BQryt�h�׿�:"�\�Ǎ:��Z6�] Q�j��P�����	����:p}�<=^��t����fŔe!����_�[ +��DW���7�x���?{/Z��n��q��2��v���5���j�A�͈(��i�͢\u�h�mTJ��J�s�y�J^�!�D�,#P<;]���,�>���b�B����͑�c����Iv�V2�������nl�����^�`j����]��Ȓ0:��M�f�f�]�Z7T9_���/���u�D��|,�\k�LiX�R�x�TN!z,�7
��*�D��k@K��0X�,�]]O��w�[1e<�4[�qr��
ҧ��%�wU���D���WX��vt,ٺdD�r�w�Y��^��ėY�VDkI��;�W��g"1�{��z8���u:k;Ayg����Y��&VH�gm"h5q��;7�Q�{�ȅHܙ���H�XL���� 3������ڟ�=?�v�.��M����vily
N����|�/�	*KԮ���X��,���Ps�ŭ�¢�@d� �	)����\�l��~g��6uz~Ea� 3a�����BZ�r���^ߩكFV�}
��B��C�?��^ZB�=�|㙦&���r�[>sG�7�=�y�W�0j�nm:�����{?}��[�,���[�~��7uD�ɴK�x���6����e�6�2J}�X����j8�� ��?�V@!� ��཮?2u�(��Ågd�Gn�7��o8Շ`�BN~2Ƈ�3U�7j�뮳T/d������~Ah�6�5���'�rе�s��*>7�W��U�^�5�c�JԨOl��!���WҲr��$����xE��8ĥ��"㩈x##��� L��p/�=	�
uKҲ|��YC '�K��M׹�T�<�f��k�t�j�+�ۡ+{}��Hl��6+���3n��ق��q#��~�Uǀ3m��_�t#:a�[����b|V���vh���aD��<�@dg*�����?<��+�1��PiW-)���_�U3.�Y��烙����\�	MkV�ۀ{hK�rU勇J���@'�Q���52P�S* �����/"؄)%����V{EٌV����I_�4(������_�=�&P��x��<#�i�TZۘ�X|��ɽn��$��m����������imK5��Ο�ιH^5�,��g��R���dm�Ǚp���dθ1Ȃ�a�HD�v� l��&,�a��J��׈�!c�AOM9���L-���S�a)���S��C�p�?��Ø����SC���J������1X�� ���Lh�9Oz9����՜���f~��~�"3�g�p3P���T�
w��#9���qd�V%$p6�fW����1��cd�i҈�'�䏞Tү���csW*:�r/����f�����
�N����謾�AV�$�{��$�	�U�DY�u�|
�-��J�0r�3�9l]G=?���!T�S�f�����R�t#��n�2	��c�[�(C.m��ge�Q�O}���V�<>��������E��h#+�{?W�so*�7�ܢ���eCțS*ԑ��<��s5lGa�# ���n�
����J�}��㞋·��.|+�օ<���K�zVY�k����a��\��Ys���ğo ���=��-�����j���H�*�;y�r�H\P	�UT�3N�ᛜ�J+b3�D���+T��#(��맼�5E)��d��u�]��{�OF���oF?�>Ϻ�KS*���t��7-�x�w�����	>�s��\�Ԭ��Fּ��M��F����8��,9JJ�
�
���wb��˷ٸ�y:�}\��9�L$��7��"3w|5��$�w7Y�$�@��._�"�3lum���}�YNq�(�+ڵ�N5�09�KVb�C�cs�:6���� ���\j@-Сڞ� '����?.[�fY��Nt	S.�޸! ���Y&n�P�k��G-١�#c]r����7��:�����@Z���wt��n��~u�l[G�sM��Ov�'����k�&T(ų��ՊI���/�d�'s��:�ξ�V�q��L!B���{��ImB�o.���P�]y34X�%����Zn���)X���q�o��B�����Bk����;
;m��4�~X��;�=���"���j&0�O�Fn����(�ǘ1�LD��;�uuJ^f��X������]�ȓTf�kd�V5�E��vJo?lȱi�G.���5��f�)8������>�A�H|�r͞�)������CGF!�ޓ.�<��������ͻ:c�o�1)�@��ް4ˋM�@�����V��t,��̧0�W��3ݕ#a�|��2�o�6M#�g�K��*#�
+��S�xx�, ��S�t6d~�'�k�d/9�9�ŅΩX�{��ԭ@���`�iU�T��
�X�|C$�d*��[��W>����-.����C��Bа�.,F�_�AU+���=@K��:��{E\���T��IY�/\b���{�u�pp�Du��b%UQ������4J'j���)�8�:�i�xX��@�ػǞ�K�5�B�
xH`�u�rc�*���p��w�3�Hx|C�������t�=mH8���(���k8�G͵��W9p��{���M)�Xn0wt���7`���|�/Ϻ���M6�D�t�s��S��>L�\M�ָ�C_-^���~�z8�'6�C����EKxc����L����At��I�)�Y.1����*�p9��d��^Vxf���}�M3��7l��0T���S�Z~����L�^���2�Rԁ9�hP�x.�������M�^F��X����{yD���j���B:9��"�]���t6H":1��o��^n�H>f�$K��(���:,"�`"(����*N��%�JGGie\�P�G<��o��/���uUB�×ĺ�!o��w��[0.y���Ԧ�{9�K�p&�� H�QAC�JDX�
�!�=t�4.�#���%��]�Δ(�tFh���/��9D�������I�Qzp���y���d�C��Yp^+>��9�D�K�
�i��~�N@UJ��;_��*%ߠY�7p�C����`V��n}ũDt�9����W�o��'EĠKtE?NJm��}�!,�o<�_�]��:MS���
y�D��Y��$�"��'�؂�ma3���V�%y����d�&�4�~���z�4��l"7r�7����0$�sYu}+����@��bV��F�K�ci<�s���#��9�{`9s���t������������8�؝O�e��?�Ydi>J��+�����JB�N�EZ���G�~�{�����C�9|z���a��9������C���,6�
,��1���2>��!��0����3���08V���q����-�-���(|�^�A��=4Qh��g�D쇩3~�/rug��T��̎�ZQ\��A��W0d�'���x���jW'*-1ן�;��b3S�G7H�~����������,����h��(�jܞ�|��T���Rd����/�&�S�q��g��h{�4?�8�-��O�{�N*߹O�/Rikqϼ�&�5N�`�F@��+�|�&ENb6�`�Z�J�)���o^\�ى^i���^�ʬH�P/?S��_�'[��0���2��i*�tn�g�mK8�W�2|�5أ�����ᚘYӔ  p��yZ�Zaln}�C 5�F~$mR���m+������;�������:?��9j8�e��Bk��%���gn�|sܕn;�C�8�됸w����TX��l�s����?)���g�����wW���QP{yq�

�gj� �Kw�����w�|��8�Cg���K�'��΢�4���`BBԏ��q��Ϸ���hWC	�h�A��ف�d��O��Ċ
�"F=��u�]uâ��m���KX�V�y�9�2�#�~�?�f�"������P�X�|���|�_�1�����b�Q��1�$��}��Ie>�v�h.-��q/Sr�ֽ��-2���4�^]�?�w���fD��%�\gr�O�e� ��%��El8l�龞�}���g�����e_]�b}� $b�.r^]����뙫hJ�z�(�H�D�>���R!o��(���!�,�`�ځ�o'���g惋w/ޭ%)�M��ɩn���ތ4C�uAɓ�١fl���/ΩwN��;{�´�2��&�� ܏egu�?�1?�qy���i{'��t�p<�����3�jR�$٬D�K��V.j��Rb3N-rя(�ջ��Cj}���'�ԫ���i��*�^S.?�*�>m���d&	HD��0�ٸ�Z`��0�w��/�Q5�9�f�S&(�g,z��Z���08̵}y�(sa�"5���C��*����=�c�>������-��3��w��	u�~( �mo�Ta�OA�M�3�!#q0�P+�C��7}_��?�V�T�R��g&M���Hh%	�`Ҋ5�%.iS���Ra���L�LJ����$����-ք�E�Rl��TS�o��BHC��4��G� L��2k�F�'�$.��;<�̟3{н����p�9MxW²/io@���5��F��'�������^~NhpyoE9����������������MeO�NK�If-nދ��'��$�y ��F9��0e��d7��UfW/��ۑg��Q�5`͸4�m�i�Q�n�M�:ת��A�JU'a](<����>���O5����s�x 5ӡ]�D1"�[�)�*���߇�pS$��W���Fy����:Ph[��5����35/Xy��B��#)��� �!�)�xa}+P|I*o�����m�|�˘H�K[������ ��.o���&J*�>%�TqԀ�p��$��	C�>:�f�4�*�ޕPs��٣����A�Tj��L(����3*R#���M3�}���
҄������>���*��ư��Ͼ��ZV��.�7�g`)�HP�T���ba|��|E�6͟�@���ơ_5�ST��O��N�l���t�>uP��*&��+�#P�&��C?UBN����l9g�XC��2Q���5�=��0�#�1P(8ְU�0>�<��a�gno_c/���Hp�3��: �9�g�'y�i�
�M浘ؔ��!|�B��Fym��[��Gz���d��h����n}��(��evV���W�y�LLf�QUv{Շrh7�b�dB��S��� 
��]��%%-����T]Hi'	�}�]!͒%2r���ͭL�,ꕆU�3�����J<[��A��ޒ�f�W�����xo�"WWcfA=LW��0Y$9ad�<;��S��'Na�Q��[��1PD������՗�^K��0J�w�z�i��� ЃKk��؀����$�,m�b��Z��(Iy�\���٪`��0`H�B��B��7�X����:(����HI�D��3��2�<4Z�q���yw����Y�c��̎��DN��>g.>��i9����x'_���A�&d6�7�/��U退��@6q 6@Q�<!{��2��e��	��bN�v��e�����_�U��04�m"Ɔ��'$��XD���%�����8^�}�8,ʓH�2ٖ�F��3XƆS�n"!Z�.O�d� ���M���o�(���M�%��7�Ѡ��:c])��&��"%�3�QKh�(NF�R���X��_��v�*S�|x�U����cS�����"���F6�խ��X��U�D��;;����{y��>y�0uN*�pU��qF��{i>��g��	�p�&O,��������L}0�*��o�f&
\��٦�2&�\$	#���'	��<�硥�r(>dĢӉ��(�� ��������~I-�N6*�����9�y�����'�S��ω���{"]�KD����*����̙Y[:��K}]12��{g ��'�w<�`(�k��Y���Yo�)��x*�����'w��[�]��L�"b�U�7�6F=�7�1������BZNs}:�:h~s��b�98�|~��A��P����Jc;=8��:����!L��C���,��z�v{"�i�<-�W���'ƹ=� ���-6WߠXp�v��6��T�"Gs��f�*?c� ���4��
� �z�>�ԗZh�+ڭ�G^ig��2��MAAPA�W����|md��&  ��P�P����c��@�_D�m#%����h'�ûQj�)����Lp����� Yk���4!r�n|V�b���M�� `y��epg��⤉)�s)X���P\���)�|�*{��(���G{�¬���dŴm�`y��ܛ�ㅪ�b�
5����Q��Q�4n��Ҷ�5�69l�F$��m<I6��Mޡ0i[X�7��[&4r����L2���;Ke�խ�M8�M��2:̞u���MZ-�%��!o�,fx��3И� |"d�Â^�Y�p;�X��b��;����A��i�6���.P�4�3�vH��m�����@^̟
����*��|��O*� ��u�[JD@�_�u&�a�i�Y9:
d��m��P�DN�(�����j ]#kt�'JM�)���i��~�5	�ɵ鴊ӱ	�c����h�k�I��H_"I�4�e,8qKI���f7F��o���+`!���1��B&���K����b��u��A��[4Ss�{��v���n�=��[��/E���w�R���2Nq���x����\�ߧ�j�EP�]����*$�s4�%�X�� �B�`���<p7&�ǩţN�B��8M�&�"!Ȇä�:s\�u����[��H���ÅɃ(�oQ^b��v�|䫟�
��N��9&�T6�yK�Ƅ6�������9"c�c[)����1�9,�8�M��m7��%K�;���ug��&m�/�R�(�F�ii����ʕ�-���$�9�j<tx�e4F9���
�;��i��O;ty�s�+�gIz����2`��_Os���/��:��Tٟ-o__�>�ڞ��3�/��i�$�l��tyhA�ȭ`W"K#v�K��?�J +�y8����5���i ���&+�� C1�R��C�K]�+�UN�L�`s�Z��*�v^òު�E�'}��	5�I�4�L�\�2^���>�Ǣ�wK>�.��_p���B�"YC��	2��zC�LT��Ҳ�V'N��3�����{�a�����iS�P��9��̓@[�K��d�L�4@����|��^lPe��6#�h�z	�����v9��฼;m������E��~������[��.�g�zx�!��CO���5ql��ޥ�Cl#�~��"EZ@�G�0C���pU&�xŬe�2�T�ʰ`���w�h1������hO��%�':�gӊ������u������&��w ֣���'�1��=���<�Ao�?����,��IR_|f죯�{12����0�]3�o۪��攽��D��E��l�}�4���==d���Gd�T2N������=|!Ul)a��p͏I��S�3�c�w�9�qT��1K�eW�C�(�F�Lig���}�0�4��0��ޣMpy1Z>Y��SZ7�-t�ُ����9>J.��d[����X��բhF�fw�������&x�������p����t���#h�3F
��C'��h�g�)�Jؘ��yA�^Z�J��cVx(W�H����ҫ{�4m�k��Vpv]�᎝�~�����>�)DA�^ZV���sq�&�TQ0y�����9u�s�Ltŧx��CO��_�3���ڗO����s��=S�D�i�pq1�H|���Zm��OhS���h�O� �Kmݞ^���0�u~��]_���䩂�9@�.��+�i��Ja|�Yi7z��� V�sWp���>4����9oM��+XٳC�}��p�̂�f$��V|�h��	b�	�b�b���kLM��`�W��p;����X���?����箛�f,[u�[8�d����9+�+����E�m!��=`�
>0VtT��R݁�s
��v�Qc,�|�^�봩��������	�W�I
�6np���V��Q��.*pZVNy^mk�����Z�u�0�\��4b��+�t�-u�$1� &�M+;͖��@q�#��� �![���m�~8���0Y�e��3�]7o;�m�$<�n�����<.�o��#jm�R2���J�>82a�y�� ݬ��X�R���\Q� ��f��V|s��ԍ��>�i(�y��Qq��X��;�$vf��BC0hT�^������t�J��ݥ\`\�nbٳVz����N|Q�6���xh���F�<��C&��h�\6�r���HDߵ��IT?���!�yv�uZl�աn/���%��-�҇�ur�|�nx�5\�Y~[�ͧ��d�<,R���EmT:_󤃦Y։47cL�����y�F��
�weR�7}^�q�Tt��0v]x����A�v�F�-�TV�ֆ`��m�t���7-����%����$1�B�N0Z~�c"�5�����A�&�M��JD�����d���٬����XJ�l��#�4�ڗ%�i�IG�舝� Xk7�nx�ޠӲc�����Nc}��$T��#��#DFrS��n�v%ܺ�,'���A0p���� ��%�'C �0.�"YFXұ�eK�Gv�8��Tc��;��4���4*|���6}n�]eL�폳ѥf���W��.�q�	�Q�4P3c*]4\��7FX5��A�>��u'�B'Mpp4S�^b�G�趧0��FcY���Y|�w7���˱��դ�K�>�Q��@)���,?�_�"C/��"q���h֚-&��U�]�k#wx�$�_[1wL����m��҉�ڂK�Y���g�ړ���f_����F��1�m� <�M;��0��p3,r͋ �S�Wi,K�l[,R���d�s
����j���YU�'ٹK�4�h������=�1��|��W3����b�o|�Hu��؋��?�޸#�K2�R�ϒ�A�ru�!�>Pq��1WYN�&�ӌ0h&�U��t�y2[WZW~<�M�5R�=U�ʞ�ǳQ�ܶ�{�\xҺ1�,ϙ��o���lĽ�&���?��dH�CCF�p��,&�����@�7��@��̼v��r�\�ASt�s/~�>���	fn�g�d[�Ό����c=�s�i�|_�~���5�DW@G������P��cbV\�i�O-�P��ь� "
��F���^�ƛ�ЫP�����{�b<�m��� m5�&X]�f�Y^"AHM~{W!���EF$�A� {\(\�PUH�����9k���0����4#��,�Q�}��d�׋6�<@#ԩ��z�0p�	ʳ ��I&B��[!)��5=l�E3�����!`g
ބ�VUK���u�(i=B�w�c�W��㵰�sE=T���r�^��F')�ԫJ1��pc?�B.kPF�[\�ӫ���� ���k�v������q������"�V��y�Hž��RK���NǡN��j�'���j��R�!�cN_2ԣ�	��-�u!Ll�ɿ޺s�Z��'�اU�dT#Y�/�(9ߜC,3t�8n����ca�Ȁ�J��d��[����r�=H�Ki`�v���C���WK�-su�]�˻�N!S�֖U��˱�\�*��5��8��!�ǔ��`��QD̳�t��V=`�� ��Ϛ�q���:NU�^D*_���ٯ��:��ԐK��|��KHN�Un�_�Ĝ}��ecz�$%EQ�d� ���קg�,��I ����=� �v�C��?ZW�@�j�ob�5�7.>�o9�aw��^��:!a���zJJ�P�i�c��;��<J�܋;#I�Ig��b~�!�%R�f��6ÇboѢ\Ѡ�S���,�x�s3��W�6.O�������EL��͹+�5L��=f'��+}�N�����$ļh�r�$yul�]6� UXX�Uv 4kT��R����L��4����ٟ�rz1Nƍ¦
)H��w�h1�M���V��]�J�w�k��c��'&b�������n��iNh7�=��h����Ait�Gl��pF���KW.j��f_����Q�dc�7�{]�e$�-=���dL
-߲&n�ķe�8X�`[����.�v=���4�VR�t��nC�sU���Rm�G��̺�ߦB����4��f�E�ZAwrO��P^��D��9X��x�� g6�]hH��+��>d�Po���r���R����S��@��p�����^Ƅᳬ��԰n 'JKj�#(-�*U%��b�>��x����<�I�	i�́Q�B���8H9qn&4_�o�7�L����G�k�p�	sS,]b0���{�'���)��<(+��#���N�9��`_u��1��;U�SL�T�1���xeX��,#'co>7��w{9Y俭%���$ɄA����+�%	�/м�ǁ[��D5�&���@aӚJ�f:G��� x}���&I�T��)���̊H\�}C 7��J~$��d�c)���	�qZ���C;%�g��n٭QSKCzz�q��Ιǿ�wԡ'�\`b8��f+����WJ�����S�&��p2��L���0�hS͘`�d����J����1r���%}M�<l�^�ZM�����iK%���x�5�@�T�!��	H�K� c�^@��u֊^e
sfX��)�m����r���Qq����\zj�d1C��Z�����bR���Ϊk[�d�@͓8����)ZP�1�\9W��?=e(��Kw��#��H���L������1p�s���N�`���G���w�l/�(8��<c+�E/R��E���顀F#�Xl�_|�1�4.�LF�`�[�̟�lT������5�e/eD���������gA�l�Y&�ި��`#��3����]�&�B=f��a�M�D�x�u���)��n�__[�����;�S>g����b���+'&f���|�}�
nU̦s}܈_�Z]���lqOx���'�r��UO��r��- ��f]I-�	Q�,����V;�u:F�D�����Y�
���^&GT�/{��M���G�[l�4�mxE����7�R�It��-b�/�&& (X8����܉��v^�r�?��,��R-��a�+�A�%[��c��V���+����Yg�����#����t��s��P���-F��4�d�t��x����
�(r�;��0{;�ZR���X{�Z�����S�s��=�A#�!bBo��A�O�qz��!(��	��[�����gz��or��3�٥��f��Ii0��3r8�rL�_��f��dA���-�:
��l�YT��bux �x�Lt��*|w	r�����;d��\�A���We�N+aִ��=4����r�aΈ����YhЖ���x � ۢ�wVQ�(hO�Z몡�����X� 4���F�貴֫#��~1�����~�A�I� �ig��P y��#; kʃ�Ѹ^�V����>��Oڨ�DD��ܘv� ����0&�@� �Y�r����}��f���Z�M(�3�Fw���Zd��f����^�����`vR���ϲ�-&jJQ��1��z3g5#4�Q��㒿�b�\+N2U��!��P�U�}����9���ALl�G�&� #����[x�Q��qe���"�Cp���`.sI��q�lx$"��N�C�ŭ��G�����)n5t$i0�4	\�o�<�Z�>Y�����S���.,)�p�
T[�4�Q^f��`Fƾi�!�5�����A�(r�cr}b�(�Vj�� ^LA֦�L�3Q,��g81�_ߜ���Ǌ������c��/����!M��[�l��m ep6�������uo���CR8�!��������I�ۗ� 3Y���O,g
Xz$�{�����L��E��l4����̷�峾�]W���vMV`3`�VF�XǷ��Kw~��t}�ٰ�w�nf2P,�f��������X]!��!�=�Q �4�^��'���F����m�(&���{��2j�xBhN��'-?��Կ���,�̕r�(�Jqs� �Z'r�Db�5g�hG}� ]9�mxı��9�&��*ױ��#������6Ե@�%�&��i(b�P*̠s���ܯ~�2U��9��!n=rC�k�<GHqz�=R�Β�����M�a��1}�#�j�DU��@ﬥN��`P����S�@��j�8 iʡ��p_$�q������T��/��FuK��b&�?<vl��F�Ψ�i�3��x>�����(O�@�r�nڡt��
���F|��,���| �5)8���@u��L�ϭ7uSt�:�n�m-*�0�II����tɁ�2�핟;(�7�׊u
��Q���QE�e��5&�� �M8̒���Ǚ�ɪcg`��*O�xpJT���䆺��T&�-�A�ڣ��q�Prl��f���A���pS��Ehs�VG`n�!AQ���ĵX�-�
�%���V0QU�#�1>og�/�￢c�<}�$���Ul ��Ou	*�1\���	�F)�"c�f�s`��SE�K1C�={��L�5-���M'�T�9I�5w%��{��M�
&{Fk��)��-���\��AϿ&��k��
5o�x�xzW�Ө6ũ5�)��F����v?���SZE���]�"|P�:��s��v��P��kb�Z��Lh�*��s���I���H\�Z C�9��sJ�3@a襜m�)-J���O��@�Vf7$���Y��{�Y����V�|�xX7fkO$�yQ{9A��n�JZenA���s�gƚ���-o���e��^y�� �.>_ �rp<��g@��k��S��Z�4ak��9�Ye��
f}a����#�+8�،�#[��7�̡n��2�37�����!'�l�bd*k�vg��@��l��p�e���������	�V�%w��$�e5�Ex��e�p˰w(�Cd����k5U¸d1{�)�
��w��-`�4K�xF�m�������N5�S�#��D#`�!�R�f����!y`H�xq�n�Ч.�!g�{W��ˌ�h���1�sc�E[����9�ů]�VW$(f<≜^K���Y��?�������Ba���t��pi� l�^���jy�-c�Q*e�l?i����0����d��?�L�{��[R�8F8p3�<���q��}a	�V�7j7�Fj�B�2�XZB��J�\��'������q.d��&�ú\%��:��^,�&�0.e{[\�V����&�֠c��f��m$�B�Y���ԧ2W��w�+��=v��M~r���p�*w0}�jf��G��D�D���7��|�|5��aW�Ycx\��!��Ӄ���Q_�c"�ch	�z��Jh_';r wWo�}db�)-�=���dK/�.�{�Do7*��Q� ����_���;����=B�?":�N���W�2I�S-��"jhm�M6-��o�9�R�v.a���H:�E��L�ì
c�IE����PZ�&]!a'B"{����=���h�-��i�h��T0BUs�Zr���E�Fwa����}pX˴��(F��L�9r���k��(��	��}E=���Z7U�����gQc�	GVY�� G�.z���O�������0M��3CT�қ�S��R�?��Xnآ���2�)��D����Wi"�a���� ��i���7+�$�psP�2{�5d˱�X�П�s�>F]#�M��a�]į���*ߕ`6A��7�O.�a�ԖRgwK -�����K�
�?��u������_���d�^U�'M�6���8��2E��s�v/ٜ/qOQ��ʰ�3�Ңn�Hk��]Xđ�W��տ2"�5�sBh����1�R�'Q���1%b|#�\0��8%�MZ�<��o��d�Z�-��>������Fe�m4���4NG�դ��?`�@P9K���V4e�Ґ��"=
Z�8'|��H���p5R�H
0(��2��D�lr��-v����C�S00�MX&�����C��ZZ��O����M��f�V;f�7��͈+���8@
`+�,g�o�$`v��F�F'´vH���=@���Z*�Q`6��Λ=�^�ffދ|�P��T��W}O��]���"�?�hЉg�#�ܝ����c�qJ<�ZL*:����B��A�F/oٻf�X�t�b�E3����D�C����Z���~є�>纡� C�|+�q����v�}dbA_��΄����Y�մI[[�R,}�l�>(@÷~%��J���(�3!^z�8�9����*�4e�:���u]*��SgD@��r�,�h��{�r�t�eb[l9�Ì��	���e���ܺF	M�O3jB�¿�L��Q~�(���R�ՃN���){���u&RrF\&�輽���]��z�Ձ������=po����{�o!����F�l��G3�`��PJ��hz�f;��>���^y�G+�]	!��$����b�qLW %��� "|�:�1�]�#*,���E���ﶪ꬟F��<s^�w<�g�x�f/�)�Ƈ;�~�H7�eqS��ү�P*�>k�w7q�����x���1"�a�{`��,��=/#�[�g�M��%�P��` ��+A�zU�F�2�Wea��|��6䮆�$��0d"�Z�k��UB� �8���A�lM�/Kk{�B��e_�e�|݂�m�#UO�4�Bs�V��X�b���)	pڑX����A5E�0�7�<y��~���cAd: _
O}�:r!b��d�N?�N?vF�[�3��ك2��:�>���-�d�<*x����ؐ�҃WD���|�}�e����=[	�b�~�WEi0�^&b��1
z-t��
�H��{D��0��SZYK)�	�j+K8�>�5���ڸL9���>��u�9tC��+uX���ө7���ϖL��Ek�ڎ���dӺ���6f�R����곂�&[�V�V�T�h��:���x<g�sX�:��W��U����K-�h(q���2��_j�%�Sd*�^��G��( ~Џ�Q��Gm�e*���D����]]���9�-8'��gM�T�0��#��_7�>ٗ�-x�p���C�M���$Ǆ^�d*0h� �����Q�0��-�#ˆf�i����9��9��� ���F�˛e.r%9i�:e$��]���S�Us�8'�`���/6��kF���N����ԟNv����`T�������S&��lp�I?=��2�V�r\�:LXZ��V	_��S��Y�]�U�&�^��4;t��4�^����?�;�����%�d�;��'Ȇ*Ǧ���?�Ex�>ڒ�Z� F��۠vN��O?��u�i��R���̔�������qW.Di)��"L��M/�����辜Z����(�c��t��=�nS"�%H���x䝽����69U*��������~��
CG��%Y���/��ݓ�������k\	l��s+���V�U���Z �rX���<�R�/�I�hd"n��>��HL����6��+QQ	�!f��2����y�C�@7�n�Y:=�O�|.ٷ[Ec�t����N[x3ͥz_�j&*��9=�ǟݬ�B{?�� g�K|�z�4u�]/��L�}ib�o kH2����Wڟ'�9����3u���R�7��d�	�l��T�M=�1ك2h��W�딭�i�>
��?V�	����NY#��)�r��7���������M�I6z�Ψ��v$ ��<u|��
	�ٓm���d� bR��	���/"	��y�^�ʞ,��E�E�;�kd�e�S�Y8��|{շ��
ɖ��7u ��Y��U�ׇ��,�(q�j�ئŃ� �I�c��`z���a��1�*�C���� !��� 5_*6Jڒ<�ţ�F������5O�.2��o]�0��<lw/|����T��-���0ª�]v����T��8X���+̆ɽ����	.���,���0U��?$}��&����L���Bcp�wm���wg��j�ܪ�b����b�����ˊ�zg���a�	O�5وRګ��RQI�K�o>O�j�+7�z��afPK����ֶ�+��M�]VT����ʓ���G�c�8Y���f~�&����;үF����H҆=��jG�y�����!_��V��	����.NF���������@r��{��2�����3T�����^�ʻ����.���3����vf?����\�Z�z���� ��+0�Po\� 4nib���I��s�� ��Q N_�2�������Z ��d��+J��y5����j�znn�f�X����%�#�V���4������V8�����W������N�݋��|���a	�S��0�(*t���?P3��0a��5�C�b#�1�8$��QW���6���끁{�`��]��K
7�:�=�i'x��w��[v�>|	�7��ۥb��%ÖCj������f.���g�B����aqf���#������O�~�UZ�w	����lX��Ve���dF��J�Ud���K���
�������w4�Gbv,���b��u�vAW�y�L�owO�H�ifރ0TE���� ��z�Eߵ��T�/�
�'�h��q�cs���	�f<8g��Pt�������H	4uy�'�VUN"��>�t|.������WȦ�#`(:�/���d�q�R���ocUZ�)��,���a��sZS@Ms�휪�8��V��m�3q��1����j�N�MNf\){z�!�su(�m��[�߄*�Y�%UZ�)�N�~����<:.�M�U?%��!߭�Y�b9����$�K�
��8W��\}�"�3)��(�����6`lǦ[8Ψ��E� �MI+& h!zi)����X�x~���I��ŎbRa`Uy��i�
�瀛�����7��w��B�����yJ|GNZ�٣��=�eƊcE�4�҃`�g��R7���4���߹���=;Md�\3�Yc�a�c�y�2٩�E }��̻��T�)���6��Tv0���$�s�53�P��'�$>�ǯ�g�VWP5�*��jC�Ieq���	���<}֧}F��F�>��C`���~K�L�����T�+#v�̮G���vD��q!�>��d��I6��I�[����Oj#�۟�S@0�]�!�$C�Ǝ*xf�6V����{�$ߖ�O�a���9�ɥ�Y�rN�R��L%d�:���I�/�Jƍ���x��R�ג6�Kk���qpx{f��kW�R�O֑�̃ܙu����EG��8J��h�F+".����"�\����&�^GL�l����9�g&�'�"�0�P��(k�t��@�#ۻ+�Qe�;�<��줁�E���b���b� ��օ!���DQ�w/��2���n.�Nx��o[g>
5�%ؕ���<et@����?p#]c�8�?�� ���C�SO|�'��� �5���Bck�2�H��h۬7��۾��e����]�����+�](0����6^�����C�m�l_Kݖ���P���?�?*ؘ�T��SE*�8Q?`�K�J�̳����me,�^2VH�m<�k�����D�Ɲ�I��f^a`#���r���2: !Q�A��vy>�z�^Y�ب���lXX&
(�&�d�K�}�u�w�|���9�]m��qe����^<[�	���I��Q�Z�p���w��b:�9,�����0A�PP�/��Z$�b�5ӵ��U���t�gðh�� �rAoX���X�n��=k$"�@��.��;��}ۍ:�gg'7�������	�l�f^W:�j�����_&� O�d�z�v�T�&M�	��0O�y�Y�l`0�b����-]r���vJ"><(�Y�^�V[J6�/�x���̬͑P\M��9� L�9�k���p˃�a6��O�^@B�|�'rg��%�j�ʩ�����a(�.���>2s1@4��ێc�߼:�m�]�5���z��u�� T��jL��K�kR��ͱ1z?ݲ83}`�+���E �D�~V�	�����NΖ:mLƚX�����Tx{˛���3�é\]��O. %�ͬ��'��tֵ�5՛'0<F�p�i�Yǔ,��a�5BpC�!�N
�z��r�X�j��A�#�0$�Hv4��f �b$b���*&�z��ROY�E� �+�mi�R�E֖6��G%@Fˌ��O0�3�2ꎆ��b��'�j�i���[��r8I>�'�ߙ������"i6����tڷfuܥ��duK�	��XDV�G  �4�	�m3���ٔ���A]��QV����?��%Vx��w~l�<�X�%����X����,,���R�����c~�F�����,������@��PW�t���*5�-�su��H�l
��bδfz=+�I�G'u���~��A��7uϧH��X�Y`�+���J��`�:�+�"��mz?#%���Kp�������"L[�8���u� )-݋�����#h�5�?\R1,2�Ж=D��)�E���&����E8�S?Oq�����F��+��h����6!�)e�9�l�X%���ʾ� dK�;�k��H�h8Om���E�"Q�^�@}hw��(L�������