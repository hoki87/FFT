��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#�����~H�����pl�Um�v:��L��Q����;�~��?U�b����1�w���`� �2����:S���Bq��6w*��v����m��<�,E�H����,�b�M��1>k�^��&�SV%�n��b77� ��������m?��8��O�07�����v����-��Z�h�-"�f����v�Lk��em.������~A+@$���V�����z�K�Ex�;Q�2���Ij0�P~�ZR[�J�>��As6�a�!9�D0��c7�w�䔋G���ITwߦ�8k��i\˧�Ǚ��3|�İ^?��g!��
&�GCW��'W=+4�E!X�m���,0b�f"����h��D�z*�s;C�w ��j�4����w�c�3-[���:}��J�0���Y�&�ɺ�ӗJ��z'��;e���捦_��� hh:�z0qY
�P,{H���y�nS���a".k�F�p#kN64�kjt����^�����?�R��u�0��P\���'�R�+�8�=Z4�o���+�&d�0����x/d-0�rJ�'�a�v�f\�%�e$����D�ɛ5nq�Jjg3g$��4w1�:��a�D%�U���q0'�"�^�!7���^��bKU�;�v�}���k�Q<ⷯI6Tl����C$�2^�t��޶���e�����]L��e�P��Hs�6��ꥉ)������[�:���򱧇V����	W#�=��؉�i�{�yE��B%r'�P7U#��soe�f�x�}�v�&A�'��#ˬt�q��_`6��Δ
E�Σܫ������R�{�8���`Yc�.6H�Z?�^�9ҏ�.#�����E�rE�T*iD�0J�#����Y�c�rT�3��K\SO�������e'f¤���׃mSU�b�Y�߬3/���A���Μ�j�!�a�ڻ#�K�8�S]�����iR�J(o�l��P���t�����\� D���"��NlA��3>̵Gi��T<�{��h䈚��In�����y	FB0b�}�ӯ*6h*}�3I����z|�eD8���ȇ\3t �Ø�f�?�JPo�p�#f��3�k��M��QXAn+�j`��A"6�үa� ����Q÷U�{YK`��_B`�����-���*�����~Y#_R��u���������.54D��D�àM����dB �(�V�����%�����5 a��gQ���� �1*.�~�+>���@de�JM��$�|�+�}�u,!��WR�?��������r������BC�B�^Z:Q"n�R�	�� ����(�a��=���UlQ�����F [��E?t� 襢�*ɪ����Ƕ���T��-��Y�������!\�����t��O�?���])�S�$�<kG�R~o��3_�x�1m6��׶��cBZL$���ʻB���[$r������;|Z��ʕ���M(�|iqP�8��,�K޾OHtԻu�v��z�?�xQ�)z$jH��p	 ��8�dL���A��U�]T�4�݂�������;V���}yd��]�*9wZ��х�G���������HN�����bŅ=�!ѸX��T���Il��[�LkS�s��l2хo�I�c9�=W�G�����f�W�o6�^����[X���������@��k߁���9�<.�d��ϸ���$��x'��'�Q�
kqe N_��Ƌ)��(T�I�%�t�J��p14����N'00���n���sE�-	�'�Q�6���������B0E�CO�ߩ8�P�pW�aW9	^����_��6�UFj �S�j��w��5�����σ�k)x���}k���(W�=���E���W��V����u`���=OQ�����"�o4^���릕7��,ѭ�g~�?UHP����K�H��P���齩��J�b6[y��o��P�e:T�jLF9y��^+�f��Ǡ֡<(k�U��Zb�l1����}�|a�VVHx�)v�b���aM1y�rԓ� 6�h�&L�ӝ���*�}`�~���ڑ���6�n_k��(��X�v�%,�����%���~-�$�Du;�n]R_��$�}�����-K]��*�f�ǒ_��.i�>O4�S����R��C�܈D5N��v3��	��vy'Kp��(̄��Ё��D�z@�=�qa]q0p�T�QB9�A��՟�?��+�b�P�4�*|�33��ܦPIc�(�ST�2� �9:��i;��<���
+7e�Y6LeDT+h'ʟ��9S��2�g�B�H?E���H�rԏ�Ǿ݃3�ڏ+pJw�HԹ4k��3���^� nx�B�QF�0h�'�Q�w�K'��e��B�d�n`HF�	�����J{d.���t�?�`,}WS�`9	��Cv]����-��2lK:ὑ�<�<���k\x��(U����ڲ0�Ayb�cHFF��YxS���'nݗS�V0�<q���ぁf{�*~����f��ğ��?�2Ɏ9��2&��ȖV���"d�������هyf�T����g)��!�y6�50}����z<���wY��f�
;L�G��{I�=�r��j�a��R;D<%AGl&k�,�����؀�	��=����v���a������א�6�FY�2�%ٯ2�Ĝ�c�k[X=~,�J^��t���$)�v��U^�W�P��k��}z��z������j�r�uFQ]ꦹ��.�K��ͫ�J���fe�BV�R0�'G�3C���T���Ӓ�0k;��yi�uP�O�����ɇ^����4E�PzY��O���ƈPz��l��{r��h@;k��y"%�=
�?v|���P!�CѪ�}�X�0��.���6za)Bp+�wL���rk�6I+��Hu�Ip7:��F_&UL�y߈m�_��{�qNl�n�d�)��<��Z<�a�`z}44�VE;y���c�X�@	���j09V������5iZ�e}A7���Tk<�PM�� �]��
!/$C8�#��v«�=�]��t�����S�<ة��<)5ct���7������P�ޓɺ���I����}Om�D�>�=8�NY���u4o�z�ޑ�]M˚SJ �P˩*�o0��UOi�˖}B:Bu����K�1��Q�<2Tkr���4~���;ԦuTߛ�p��+4���ݝ�v ��}��D)�/��p �ڠy�ZO�!���cE�y�߇k��0o�~����X��v��&9�J���Oѝ��x�H�;�s!`;�܈-}#d��0�,��Z'�7{�Ȋ�.z�~����1�.�fv9vD߈UQ��6�Ї΢�����`�� �=�d�!C0G����:>�D	!b�H
5�;� &�2f:b��å�\lvq���Ϳ����"C��g��4�򊏇(wd�4$$��ERv+�/���5���=1��o�U��WeS���a��Hл�i�����X>\�L*wk�P��w�i@��Z�fa�깂јH��9�7��0m!�o|H��7������55�J�V� 0
�Ǫ@
������]L��a��;�jѵ�	)q��0�S�X�2tC�/1�!�2i������	h�j)����L�:���yK�;M�ż�W�O�x���y�ٌki�z�(�5έ� Nf�?�ư(�Y�G�9f���A��~�O<du
s� ���`�����C �	�%Ա��ਲ��5�����B<�2Q�gW�~Ψ�;�u��И�SE���d�e�v��6��8l���3Ƀ�Z-��J%Ȁ!Q��K�ݳ�G�
�k��a�D�@�F��g����M�g�?��Mx�w������Z�@fUb���9(��[�S�3&.K?�;zxm������f�&��Z���� U���L�2�<�"�q�,$5Њ�=xD�@e^�m��EE�0��
�Ba�!���t�����|A�fպڢB�����˧ǆ�]�b_$���*(���Y	�{�L���2�@$�eu���aF�Ơ��#U%q�k[c��2��*mU�ي����	T�R#<�~�!��pE�Pf�k � F��uF�`�:�L��C���Kq�O��	���/ ��~�Qv5����Ѷ��@=���|�/�(���I��6��"����:u��.Y��r��C���喢�K�������}�zb�Z{���E^|S�?���],��ОPm��|PӋ����!�1Q�4AJ=nE��Nn��`a2�);��d����C`~�Z�F�N�H���7X����"@�~J��p�1��w(�8D!������=inCJ�cY�>�T�6�%�!��>1A�r�m�>��O)1,QC|?]2&��ݵ0��G�I����bP�V{a>��w:���5咸v��yCB{4�f�`{����>��2Y�Ul��F�1���4�xi*�0�;��O��2��%�m��Vp޵>{���\��g�L6%R��8�܄CkTs:h��eV�Y�?��~�	@UB����S����AJ���G���f�a�'���0R� ��}A�Q��	���Mw�Zʿ:���0U�7�m[c�$4���ᰫ]�����m����! �zW@|�1�����!.lB���@��Чf}nzXQ�ʋ5�7� 4�*w	0��)F�{~8	;i�#J-yfl�xy�HҶ;�-�6�v �&�~!��T�Ą-� ?��fq|���1[���ѧ��yZf�����?��!v�X-<i�u��vv	���`�l[���Ͱ�:PD5���3M$�y@���U��'�Q����7wM{���U���yށZJb)4S"�e�]b$<�=���p�tFl%���xG_!9g��d��Q��~��Ա���
��J�� p0��V�*��I�Z}���,0{X������>�'�d�M��#'�k���U�|�@�ޡn���"��2�=���!�.�$R��}r�&��q�4��pM�65\s!�!�R�0����-��1�
\�q&��2�3u��b`,�4�k3�f�֒��^�d֪ԅL̫jaza�P��+,4��B9�\������fjs�W�]�\� �s��Y�Է�k���S{�b�2@ 4�3P���,��\;�H,U�P2��w��%tL]ѿ��3\��B�/�fz�o�`�j��=����h���8��-$��Ѓό���@z���PD�C8h����jϟ.r��S��h�~� E+{q�8�m#�Q���'��Z���{�E;4�������V��?��Rm�A�ƹ�]Gi�%�t��'�e���
P�zN���eŉ�M�ZF�*��{�ԓ�����l�ȣ%D=�Z��dE���h��-����-7�e�oWi��c�[x��ő�2��<�����h$@Vd�yG��[{���T�_!����8k�]��B�X��tn�C�Cڶ�=ܪ^��+رR��`[��}.hC�ӧ)|��>Ƙu;Ǜ�����\3�WrBb�A>�J�`�� �;�C�<m�	�4��#{8��WeA�����<���������w!��&1I�N���2N�nA|
��m��!(���� ���7���T
LЂ���	I�}�L� $�N��wN�����5=�0}�D��6ZRe T�� �'�/y��r	~vMqx� �A��I���0�� ����NH$E�_{��N�({	]G��	"�a��1�[̈�_xؕA�v�_!���α��0���"��:�M��6�'�b�����,#����l0��������	k���׷���wp߀E&m$f���(�U(Mtz��g.�
̓�/`���4L�|]�:Y�^ڄ�/��+�KV��*���U�ĳƏ{-v���b�K�/��*���I�.nRX@��ͻ�O@�~�,g�Y~U�ö��8"f��M�C���*F_eT��ڒ��\v�;�t�-� m�0��g&"|ڂ��e��3P�~����|\죆��d�� ��&PR).O#�����@sK'a����/`en��V�a�LEs�c���!8/�Y�U<�'��z(��������K�K�V,g��]g�`���3
���i��]�j�&��b�Cd��;z>�ڏ��Ӏj�
7;P_�7�<�}���Jr8x��C����|M�]~i��8�ea �����F�Re;�2��g�	�n|S��#���m�D%9�!(&
�����nA�^��A���0�}:��"�<f.�2I�a@/�K���,k�.i�������Fr%�,��ݱ�\�g�еf`��<�~�CcLL��k��)�lw��_X��VV�J�O�.���ϳJ'�e�ڽ01�>�G����,��V���.܅Z]�3)&Vca�us�	�L�l��"zk�u�z&�-�h��)Y��=���6�F��F��q���!��"��A/S6��煉:��f�^P����K��x�/���������o�~x�<����V�3����-?�@4�����'��NߨU<bz��*���Q�+�G��*�G��W�9�{3�H�D^�$���ju��n���;�uB/��.0Q\�5Ose_]�����e�X��;�;��>��P��X�a�e��>�dH��퍴��9�ZΡ��Zj�� ��ˀb�r�(�@Н#�+�'=9R�h��j��~��V����9� :IK��0Ձ^o֦���#�#��m!g� �ˁ�li~X�Ī��~p�Hr+�(p}���H!��f��c"|�/�=y���B �2��"�w��љ�Evb���1����NN�o<,����Q��@�(��y����u"��?!(W�+�}]d�L���M6����28��UQ�6u_��P�L��g���Z�Ny}�м=r��B/��4Nd�o�˿�>���'[Mݴ=��=��>�X���i� 	p&.�ݢu��\W��]ǟ��8潋~-���N�1r$9��Z��[H^�NV�����.<"WGgH�%�g��ޛn�5�$��4H�A[���ům�$H�y/Wp�ע׹7��7���Y Z�Z�C�=�cD�j���>;wp� ��z%F9����p#�F\��^���Q.h10 *Gbv�>���Y���Yd�N�]�ɭs�k�'�d{�&;m���]� -b4���XIL���e�5,�*cnܱ�t�{ٝ ~�����I�6&�&WY�V�\��N��l��<���W��z��Zc�G�s�oYz����]� Ю3�*{K[A�N���©�O�7S�^m��Z�3��%T��F�p�O9�Ԡ�gRsE�Htf��h��.4'������uz�5�{�Ǫb��,yԩ�7p`l$����ˋ&��y2ڥ=�1��:q�4��[�����~#�I}��Sg�}���~�j��@xg��hȆ��1.�'��yr�c	O�b���}�J��zNո�`��!��/���ߍ���[���p���4�}�*�p�?���.�������o���eM���V�U���oN�Uy���S3�g:�"ɂ&e����=�Z��I���)��AsM�Fg |���P�7s�~@�DՑ������.��q�1���1���'Iw�Өɝ��d��q�0C4[��u��a���nQO\�>�\OB�n��5��,�vO)i8&-]) G�Gv`��r�Kg��C��Y��)����Ǥַ�o�Dn����ǹ�Ͳ볪{0��^d�Ъ ��S�l�IM�6��A/o�����ܪ2M�&�п}�
gsb�[솦F�ƕw��/\���v�1��}J�V]ֲ0����s����CC�m��-�v�;A����N�p@`�զ��K�WU�Wl�p��]�jq��'Ru1晍n�N�E�'4͹�P�;y]�l��"m����pT�,G�ku!��&�h�]k.���?����ŵ]�1�����$��Y���p�O5�����ѐ3���ز�!��ׯ�؁Νl[�]m�r�@�buh6.g`Kz�!o<`�Zfqʎr���B��I0��O-!���܂���[R�N������.#:�n.�|���gc����2�&a���	��d�N��8|�%sM��S3�I�|(FC��*��ǃ?����}ߢ��aS�Pt�bP	N<-��i��ƫ���ƫ� �AF��2!�/�k��5~�,��t%\`���j;fG?+2� �o
���'ϼ�$ĳ�LքC*�綇q�IG�)r��X�L��s�BP>�殰6�l��&{�B��l�}Zm'�JW�4���Px��Oc�"j�zؖ�v�Y��Fs6�Y��4�������/�����4�k�1�h���A��Lx��We���GX���,0q�j����~���Z&������K�3��� ~�2�]ems��E��%�q��=���^�cd��H=T����ʍ����"�F~׌���S���^�k[�bd���Mj��%��F��tue�ߑ�I�V}��?㟶����V�OT�<6E�չ�r�;���y��Df�D�*��=��(Dt�~����Fo��<�H$��W��1��k��-e䷷�p���]�w~r�޸�p�Y�VK,��D���5��τ
�L8�Hl��37��E��f�&0K[�7�ڳX���E�ɾ �B�#��&�� ��i�qHU�mh�)ňF��^psT*���?z+��)i�������SU����#�|!��&�^	z�6	�&̓���1�>v1r��?�ə��� ��=TO��u�{�No_�TNt]�Od��k ��J���@�DB)���P"�����[RP��g�b^��R��.�xY��,`�5ВC��zc�n|j�5(��7Q.c�Į����Y?cjf�n&�3$:������I����~%�#�~�?
6�Fɪy9C7�jFP���猱|M$3(�4,��L�j}sn�nZ�6@�����i�Q�����-��s<I����s��M���6̍phX86�1�\`bv���\�`F}�D���b�ӯ?БŌ�a�-s}�jҦ|WV~	�c�����b���%���ڸf���$i���&�tšlɐz=���b��q[�`5��$ܜ�n!-��#6�v6Jpmz� ���f�25E�`��aX�x4(R|��ϯ���m��~:��� �p0��,-�;�
r$��(����g6I�=:���W f�7�����Pxu�6[w#�!�v
�Q��|0ceXC�y3����%G<g�܏оH�[ðҖ�m9M2οP��aIG�����_4ʿ4���1���xk+p�+t���V�{�y�h��껻�ꡑ�w�_sb>�G�1|\X�`9`
C��]_�򗬏Q����B�j�0��/��GK�yj��`&�g?Y�T�ᕈ�T��{4������n:j��-�ۀ��U��O�WɵY��e�|k_\��C��`�����-/�q$��&��I^u�� /����u���"m*Gb��U���f�W�sѮ�	�k�:L���j߼�	(IՏ䑛۬�/��Z'��D�Ր�E�o~V�t�#���">+2�nKq�C��l�Y��a���N��de_aG@}~&�/�ٲ_[��4��q�^Z��B�ϳ5�ab�'��ۂ�J�w����K<��bk����-F߅� #��'$ⷊ^����˄�FE���|f9�}���ԐA�����t�5���3;ƱE(�ߢO�Q��ftZ>HH��(�H˛�)��
A`������9�O�n���5�w��> D�r�m�oP�=�c�#	i�P�]�Z�G��l��J��c��9fF��օG���*]G���3���+R�'��X�<�IXH�[��Uݞ�5L%4��@�����I�H��n~��B�}�0��4��1�K1F���W�2^* �����t��YX���=퉉:H���Mj�n�s��g�>��e�-zU!-7�m�a�&���?|o��4��ο�V�Y�3��4_���������7&�YD
HJ��@���0�ƍ�ud�x?��(���T�Ɏ��0~s1-W`ִ����A�ͼ��߇~����d2y,�E�o��Q��?���8���z�;Ej�TƎg�xnw��gݱ]z�(r��zx�#�@���~���>ݚ|�Ӭݽ�Ơ=zeٳo�D�e4���*�M4��Xw���JN�	9�ל�l@ +̓��U�Cڧ�b��)���ג��<���DnJmRyxp٣󂱔ǟ�P�`[����l9� ��C �#��ȭ��_:�|j����KB+�! 6��q��:Dhl�fC�;�lC��Í=��+�-t�9R�@�e����4�<�@ζJ-�oQ>xM���p4�y_m�A�L%S�QKwO%4ӝ��A7�n/�jA�j��`����Ij�X^]3��5�)z�g��l��}�j�s�N�aw\�8��m�<������5m�����/��+�,��3I%���e^:��=(�k�ח9��\��ړK��nw���28Վ��М�N{���Ͳ�dF��{">1 5A���Y �G�ë�r_�q�K�?1�h�=��y��9�/�o p�ߥ�;�e�D��#5hy�1݆ Qv�DF�WF���,Il�H��U������u5k��ъ�<RDD4S�[ڭ&Ce�pd/Pt9Л��Z]<H:9���6�����g����$��g��9�7�mܿ�{����)�6������^a��*�U�fB�L�����K��c�y�˞�\=2t(y�XT��fo�0�צ�H�D��Hqo�6�����E�2y�K�Ҁ����D�Ȇ�w�Rx����Z�����+�L�h�Yn��d��5�lxY�X�w�L�  BC�����(B?�h�u㞂��d�'� �ɹ�l��M�G�O�\=���m^_XƤ�8j�o���+�v�݅f����"a)�d���ŏ�Y���$ʯ�RV�e���N��Z�xb�L�V���q�B�	K����GV<��O����)�5�7�oBޟ�`�K��t"o[���s���B���P�<�=���6bi����{4Z&]E��h2F�~��n�����ٻ��Ǆ/++���ْ�B�ȒyLP��gBsX��>���b���i�������%cH��7$y�$�*Yq��m�J��Òd+�Hu{��*u����1>����:6�/^FB�"��VN��֜�_�2�-�n����ۯQ�:�~3�]pd�CXƴ$�G�$���G�QO@F�z�D�+_��5�Y2���M.��ϭ��ï���ɠI6xݖtY��rļVs�8� �l������]潠�c����!t���;ڔ<#)LU�[��X�G���I�}�>,�iz��;��(uE>�m�\}�L��a�Y�j� ��h[�ؤ�BBO���q�Jg���(T4�24L4z�[ԓ��5�W,�W�&���^��-��E��$��Z��-�$��N�/�������2;�C?�@X�-������p�Qd�����c�(4�ҥ�V�#j��!�i��>�v�C�R�3�}�n>t��{�j&Z�2��B��˼%2Q��g�M�ay�o�Ϟ_��
���>��0�}UzE�P/��ئ�SVV����d][ʣE�Y�Dk�k��&�D��칿&��f #*p�����^�8	\G%񤳣��,C��O7j����QQ͔te.��pi,K"8�8���	j�M�_o�P���V�
������MgL����=��Hb�||:��	{Cz9�Y �mx+A�)˃�WʫAڬ�y��}`�����"a��f"�\����zw�t�����-��7�vo �f���7��fs��x�fǨPZ��R�� �wV��9Gr'B!:�^�*��RR`\