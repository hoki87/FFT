��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�#&��#�<�����)e���0��q�=� �%e����j�I��4m��b�����u$���r�}s|Ά���EF:�t��c<���n���b}e���p�xn�����V �`��H>��L�F|�җ+x�࠳j�A�I����P�>_T��i����X`i0��9m�\�I���Y%�:��2�����Ґ�����ˇ�f���F)�X�!X}�K	�=��n�1�2�.+*���50��_���e�vM���Q�jA�;���p�w�d�e.���%	����/���}�W�s��+-�a#oZ��b��BB�&�'��A	}s�3�%b�-����?y�(XK?�	1"����f�I�����v�_WL��}�/oH!�ʼ����:%��$-��0�'K.NW�Ù0'R~P�{N}!,`Q���J8���[0&��4�laz�����+����U����rA�dovr5��[H���A��l���UCw���:mY��DT�`�v�����_VFD�x�Ǜ������dg;f��u)��Ǒ�=�T��������{�����yl!�d\�EU��Ǫ��ȩ�y\�a]/# ,1M3�P�T��?��c@�Hw-�@Ey$Du�L�G��9�d�@��|;��l����>�:og�h	�H8gBĩ#M%������Q�T��JO�Vǿj,�1�(Ъ��D���l���zӰ�N���,��A����!#7�q�r:q$퇳=z��=%]n5�U���;���I����搇�G=�-n|��|?���H���:ʴ'z֗���(���9��fV�����^Sq:�r3��ېC&"<"� Ri���%hl�jG�>&���z
&8/���	�5�J�!^��,XC:�{WS�� �E�!~2^��5|����]�*+�WXJ��^VeC�6+�C	��nq^�$���t!��'�����T���M�6g�5��"���n�N
c�]���_wf Q�d	���a�L��vH��z���/��C��c<���N�oQ�\�����z�q���;�J)���tE���@x�ǛZ���`B��PΡ$�}v1Y�2A�& �;���k�ck��W����=�g�H:,����p�ۭK.��RB���ŉ0H�Ȩ9���/�f�n�0���P\U��#���oB_z��z^��tXe<.�,G�e2�����i�V��Rc&e��6�HP�̝ 69W���	�^f�Յɳt�p��V�O��<��
.Qi;��o?���R4;���Y`BBLNN�nI��L�j��q+���MMy܅q�U����v颾�ྑ�\�?�9
���a�hj0�aZ����N�EKx�49@�|)t/�/��Q���ba59m ����i0�/�~�'N1HN�V�&��m��DlZ��xT�����ü�u��>w-t�� �����I"#�/���ȵ�_��o��@{��ǂ�3�L���N='4�%��K����/��7��.T������7f	&D���1[��2��9�嵱v-�a�י� �|��A:���6�4�{��k<�v���+C��\�0gD���K��eq���ǑAg{���׿�Q�hY5v���G��x�m�S���bB�T(�\���#y�r��ͧJq%;l�>��Fk\M�Gn��
�JJ3���R�:T�����E��.�ŵL��F�|�e�"�ɟ������ࣾ�h�սU���"ij�=�)8R��ۗ2��h+���F���"S���HF�~7��>e:@�Q���E��l*�+�������3EJ�O�@���0y�۟H{{�&1�s�i�NQ�茯m��л�t\�ԥ`���F�����C�YteDm㸟N���g�"x��b(��q4���-�wj-��.Z
��[?*��Kf۵��6�#�.~�N[Y��
|��)ۺ�W͚}���%�7fb]?B��	�
8ͻǏx��Qw!"ƆK�.��?s3����>��JF�w���ˬ;����!�îcf/�
E$j))�D�]�l�v�՘j��w�Af�E�t�nY�KJ����ceqɷ�e�Zb�U�PE<B���c�\�U�F���̕ư&YQ�8OE0�"����-}h[��8A�2�*����w��Ku��õ��+���uu���^���f���6��_�����ǯ�O��:���нF�SzoK�@��p� ��.������8G�̥j� A�.#CS�e]X������)��Pk�~	��d��}4Y�v���˩7=K@
���;@��F�WoI�����m�?�Q�]�n������Ԋ(�n�ǣ̲G����#�?� z[�;µ��
�σ^�UR.����-z���!�,"$W���)�z���?&u�w�٧�$rb�iy#�<}�q����~�̤<h�#5�%^8�lw4d��]�ɂ��m�Gh����"�$�F�o���ڽ);�Ǚ٫����n��uٌM�S>j�Q���y�(�˄�!�oɻ�Ì�5S͇Q!��2�~�����D�t`sj���Av�<9�+|QgpiO��2�m�D��P����A4�N�~�V��;&�<��5bw�&69��De�S����.�R�P�IT��GS7�j���c~�����p"��T�W\ $זgP�߱1U\�Z`�HDnٰ&��R[үD���(Gb��Hb�y.���:���Ԧ�+�eKƬ���KtU�����ث%�j3�G}&Ms�1(�A���%�g�,�>�^�p�d��+^��&�X����q��@1_f�*M%��pw�a�H�����G#"S� 5���)�6�<$W#m���B�"�E�.��^_�Gi^C�����<��u^$�L�lhɫ����c-�b��L�X�x�%!|����臦G��}3�^��k�DeA��/*zoG�^.��~��f@A�K�y�����[et)Z��_(�WmO��!6@��y� �HT�8g���]�fg3ɹ~���BX�l|!s�HZL�ϯ��Y���6�j��RϦ��"�5�g)��@dI����Q�S:�y<�Q�h\vjb��s�1�L0���j� uI���5�;����"��ߪ%z) �si��󘣗U.��e����ݪ�V`�x�M��k���9H��]�X��I (s,��	��iHj�����ΫN�\��(��D��I���� �R��� kg��^<p���M����ɠ����l!"�B�s���ۗ���<���^Hw�|�3��|
����}Zk�!� �����gA6�i`�Jù�G��B7�;�2,5(BN��Y���d�w��n��tH(���>��E�Go�U	Q+�����.sN��TW~&̬x�Q��Rh��c)���&+]KccW��
DQ�����~[$� � ������ËR�0�t�m��!'\�˚-��>ߙ�,B �n�@8�f�W�l�2WZĻ-x@��K�ި撚g֪ϝ7u�]l��v r��Ϊ�jUp���l0�%��J��c*�0/�O0��}�2/@/�-��,ޮG�[�'v����9��u�r�P�Thk�'.m0EW*��������C�]e�#'����o�����X�M[�RB���]s��Tu�M������.*��(ˬ|h7��#49���5K����dqvК�uB<O,|$e�}��HR�J��D�"�,�,��R$�Nnܱ��% B��o�2X�[�j�ŒSE�&�[����!��Ǘ��+�M�M��u�ӿ�gu��W�)��G��Qf�w@�㕇�${zT���W�w����+��V��S�O��@|ɖ���rc�X��0�U�ٍ��_��;��ViKd���qJݚ����� �c�_W! O6�Q#B��G��]�B�sP�ַ����un�G�G���5v,��@��y���F1e�	�{C���	-���o����Jh�<p��-1˄�yH0T��u^���H}U^��o~-���H��g�\UO��]W6����id��H|k������ݤu���;M�=�)QR�;��1^�����_��]D0}�@��)S�d�(0�90�"���-[@!6Pn)7�pq��� ��A��<�Ҝ��W���^}�էM�Jnu�i�V�?c��d��݁�{�Ϝ�)�X�8�"
���5N�����&�h��1x��+n���~W���� ��Brw�[ݯ���CO�����∽����~�64��3�G��l{m9��F�gC�.(�wuА���F�4����;�W�h�>RtMQ��I�)���A&�����к|�fBd!/�yA~�'!3�x�fH�O�� ��Gb?�qc�W j�"W��su�7���h�5�qⵙTA�
��5�� L�CvqЕ�j��"Oc�Ű_O�~��W�-�mr���<�HEסE�Ͻ_������t�w% ̀��"�M)�=�M�C�E��-M\<���qvP���0�W���	����z7`�n�w&�����!0��q}�'��D���8h�/����1�%M6T�L��S8���׽�LC2������Ts�b�oK��gD��GQ�����r�v�Z2��L���P���(����A���d $x �vBH3�]:! � 缟�g^�	w��T����d!�2U�y9Y�s
#�� *��z\�.�#qBTE��x�$��Y�<+YC����C͎�ݝ,t���@���C�[1�?:N�7�(�K�bTIˣ��V��}��&�C���]D��"��Ը�eэ�&s�e�����ǞX2�}y�p�g9��r�å?�%hNf�� �����0Y/Xi�j"���C���t�����ڲߞ֝�2���h���Х��7�;�]H7\�u�^�:dXQ��}�{���:6삛��n}D��	��.�M��H�d�K���{3P<�X�pW��� Lۺf��=��D�g�D϶���[��٩_!Z�}����'
Ӵh���Z/w��-|C-�x_5.�s9e�ms�c\��q�E�C�2;�M8����{��#S���Nb�a!�m�V���)��g�2*��e���uʟ��hV���A�fFg����gIm��J���۔�.���0�k�裀c���v�#���o5��]���m��B�_O;A�F��\�׆T�H���%!NVO(s��thq��*]�⫵O4T(T`���No����Eߩ�!h~<i���E��u���!b����=LT�Y^���o���3io���`{Oحo�B��l Tp����Ϫ]��O)d�F3�A<Z*y�:��7u!�>�8N��
�ƽ����)�"�2�*���*���&̱B�!b_N���YIx�X�2�/�H�ޞJ����x�t?v$۝@ޕ��������?���p6v��٣��LE�;�������Hh�WbN���1ړEz'�b��'��~#�=F`t���%�ľś�i�::�W�������
�dnxPC�,�{��a�ҷ����8�x��Y,�?^�/+�-Û�uǘ벍�k9�y�AM�|z��~Z��l䕈{!����1��?hxr��{R-��6ħۉL��YX�~q��2�Ƴ��I�;���O�~:W)L�u����h���|Ē�xOw��B��e�Zfܫ��yF�4�;)K>SK����#�dL{�P*�]�ZL��L��B3eR7�3�W���0��X��e��*�Ǟ�9jr@�/�^��/�!����n	���O�mFnN4�J۸t���.�8遬;2�[�o���������8�3�+��;U�S`�'��O�nC������š���T�����!�F�����g��M�4�����'e��"uW?Ԑ�uv��l��YTu��rt��>�_b���K6q3�˙�!xk@��yo	2��8��K-�)���ȧ4W�G�8��d�:0c(	���R1������]O|"y�ۭQ���f��:aﵬX[���6'�X����s?G�h ��[|0�6�vu�� @y[բ�@�CNx�'_�"�� ^��f��1f��>%��WM��$,�2-��KDb�B�)]�O�|�A���l)/����7It��4Ϣ�r%�%�P8HXn�C�7��S�IjQ���W%�zr�0�Qo�wӊ���?f<S؇Il�!ý�Q&A������O�e+��8.�2c��w���I�P�>����=S�J�j�K S����R��K��w�,���k 5�[�'�@!A
ٯ��]�a�Te(T��"똃����Y���l8���:���&)�B��{������<������x�Y}TDɨ�e������R�؄��(���Q��4R�Ѳ�L�D��(d,�3{�k�c�؝���4��.q�Y�*��Z�$r��6�	/��?�?1Q���>W5�,X��Q�a���e�3MdqAZ�\��^����eI��呴ﮛѭq�B<@�fy��!VQ̚�Y�́�ێ1��P-�������#gjk��t�3�����Â9�Ǘ�Z�l����V95 ���@:w�F(�y�u�A�j�"#�!����˴��G���sƅT���	�q��\���A;�-��y�m4q�1 . ���<iJJ���͇v��hdqE�c� �6ݻWj�y�J�"��E����'mZd�,���]�݄��Č�q5�?��#B�}I/.�^�_p�7�#��m�bP����c�ܐ���;��~�����5����U��Bc�y���|��5ڢ�J ��:��ڎ �s�6���Qt�&pv}�%��9TE�o �4�2���͟�sŚ���,�ϰ2ݪ%M.�>j��M�� �y�� �@퉢C%�Y�;��a�ղ�
|qtŶ�?�)1�$�R/��+-q�~�qkN5֙il��@
NdǟR�)O��!*�q�Og���4E��k�}�m���׷6���o|��U=��l����Z~(���à��Y�?�s��{����@�A�H:��E8���64��A�W�Ǯ|%~�	���F����pY��L��٤W�ڰ-���jR�	�nB����NL�J@VG@�4�s���ql�x��}���X0NKa����~\H��xh,�A������.d�"���<����h4(�F��'�˔&}�7��Jf�w�؉�BI� ҪX,��?:^r�ҩq���\��e����)�B5*���\CA��Rt4�lGq`{��?A}y�������U4P{:�Zu�;~s��\�&��i0B�2��(?��1��d�!V~��͙{�/�F��G2����}c��;�@�ڣ��K�!�7�I%ɪ� p��	���+����b�kg!�؅x��M~n�+J���uWkR�y*��	J�����Mc�|MX}�����&j6p��ĭY��,](Vݩ٩2;�=8��  D��⃜~[M��U3ŝa$�����yǒ����n�^d���mYA��'F{20�:S��d�u:�v��a�i=(%���? gO/�chT���-Bd�}l���n2�E"Zs͝a�JC$�#��/߂&5��@�Z��{��z L��W:��hj��P@��+}&U6����2��Q�=E�N�gO����˚���=2�+T�f�}�ksi��_"���I,��m�L��c8M��u��%֤�����I���MC�17!�;1��9�@��c3LW��A���UO4k׆9S�����y��o�sr�*nS���TP�5�e�*���׮gS}����G5�����M�R�rr����Hx%{(�r�)�.���耶���E�]bU�37k倘q�cY��[����u{,��QhW�� �1p�i�	c�>f�b4ߐRoG�HlG3��g���fi��[�*���<�@�H��KL�p���-	���*�p����u2#a�p ]g	<��!t�iǻ&Ҍy�����7&���i�_�@�=�o|�T�Y�\/<��I���6�����P�~T\��Gӽ�P#/d��E�<ԥ�D��?������F����ë�FQ�!�,:e:�*|��0�졕>V�Y�+�)�6�����-��D���XN����*�Rs�����kT�C�v��Cg?��ēh[/����s�,��Z�f3ֳ	q��jNi��݆�����m�d�ݮ�Ƽ�:Ud�(�9�}m\Z$K&*��^׉%O���:Z�	��ߠx�4_*6�e�i��S�oo�0�M�##�m�*�n:���^��{������b��db���]�f������̏�8����V�G���%?�UlRT�����]��e����0��9���@7?��yZ?$)�2f_x�,#�r �Bk?��/,u��|�m�#&.)���`��ǻ��'A,*���K�S��s��o���B�����������[z��DMن�3�6��7�[����n�����\O���n�c;l�U5���˚X�F^J��غ�y�*U&k���)n���t�c��⋌�g�Y@(Z���$����uH�` s�����D�CZ�#�n�h��&nLEP��6��]�d3�L�v�Y0��]i�����xm�?�1#y�7���DO��! (0h����2�=��\^W��k��r��e�?��X<�n�t.s���H��> �%��j9� Q�\ܥ��W��J����dp�3=��h�Đ���cХ{��6��GX~�p=@�z/�"������@���$���0�u�����Y��W����	wTл��t�v�=����g�Y�.�����*x[e�Y����7Ww&wo3�p����,%p�X��Ng�O����#QL����������&Q��eDL)Q���F\�� �M>���}�Q܅Fʱ]�v�aĪ|X��%X]c�㬕�>S^��]��?l;Xy5�#��a���򉟈}�љw!WK{�6��'��E4��G_�aq��e8^S`������o��n����aN���Rl����,�ޕ�W_Q�X�J�̕v�Հ��Y?��]�8wCf��ȴg���~e���TΏr��10`����.�6O5�Z���
;�AȰ�v���?�M������c��KM���g1r�8C{�c!�#�zz�\�,)�;���QU�� �%i�~�M���N���:�+N���U"F�ڈ �D1U�R����3�����D�T>���d{:}�2���M+��bŨB���j;T�s��������[ߑ{L�*��Ny�\��`$���@)~�n�F�j�_��q���ޝ�x�E��j�j��p<�x���]�Ӣ���'_�@L�Y!C­�'�T�0�]�0�؋]�j�?0�YZ�K !��,h�QT�!u�R�𫉋}Y�e�&0d��[�n���2Io݃������5��ā�������:Η��9햛4��>��к�x��P����n��D&a���:]���6Sq�
�Pv"������+!�Әh�^(�,u���u��L��{�O�lf�8�������W���[O��'����9x���`e�1�Hm�5�@Jd-Co���?�o_(�	�({���W<�t�j����y�L��E���`?�ە�?85UIAV��b��^H/ì`\r��o���7]:�-�W���	�A��Cw�fjO��V_#tH-#0w����h/��J��s�A��f.=/�~��~=a�A�?G�]�@s����'i�7��pl�)�
 �lY����-�_Io�f�M�{�k�L��8db,���ty?^/��L�9�SFg����1��A�!т�#��:��gRb���0J�#q7f���Z�J]�S25��_-Bv�N����W��b�c�CD�W����/}w����?"pw�C�LJ�=��@�zeL"Tvz,i�[mQ�����|�Q��k�v/7k9�?m�{Ўz?G#�?L;�!yc�6�7��O�.���Rn�&P����J��kB��T�9�l��N��t���J�D����z����Chh��A0~F��'���<�hV�۝,g��Fb�3�z5J|��;k|t�,R�lS�epH���t�"��j|C��B����T�+�p>����W�u�u6������f��l�ipY�^9 e�ɜ)ĉ4<B8b���q����IYF]V#������t)�0K�����`��UY���#<�ܬoS����.��;
���7ȭ�}��uo<qҗ4�+0��ng��1��c3}��������%��.P$�%o�x�q���F�+-W���0S���:|������6�G����?{E�.���C�]�ašD݌c�.RU?�M�N.;�	��cR��8X?���l�@��)#ze��ӟ,H^���G�j�DiD�W=.F��68��Q��ǝ�dDQ��7i��k@�O]
?�}$O���Ւ!o��}p���7�>1J�c�U���C����O�+�͊!�h�	����=�+�PD�!�8����t|�X#�m�H�%�/��z�F&ϔ4�V�~�g�����p���dU#�x��s��hh���&�sl�ʊ0��+��Z���r.��%���W]:rB���y�j��R1ϵ���T�������M��pD�`"^.9Q{߽"0/�@�"@kb8f��ء~�5c��7a��V<���h��>x�\"�Jx���ܵ�zõ��eٰ��Z������{{�?���3{�B�)����/>������K9- ㈍+�%��֪L߼��.)�r�
���|	2Q�m��2u<7J���3�X5�}ZR!^u=q]'��'��/�2�*�гe���<0��aDj��:XQ�wC|�|k�ec7`����^\�z�<������G�j��縈���h�m����@��������