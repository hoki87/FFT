��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ���������,C2Gz<n�9Sm�i'y�������4�н|�	Υ����AȤ�Q�O��uo�3d�YƊ�d9מ�{gJq�A�m�����g����r��r���ں�}a�����k�Iy�@b[W#?�ߎ��(Y����9>�Ej����
8ǚY#�5cG���������D��awAbm ��2�[�W؟���ٙ1�?���c�OQڸ0��c������� ��m!hU��W��z�������Pcq��*VD
�;�p�b�y�W!aU�i���H�jdT��ɉ�D��-z�2��#ms��9���[�!%��h�)@��W>�}=�B�g�&Ut際Y�߁�\��1�ƴk���-�ñR&��B��y���ڴ�N�W5U�����^�]=0���������F2��'dFl8��ޭ���� |s$N���z4��y�nM�Xq�4�� c���fa\��t4��5Qh���h�����wK����:��vmY2|Oc8��.�:jHs!bda՛F�J5��Am��@���;������0��� ޣ҆�^��$���O�Z�N�5;r��l�0�R�Gʣo���u67o�� -��je�l��n�&!��.�E`������]8�#�=��T����� U���_u#�#?����AQ������6��0'w�+r4]���sy��>���	
�*��e�]ډ�[ ��W�Pjpc�ҧ$���
'�&��ǫ��o�m�@�!{�P5���JU�k�w$v1nUI�p��/�)pm�LM�ĒE���	u���q�a�@!��׽Y�����[j2���o�,Y�§����MAcM/�7��4�@��hMQ"o��D*��[�G�f��r޲�uqUf���,5�9�Ruh�;l��p��9�Z���²X���v+U�g;����R"�|�ŭ�����q�Q����{���zi��k�� �:�!�~8JPY9L��ڟ�o�����q�$<p�1S��h� ��4�F��첍%\�F�ԮUP��ku��ʦ��c�>?:�hy���1rO�ԪF�����@������1�!��%�(�zd���,K��<'2�V�OϺ�H���"~+�p���{	���0Dd�4�V��;�v�H�����s9��(/�&�kv�x]��L��h��"��6���'*bD2듵�ě�4ا�Q�Dz�;^� �"䩧A��5N�0���X?�ہᐃ"�h=���&�vgI���k�����m\C���d���i��%��CA~�����9@KC"Q�
��j�*=r���d=l?5U�7���6��Sw�a�mf�o ,Bs�t���E����N3��70:��@��ο,�!����NT��~n/R��Q.����w��m<��_�^�C��0�`�඿L y�4�X���'��/�u��Vw��&0�1=đ��.MXUn����Gd�p)�q�n�O���Z�p��:$�ё#����#��6z�'�n`�E�߰U���T��B�'>j�Ri+�q�I��hs��*�|S�hҼ{]�6���H��.�����="bTi���|5g�v`��F��6�Π���ECjZ�jѦW��N�FnZ"�{����rj���[6��03���m�̛��M�PG�	5���m��yE������r����_~�W����w�XϚ�|���}]閁�DP[\��d���)��\Eۼ:��5��wZZ�-�����J�Ÿ�?'��@��=��q��EeG!��҆^8�ybI�2<��0lx�ې���(�2!�x|*]v���N�U�e��������y5�,����G�.g����X��{�-⠀V�~:��.A���0O�������N�W�/�)-"����)��l_S�9�)j/�E� ��|RM[/u�hI��O�]�2f���-���bȯ~'��»d���r�6�_�(#|M{ Z��H�3���'���ߐ�&.,����F,3�Ä���P[�����ʆY��ܸ���v��<�p�����N�|����a)O�Kv�.�����V@t�R�0����V��fYF�~�4���R	v�p:��y<���.bTV��g�{���"����<�р-�o����w,�T�8�0��(�Ke��Q��	����C�/HJD����8��_O�)y^1��n��cOT��ѠM�����y _nQ7��BL4p%�Ps�h�oq�	"�x�x=����I��=_<����fn�ť�,������'=�K.1a�B,HU讦!�_�����s�J�Ԛ��pD����� �Rk���̖�B@[��V�r���%��Q��ˋ��r�`'��^��6a"HsK��#�`Nє���7_<>�k���8�&A�I���	I���!.2��R�o�B�T�p�\�N��$��<����(�J�T��_�������!B���)?��q�}��-}�M.��\h ��T���Mj}Wx�T�@���g*2�����߃��-]T���*%%��z8��_6F��ԅ�\ۀ�\��eb�r�*��-�s6�AB�FA�!��6+gO�����ņ�P���ԛ~���2z�+�?>��C�Զ=r1�O�B1 s�,����Q�(���HM8*zb�~#�t�h ����]��U�xH�b6� k/#$C5 3��H�i��n��Lz�̭��@�o���伿-��iҽ���p�b�� �V��K@"��8_��VB%�^$�O����Ϸ]� �4S����Z���yo&�����d�Ũd�D��ln~D'W��}��/P}U��OQ��Bˑ��cN�_u#�<rc\��ԺnĆE]0��o��9Kߣ)y���I�%�V� 8<=��Ct.�/����������+�5�^�+�뫲��{+2K[RR�{~�\��yx��<���5����`�����(1���D�p��o�F��vYU�ffC�'J�����Σ�y�'iw��П���g��HE�Y��q8��8�`�I��gM�=bv�]Z:���yN8�B>��/�
�y3A��5���/7��6g�w�#j�Dlw� ~�u+(��k8����_��(��*���T�(
b�~�i"� �RU65����J��ؓ�čp�1x��sO���O*E�;V7��Y�gsrQ���`�~!�/7Cہo��Q�Ο0{8�ѕ�iڨ���(Iw(���X�!5\4�ێ��"�.��MJ��jđ"T
���͓�^�l�� L1�MY�a�ۗ�\vez��SA��?\<�rD�Y>�h�u��%�������}y��! ��R�����L���B"L�����(�WЀ�R�h��-L��b��yXO���"�D��֫�����=�Ƿ��Iq�|�"�1���ad۬a����A�eG���w�H�\:�&�ǐn��\�bEȜ����l�����[W��{`�Y�)^8�5.�#�h���?�q��p3, ��Wn:���8e}�#u��)���%Đ�����K:��`l����K��qٯ�S�FO&��
f9ZN�2r����W(�`��6<E�_��޴���odJ`ʤ꧀�a4��R�W��0�>4,�>�$l?:��Z��l�͵D]^��M�~�K�la9BH4Z5V�L�QaD�p�ҴH#J(^��w7���@X�n�xبٷC��n�ް���M'�`_ g_4�*V�c*�?�8%��������UC�ZmG�W��9�_�,��֞�*}�MGX�E-pt�@>!��q���l��(���{Ļ[����Qy�ڂՀ��D��7��~"�bȝc
:�g&]����P��?��;0�*W�2�촢K3���Y�/q7�f��p�k�ci�BC��Űw�m��El��Y_*x%��y>����(3'���I-ӕ�6�7��A��F�Ժ&���E@�	OygR#ff�^9���!��I��.�d*�c�44&O��ǽqX*b�o.���=�@b��[%�1i����ҥ�`nD��Wِ�	�S��Vm�j���Oܺ� F�5�j� }�x/��Љ������4)�������G��vP��V,����4��&7%��,�o��X�@bM�u�(��G޴�7�N������^s]e$��{av�l������0���v�M!v]�'���K�D#X?��3� \_�){d>�)�X���e#����0��қ�X�*����RL&%�.������ުE<��C2��û�fZ-��!�
c�Fqq������oZH��y��$|�Y�"��@��ΉХ/���E�L݋��B����0	'6��d�#��']N0g�j��D�����u�-�ԪNɫ$�K�멠�kr���b��jd�1=��e�R,��~��_Y�e�	ꪕ"
>���� )�y��:BX�Nm�&m�[lT�*� '��>.r����ypa-I�o�#'Wkj���?�ER	C̢P~*HE��ő�4����{�!�R�^�һ�p��x ��>���.�(�v#�b'j��e�gм�L�gEj�=�'�-F��]f������r/2���:l2Z+VZ_���	_�R�PGc.�ȼI�>^�S����	�dd0�簹���-�}:#C��2�^��0���(����+U�p<�?�f��,,zIKò�ȥ��p��ȣq��]�(��c69�1��z�V����q�0��4�V����^d:9�d���^�q��m ܵ�T�ߏ#���9v5^@�l���O����G&
,�,���Ϻ�h�S�!��ݔsȰ����F�M�;�쫯���Wy�����N6J�4�U;+כ�5D̐xvq;���js�0T�K� �X_$���~����w3�&_������m����Ͱ��("Z��M��эA*I7˭/��`|�+18̚r��6��5�_'P&�� �_���rE�7� �d�0�w�"����=D/_�z�#��JEu����Pu�R��u�#�&��ߵ⌣�[?�AG������\�QLR������z�q�i-��̶YM��n�j����?��-\��:���}�L��0L��T�<g�L��T@%RdWn�Ԋ�[�w3;@����P�\���n��=Q�CW����;��̸������%����/E��.#� _h�Y��Q@�D	I��������zH����7]�XqBБѢL�՗�1���1eYE��!m�o�B��	���h��醂b+lժ]�aB�J]Asl�`�i.|�|$j�'�P#�d}����i�(��Y�lHn)�+|�:!�����y ��FQ�-[U��z�8Q��6"�-(�d3�3���ם���m����o��|4��s7 ��<�bDI����ږ�0P��f�Iu�ߦ��]�cy %��/���ё�'�4P^R�ԑ���?]�^Ȁ'\ ѵ�R��ΐ!���y�9�7�(�Fm1���!;E���Zˠ�;�m��Đ\w�J�P����ۥ�/��0F��H���z��Z�(�P�k�+�Z�R!��|��"CԈ274�d�G��ԺzA�^Z�
�����YjZ���.�J����}���L�:���`�����S���1�
D���H�&�y�s���$1[�^nm�w��8�ݕ������ez�ej�|9��(�Ъ'����6��M���}�r2�
��ҡ��4��Dʋ�����i�L��IXЀP�=��2h/�G)z7�'C�/3�1-q,vz^�(��ŕ���޶�qx}�(��K��h��S������-@e�]�S�X�����5:�=b��ދI���$�,�y<\Z�0�ģQ �'^�A�,ҟ����\;7�26�9�g�@ۍ �8�8}��ø.�^\�&��5y�s�3�{��n��!����Ǖ�F� .XS(`a ���л�fl�嶜[_�I��������6(�|��W4-\*����y��_O���8��{<��Ϳ���BF�������mկ�h ����Qd�o-NwhF�G1D���pI���ƛ��c@�(�bc18��H�b6L᯴��r�Tp&	�G�ލ̖��5$t�畃����r�(�ٕ.��Bб�VG�K1�%HzRݣ�=���j�/�Z�4��O�6�& }�e�"��@{Xp�M���j��
D�G�.-�<EѯD\�&`���{~� y�؈3��߾����-*f
�3��#t)%h�h���2�Xe�1����O^����>���)�}z�N�\�˙�ɦ���u���u�� �60X1���%DUT� ~V�§�Ώ�������4A�R-�:�\5�����z늽�U�L�b�JR��z�cٗn9��\B�_m�S��&
aB���s��ܟލ*Y7��T����Z+ g[�Z^��g�����,Z�^��/�4}���2^DRm�+�ϴĵ����ы�u�K��%c���>ă�l��A*�0�Z]�!1Ŗ4k7%��3<�8ݧ�r�7��oe\G���35{��"�=���*���C �4�ɽ���-��D�����4qk"�I���'�i�u���Z4���q�Hi��qf|�r�;�$p�ҧW++I�u����:��m`�����SC;�Z;FA|�6��������L�MxӃ��Q�*�ż&)�
C�.Jt���Ż=*���I��El
��Ϸ�>U#��!�]�L�4z�Q��̧�^OCI+��8ʃ&�/;g��Tt������ѳ>��I�@V!����0>��:���A�w�\2%�`��5.ā�K�!��]$�z"�(!ZO���ݣط���:7Ͼz�>*eS���|���4�8���Y�?�](�F��6k6�~�:���jNL��u@Nr�k�^��e�z����X��F�6��ӂω;�*@�Ŕ�b}��	=�z )d�����@,���0Y�|�H9���<#Qp&�4U�݌�T�?1V�	C5���4w��$?M�$w��+�`���q�A�E���rτF�p�<��^�L.;r�=���P��UL'Ю�r*������:X��u��fl<��rjj��[�J�|�c F��}��V5���|�鼢�tC�#�Zp��*���E�<	l;X��z��ݾr��@4�%W0<�Ƨ�/!m��C+� �C�p�;�~�(�|���9�i۞9�E���J�ׇ�o��U��m��p�v��`�Œ�tMu��/ ӫ� �!�6�^F��5�2�c�vwLS�r���ϔ�?��='n��iU�U�Z��a%��Hz�<��E��(�D�;X�0Sy/#��+)��~�.>���	� ��#�3�B3�(����Zb9v$����4 9����4��@��7��^ws[�-9s�����%������-ʼ��(Ѫ���QO����=U0< }�J�Cq��N�K�Uk�P�e�
[�L���זe���v�X�3�xz��[
�k���Ý���O��T�:�A�2߳�d��x�/���J���_�Xg���Uq��)�K��;)����{��%N�Ġ��u]�$\���Vs<G�Jw��a��@l�+p�Ό5M8�.k�Ù�o���E'F�'��~C��Y{�꒩��h>{ ��z��~]!�`f�@���A2ڦcRd�!Teb�P5��&�Ye�U���F�G���#���!����a�/�hB��eI�)$0vc[=�=l��h,ힹ�W7��g�cL�q	?��_A2y~	��Du��J}A��_~�V���T���?�瀵϶�h�8�֝]�5bǒɘ�8|A�r��Xc�q,��+���S�I�=aR2f�_`�\M:A�ģkJ�T��<�#Y}��5>U�)�)��Y��
a�B��U����z�R���\�𡏮	Ç�fR��@� �o_R��y[{C���턏ņDR�fM0���9z>���+��@x�.� �@���C"�a�f9�
�
p)-���g�� m�6�K�C����H��㬉��^z��9���S�af��bh��ߖ�ʻR��V���Z!k�l���o�`�z�T4����{�H�[;�*�053��Co��Y4>���"�"�U�-�_�N�_Z
o���ێ�R�T�(͈?�������0�ӌ&	n�Z���_��$���|r'�	�"��rU�!��
.�I��_������qU��!y��C��ظ%fmhfǝJ �ѫ��J[�i,��}4��ҿӵu�Z�0"��<l���܄j�`��/�5¶�&KCr���p{3�> ���8ŀZ?��?t�#�a^��~�|�
g]D����� j ��#�s!�`њ��^����T:��ES^��mPQ/{���=�ό\c�$Mt#v�	���D��+����Ðyɒ����>�t��B]�+���*��Zjr*�I�U��f��3׿�{����Vպ���G�H���}���=C�=d:��ʋ�#���-ґ�g3��G��;\I����@3��>R"�o�B�:���a= ojy-�"�T����.�E�R}nAE�υT5�	�	�� ��1	ů4���q�|M��+Lk��w�=����|t�Ӥ�A���)�4�8GM�nh]?V�4@ ��!R_�BJ�P�*>��u�Z��$#aoE��G]�k�mNQ��m��֮µ�����ij�Jeb��]��׉ݔ��Nv�q��~�Mw �|�����HTR���mR;6�Ζ���Ǭ�V��� �~v�� �D��XE�FH;}�f@�J��b;���Z�8�����5 �_���;7��Q����w���p8�ÈG�]�/���L6��W�,�U�P��F���5��Պ�5��D� P�CMc���h����P��dmT�gܶe�D�v t_Uh�^�7���LL@�.?@7v�1,,�����3L���f����(D�F�l��ӥ��o@�d�7�Y�'P�l��2ZS�a�(uV�:�����C7��r)7aC�4�'x�?!�c���_�e�(;�ki�;/F�x�"�<�������Zn�E�V�w@Ayʮ�d*,V;,�2���O�E�.�@�|����q$R�56Xx<ӛ�пJ�JXdߊ�q#|�h�(1j(����ѓ�=�;t�����E��{p���s�:���&�`m,
Q����ڃ�����PU*oc�lh��ʌ����ȁ�fW:�$n;�4n=nt�E�.�nƒusw� z�ŋ-�	TBV��l8�u�%����n�$&)����0��&\B� eL����^��Ʃ������vR b� d'����Ɏؠ���b�z�f�/�~����,܎ր{��7�@`�<��h�G���11끶��[���{�`����3��_k�h�tՒwx}}��%�D9B�SlK�I(uǇ"�{��Eb:�ǫ��`�*�Ơ�M߁�����Lܶ�XM4��J���ݍ����BЁ��\b��=���P#��m�s�K�4)�wQ�W��/C%�T˩���d�Cn�ܦ�I��Plzi�R��נk4��"���X���>�<�Is�S�W4�-�Ш��c[���g�<��f�;�+d�c��2��i�}(9
%%��|��2HĹ��b��~8c�.��P���<�65�7�����2�q�`��C[��3����t�@2;�Karxpc�@V�J�Lze�bSm|�*\�Hyڂz����]�  �O�8ȐK�������*Ϝ} *$*8'I�,"M*@=�G}
l:s={�Eq���:�Ԍ�%�R��2�(�uz&�x	fV�b���ʟ{��'�պow�{�gL��>��ιTpF|=F>G���K�
�5](vD�^��2W���Ze�)iy��b���?��G��8Ô���Ҥ�p�H5���7�G����ٲU����g���2�d�*�֥��⥙��P@|��s=
�M�z�)�9!�@�2�z���yK�H�x�W1iD���u~u ���e�,m�5*�bϨ�Lx��a�M3eNv��m��\�x�-�؟b���� T����Q��jԦ��l]q?�x���[��R��V�߃%�&N��:��֋��7�y��Vێ�?�t�ԡ��}�Ћ�� 
���x�X������a�� �J&�K�-�4�4� ?�N��>��`�\�N�3�M7�VՒm��_�g1�iB�7�kK��}��?�J�+*���^�+��a��0�a4?�8c\�M�W���X���F�e2E7eYLxJ�Hr1J�ԩ{��,M\�:'_"�e^���a���I3��~�_/��ro�72�y��d84��<��d&xbh���\�`[���7+]s�t�ُFr΅��䮈��6�8�>�;�C�?0���}M٤A�":|d�F y���}��Z�q��{����N�U'�k߽���SQ\H@r��(6|tW�����>��!�
�0�[�[��EY����V:zE[��RO��Z��I60/I��>��Ϗ��肟���Cg�����lD�K��WTcUP��c�&E��G+��G�|��
ԙT7ԋ�)��_F�,������B�"��W��j�嚋��v�5�����~��x��}b��ih�?�y=�eܷX�h�o���\� �����?Z� ��x��Ԁ�v
�e'���o:"w�x��1G�f���T��9T>���o�v&o8@����!�H�g�5\V�!���B5��m埁���"7�{�d��W:� �(9j��"� ��eʨUh��[�@K%�D���T���/�\>�7̏k����s갊�i����n/R(j�X�X�8.Q�X.�Vid(w7%Jl�S*� ��\*qX�5���F�r�}/`��ԁ��c�@��!��D��G+9\�eWP�L���h59�m�|�ȮZ���t��5.գn��.��lUQ��'9�dc�m={mר�H�{i�s6���3�#.?�=�W��e��?:u�at��ȢO���}�"���i����4F�������M�
�-ݬP��M2�m^�L�U��j��KL"Cx>	C��6 �ޡ��Vg�P����1��嗯���Lלѝ��0L$1��y�����o�Ղ��lbo���eaW�2�؋�����7�MF KC��bE��a��`��ó�7�*�����v�qq`�Ȩ+�u��M��m��b�����X�S�`rv��<f�^x0������ ���ʕ�KƊG���!/w���8��+�s�#��˫�ie7��'G�?����oF)_��)p�����S�Lt�T�s�tRA��M�!4�!����֖�i,\R�� ieb~��pq�?�ј��^"������>��g�)����<�C����9w�&Q��Ok����[Ǒ�S���R�݉�3_�'�m+H[Qه`���q���E�i�V�g�g�g5;���5[�t^�jn��ϥ4���]!�0�e�\��8ߔ/�ߞe`o���������Hi��e�!	eG��Y�}�^��l�ᜩ����ua�B���mF_�*A�����	k?�c?]�:�2��G%���*�q�Ώuv��Te�M5�u�h�:lq���QP�ֱ�bG�2�@hSE3������K��Y�趽��u��z��Q�\��ӱ��L�g����ҕƜ��ۍ�:L�q0rɄo!���[x�W��+ߦ)�ޭ���KR Kz�@F���e�Y�!>���N��;�LOKO[����\�
G���\ص�>t}m�4�i<��谮��X�
���v�oEÓ�}���'�	� K
�'r=��<��!eHBQ�b�y�Y[2L��}��%�(-Vt7�1T�G����&�g\��̆�o�.�j���Y�ߠ,������_�LJw��(G����dp�<W�"n6�D� ���JK�Ez����%�6Kν{��Ql�qȻ\{�r�T�Q��|k_16C\��b�MY*�ҜԂ٘fޓ^Ȼ7�d����iH(��C{t���'�$��ۅ-�(��\����pJ>'_�o!��^Nǘ����z�gHS�&�~OE>&�0�t��mp,[*D?f)�:L焢��ܺ�E4�������5E��a�/a��.�c'�_�|T�'$�E	��Wc�ʄ�Dv��O��I�T�e�d�����M�H����E��&뗯�yp߅ovr6�`�t2@��{s&J��l��C��b!G�F�k�֔si_G�%�n�vh�6��=�����MN�T%2[3���`����Ԃ�װ����DZ�`�4��O-ZF��&��t��2�P�jʒ/�&uKƃ���f-A�nH�.������v3��\6� ��Ъ�\�q����D��<'m����#���q�LqMnN�9����R�Z��pde	��욿 ���vo[/we�k�!��Yu������U��A�͔+9΂�	�����!����I���jg���:��W���4���+K�[�qٗjţ�
(��f*a��������q�J�X!� ��,g�k��2������X�ݷ�M[�.g������ k)�7�A�n���<��6:;���_K��Ք���i�tP���S�f�R؍���@��M�%�8sƯP1��?6!*>�_�h����/
�(������G<�S���Y��y�5�mW����sE��(���|
�((��I��v��X#�
�����m�7-���q�)q\*"��[Է�͗f����40J�/~0��t��-1	6��u���_z���i�.�>��c�nh�~��,]f�5�q�t�š�_��$��#�}ʅ�p�,�>��U Տir+[����9����T���}��#?�*�e�	���mi�H]�P������7��J�,��H�q�1�8�m�l�6 #-̈́a�� �6���N����������.g��'���1,���LH}���bd���t��� �öeV�K�B���4�
}��xT��Q'��#Cn���	Hh������޼�-�%�P�W�^@-�(����������KJ��o+���$it�hII������B�:�aX�e�:�}��ƈ���A��J������l�l�v̌����&�Q���l������&�ҺkB��}J���Մ�)���h��7�T�(�k�&��hf���k�U�u�G�3�.k،�%a0i�h����?kS2�z�tMW�Q��ؚ����G�&o�/&䗥;�]���I�=����/����,+���R�?�NJ�r�3��l�)��P+EО/<��C!som���`��'��ŉ5*��?5�U�I\4p��V�Q1
�PJ����/6�������]�Jį�vq�t���h� ��RPv��݂�:_�4ϔh��jhpѠ)����-�w���$� 6|�q���W+�ȣ�\��L`�(��"�`3%��K�}L�I�-.9T ���tT�Y�������ߋHd�E67Y��|��{.m���%J�1��#Z���v���Mb<,\V��G�&SY�pMo�B
��.��<���@bH��k�D|�D�o~�C̎�t ������7K�)��Y��0B �T��> -��%ם�h�!��R��TS�N\�Am��U�:�:��R� 4DK�LH��rf��L�o$<��p��f������#R��*[j�X�?�S�vn7��-%F�)!gwp��ۜG-���&+�X��4����#���*��{��\֒���J@I6�n��Z�#����gr���G<�{��Մ>7�$d8j�O}���	
�_�S>c٣��&� ,�|����۱����*��6鞑��7�G��[0�9ͭ�1�:Up�_9��D�݄^��OW�%9�N��+ָD���������:d�����p�qvBJY��f�C���^8Mc ��U���><��p���{���/,˜����*�V!��] �g:�=�dQ�?��d�۾�n�_ٚtL�zԤ�1�U�ʱdD�!��د
�([uH|i8]#��iAyH�	'���)A���]��X��ⶂ_�\| UP3��(F��x� B�J��@`DF̸��5z�!�:`�dc���a�Y�'�%�3E��Κ�5�F�A�e! C�zx� �=��RP���0[ᲊC�=ZA�E�(󡮔�Z��%e�u0֎�G��O��Nm����;��C���a�6���� �7]�V�������D�=a�|���p_��YQ�ys(��/#��ܒ�5?��.A��XV�_'�da��7W7[��A�m/��������A��6�2�^��.��y�R�W�望�:&��h��%���~��#,&��f���Ȫa��ۡ@�HP��I��$g�O׋g�g�uRO�Li�S7�Fh�+������I�� z+YY>�]p �����bh��{��4�w]�
� �s.�ީIR'���+R�+Ȧ��!z��S�]�{[_���kUsM�69�:�*�ٜC5�P�.�ٲm���V:$.E��I4�b~�>|�PŇ���>�鈷�p:`ME<,Vō�^K�^�2`���-�\v�Z��ٔ�7r�7(+l�t��y6b�u@�����Qj��;��c�/�����c���7��@�p�Bv���wG�Y�Y��G�vg#�"����-�:�6������9&LA6�%+���������#i�B��-}N j|��]�̷_�s��ن�hY��2;`KXM���ja�
Y������}��~�A�����N�@9M��Դ!}߃y<��|Ü�P|�b����{���\	H���e��ߟ)�:
�Ƚŷʾ��}�nH�Ul;V��'LQ/�T�g��W�,޵p��(e(��M���MzX�Ԝ��cş5&�Y�hI�>���v�[���?/�?�+�'�U�x�9Lv۹�?=i		�v����%�Ig׿6�S1^��,�����:�����/6�Q��Ġ��hY1�a��Q2Ț���N�i
���	�˫���4���r�:� ���H��ɀ��V�)B{Â���A�A*�yU#Wީ����`9��ư)��Uy�/nD�t-���	�lT|JX�H�A5O!��T�}�4�3Z�`�e�����	R�� Ab��J,�o�ꇂO/O��*$����v�!�FC'Rk���KOi������\4�|�~��zk���K�`W�� Ie�IS@���<�چ���~
�'�Ɇ�U���u�g/��1���+`�֜&�o�n ���c�X:��Ԓ���/�^=�9�� �g��=��?)rqW�#��a*1s�!AK��@TIʷ�:	�����U<9��:f��4�_�f��Z%Y{���U�:>˩[��^���ğ`
���%�:�Q��bed� ,�40�Hњ��Xd[Sg�<#o��ۗ��Vm��u戀��:`k�!��+Y�3.�Ey�JO�4N�уvwG̳>S�ғ��a��#
}c����q�w���+��Ձ䤁)?�EEC�|`(��D���ܫ���8�5c��@�/!6ZEτ!��-9��=py�+���L���pmE����W�k����ce�Z���&�N�W�t8U�/=��2,L{���O(�zn������qX����Y���Ȱ�Z�L��Y��+�3q �ܦ�j�-[�
�3�ڒs�
`g�?�Hʯ#��Q�#O���Q#p�e
��E-}k6��~i��s�]K�޶�R1yH�Ŷ�gx�rM�z��+	��X�⺤�{�!ޟ�� ����6!a�k����ٜ��74h��[q81tb-Ͼؕ�5��{TU�ie����Qe+���G�ܖߚ
��]��?�
Zp�$|&Z�G;޿R��o�=�3td���j�@��e֢�u 5�@���I4Ҡ�IYj�g��f�ؾ<�b���i{d	��ڃ�B������;80�2��q��I�-&��}9���z�=�Y`T4�A��U�h�[1T��͎���-�c�}�#^H�|����|]�\�9>��J1�*�u�����F���_�-	��}��d��F-�iN��$�W���v��1,���pY�Wh�9in��Y�M�!��K�ҧ�-<��&�/bXFj�1���T�l=�z�a�Bl�wA�4:(f����,�(�ǎ/ y�W�8"g�-j�c�> �]�w]�*����gI�r(gV0 ����-yX�؜"\ڹ��Z��j�S�*��۪t�I��O8vs.����<]ˮ��ǜ���Zl�Rٮ�1#\y_�O�
yGM�^��{<9uNt�
C�iP�H�u��Ka�;H7+�$+�rR>�?jU������<X���E݅6���l�$�:t_R��"K�v���H�e��/�~�ϙ�=��ݼ��*	�x��7悲��S0�"����G�.<hR���Ʋ�`'���*
�I�r�xf�ؼ2dJ�'�sT�7�t���S�1�/1�T�,���g�~^4v�6\ �ӻdP�W}��Cp�tw0fr�����;�?ϡ�'�1�{4=R��"]c�z溜^���S�h&^#���N��%���椓ʈ�|�n�aZ�\o�A���������C��$���o�_8fÆ��zz���Eh��� ��tS�D� 1u�j��r%�̠��`�Bi*�h�x2��#���k㢶�P��N���8*�ph�j����t��+�)t�׀�#1sǎ�&�2������%�B�w����[L�&��c�ռ��Ab��f���j��(%�����Ԉr��^z�dHw*E�t�BK�l��<M$�@���B�.�e*�k�-�A�[�5Ct��~��9
�g�����*�0e|��9�',}"���F���0��͎�?��W@����:C�د`�}�k&�
�#�9�ϓ&�N�SA�WXP����=����{�s���jg�js`�#�4����Lr,�������v��mt%R��*-.�!��d�i�nd=�*.����+3
��L�x���+|;�'tc�%��B�۴�wLmu��W���l��a�����P�|'�R��Ӛkֽ�D�_;���-���mI��ʬZ�j�'S�"��~�ga�@NO@ςZ�z��P�]d;I��{����Ό(��bu�\�?�.8�l|l[^+Z�i�^�����e�#H��F����oq�!�0[��!h�o�i3�?�G����k
B��ޭ����H�dH$�f��h`�}��:q�������"��)��	����q��4@4x�:EL�|7:=(����oP_�L�q�ݺ9�W�������:�e���7��3�����y#-rΕ �aU�!3�����Ha�F��T�T��C�ݼ1H�Q�h}���BX`4��[�5��j>�&���Vn�{�>���P/	�~&��h2g������̮���C��,��X��ʓJ �d�mbB��nks^���*�b��'RIz/��8���Uj\ֳ_�߱�T�f�3�b�)��\�dI(n+Ez#s-�?�%���5��]����V�D4G�<r] ^�>��om�5�L��Qh�Xm����[�9ܒ��^�K����QS�k�6P�?�����ep#1�#
��W6�E֥�7�qT�v��dKN�[��fb�B��L�w�U`s`��:���D�:��'�h?�3]��ɡQEP�.����O	�e ���.�O��>�=m����1��Jz��BTH�ŋP05P@^�>Z8$��H髥�}I�c��8~��\݉%2²p��_�ʹF '���`D��l���ZK��+Gn��ˁ�>]��RE�Zk_Ȅ�R�n��|�m�K�ܪ��$o�d�ȵ{�qL��+/��aJ�ěvxX?'�!oe�NB\��Q� F�'��"�}WGc� �;n��e�_OJn7��:�S_tuI�fH� ������^�h���ل2	eht�2W8|N%<xJ���0en�Cc�i���૔��4U^�l[>A��uj��=L���1�S�F/6���Ҟ�A\��������-?�}�,�������<�����6�� {�ߨ�Kjٸ"S�vD�$Q�M�&5���V��cN+�J9[ė� ·���7��"h�i�*����򦞸��W��N��A#�ķ�p�FSzo��7�;�z��&�\%�������TbF��ǻھV�`��^�Ʊ��`jmo�gT�꾨G���?�ȼ�8���;�Gd��X�J/<�G�3I�W�`���)���T�

8��D��F�{���}������ˡ�F�Ӥ.�16	/�N�J��M=��g�k9��㠐 �Y?|'�O��Zwft��6�Z�ιDZv������a4�����Ot���jWێ����BA���,2{�g-���*M���nOA�n.��3裠m�]�(^U��`���'��Q}�X0�?;{����XA#����B�%�������»H7߶�J����9��Z�bh̡,$]��8�"&��4X��?K)l���Gƽ����~����튖�X�S?� �唨���E40+��c��R��� ��l���-#	(?'Pc!�s�=������(T��ꆠ��l��z���Al�Ʋ��}���%*�&��](�j�,��u4o	V�J���<s�4��K��4�	�e�^tSg�a��.>����*W��Ǯ����L�',Ame��E��(�l*pQ ���P[�i�w�~��k�����1�;�\'r�]�V.iOP��y� e^G-�bY��G{���dj����K8L>��y�6W^����N6���T䑝��K�N.�&����/FB�e����C���_jo����6�i��?w5����I�݈�_FHh b��vd����2��-���8�p��PZ�v5 ��TQ8��ۊUkx�\����!�G����̴ty4��;���v@*ʶ��'ܵu0�ڸ�p�<�g�����4�w(6�8ZK���'s����Ή�r�8�p��u���)��?��}r���c;���L�� �G�ip�Q�ĭ3�a�:4I(�r%��D����U>���r�Oİ���L�����b�����I�\O��g�]��G��$:�vG��ad��Y �Xb'��lV�����gKD�Y1T'ׯ]ck���E���/=�v�.&f�{�
�n�^�ʣ�Q�\'G'�u9��	΂����w�?���_��G�Li ̈�H������O[uΧ�o�.�����yjY���a#%O�W��}s�ۺ+^�G�Q�Yh�]�UxD�� w�N�8t�D����Jc�!�.�(��\�2�x/����W�ݡ��3Iy���H�V���������*Q1:H������쾿�jLE z�����b���Œ��T+�Ҧ/ ��s�!ރn%W�{��S��y�
�=�;g�xr��p����G�
�a�ɺ\5��j]��R9rY8�@�t�]��?���dY_��m�oj�,(t	���y���xcL��\�aE�o���5%Ly2��0������������Hd5����ҏ/b@;���~�?9�4Z��lYPW�*m��m%�:��Du*�0Ic<��ؠV�CE`���]x��rpa������+G,i�yp~	!g �I�{w�L���q���D�i�4��ʕ���A��R�~����tڴ 5���w�8>�O�A 5���F���^��x�d/I�zE�Ek��P	Κ<T�D��U�½j��/��| 7otL{f3Ų��M8E�!�7�ŧq�l�C���j�+�����_�ZH��q��F+�lB}F���:�嘺�G#
�߸��o����"R#��`J��;i�ӆEGS�R-ʔ�;FA�ˢl��A����a��f�^~������U�h�I�ek횸ܵ���#���r�ҽ_�f����,�9�#�\�	ׇ�{v�՗F���.��YMFo�S)���t�H��$�+����	�#oO�2�.B4eq��\1uώ�}��6\%ب�6��Uu��g����$�?A�_1ܐ�-�4�O
o���_���]���Eȷ�P�Q�C2Z����.�t�eqͫ�1�I#/|w�fK���>����D��*��I��X�)�US�)K�HI���8/1^��6�uZ��24z�[uf%m1\n�t�s���]���c�;$�B>X���O���4�0�5j�P�;Pf3���J�ę��-�Gǝ%�Mo������4��Q����"JqAJ����@�M�>���n͙��|��:��:Q�"Yy��O�m�.!�#�qPWɍ~&�v�Ҕ���x,X@:z����W�>{$��4����᪝��u:�N8�$ 0W��p�ԬԉF.D3�gB�Q��z��bEL��F���:�Q�,nx�?B}��x�W[�zi9Y�U��L��ӊ}`���P���[(�N4>&P�X����9 G}��cy#3z��&��� P?���T�j,w��Q�]%� Y@X�u������K����.��Y!��f���6�����k�}uU���g=&�^�:�Ͳ��<Ke�<"����U]� U7ڄ�| �G6��i�>U4r���ջ�D!U3�5Ӈ�Z8���5)mjx�>"�@�x��p�D�g�v@�5��\���JD�T~��y����w�s'
[�&,I(��渗H������yR�bG9(��b3��:���C�i��zy��m
#֜���se�Ճz�Ax͈�;�,�s�|�v�2�j4pzqJ�:#^P�zn�\��.��X��qD��	��0δ�Q1�$�
�O��!.�s+N��B��ˉ0�+w��/C���X缶ٯ��|���)*s{�S���i\����N<�K�����S�+�M0Z/	Ûy�����)%`7�i�J\�Hd�¬&+����nbF������I���>� ^�F����ߧ���%�.4�h��9�$�Jg,�b��~_��0Lj�J>�i3���I���/y�v��Y�#�"�p�_(�_J>��q��/�'=�I!ZeL��X��х�
l[�z�V�AA�����>��.��UM=�9d�~%�Z*U�
�H�C8y�/�&W���7U T�>g=�.������;���n;�����(z��ǽ"��ͩ�r��Z�rΑ����*�%O��o� ���#��y�1���ZG�Q���Ie,����vjM�z� ؉m�n��]7��I?����-�)�w��|�+f���V��E��~4W��ji�9����x���[���)�=�(|�do���hkd �=�~Zݬ���S�$��o6`T�R�R�A�:� ׽	[��0������fw�&��
</I7r�lE��x��p��"�U����2;T����n͓
݈o��I!i�di��*�o�A�o�.�{5��5�\�!�?�hj���s  ��j��A�7�t�Ks�����i��O
�^��ʋ�6�c[�\��d�z�sө�3�)lp]Y�~{M�A� t������;ڱ+�4+�#�(r�,�{�BHS�V����0�|K�a�)��l��V�
��7��R�C����؀���]����a�0�L�k��K36~`����� 3L��TL���2����x'+�Ď�C��������T[�_�b'E��
��퉺�p�����ݜ������@UI�с
H����V��	�O����k�|mI�tV�Y0��w����j��^�t��OJs5��<>-?RD���B��\r7
|Lf��JMj��薧U���6֜0�z ��$�T���X�UZ`ou5�6{C�5<�mt�4�`̛�^�G���Wf0!)�����zM�0���jYr�|�̣b%�ɀ_��Z��b�u6(TAN�_(�[CO��,�k��ͧۂ� `ֹ�����{/S�<�a�R��m�;�i(�Yto�I��;�܇����Vb�#zϥ;���VJ���N�:~g��(E\��޸o�%q�z��,��e��MC�q�Z�@sR��XOڀXZ�Z���xȿ��m�-N���q'˞��۬#�q+I�*_Ψ��#D�PǚO �;\��N�C�.+�\9�ʾO�iG�舁�r�y�r�����> Kk>t{?���c�B2�>Y���P�/@�L�7�4霫�
CCx|>m�wM�Uz�'�w���� ��<�5�`�a�u+�t.�$��׿���t2Z����s{j�_�o�v��?�Z�H٘�I���\����iw�%N���J��I�/�c��q��>)������l3]i���{V|�H�:�S��>>'�rR���&�gY] 5�x[�����
�Hno,tb�iW:^hf%��=S5�/au8F�P��2�O@x,@:j'��N1.��bj�N=C�x�(f����6�m g'[Z�~A�\�iV� +i��tԁD·O�ݱC��FM���1�-~��$�y����k	ӳmC�d7)7b����,�*�6s�/�Y��og�{sz�7�}��>;l0��������-F�=
/���ܞ�䬘���N�� _={�=��
}3��q��+���mʸF&˘�)�%i�[���8�_fA�<��N��5��퐝GƋ{tZ@�ה��n���!�@�&s��=<�6Mƌ?n�ZNy�w-J��a�9b�5:�a���u�NV{�H>��ePV�w�=զ�D��laZ^Qv�{ٖe�ь1"�u�&�r �\�Uv�?Q�\�V`�dȘ�j�p���w�"GgcE�i�S#I#���UU�����N������cCGB8�i	���(:���B^�ݎ? C���K�ֆ�L���-F�����Xt����Q��ω2Xa]�I�踡�쨣�ɩ|�?��x0r-�E�#l8��l�|p�Q\��>��ۖ�g��:2�׷K��XGW� Mw��S�:��R���������&�����hx��+�����f���(Q�&�E�^�LE��>����<�1�!'����
y�uP#Ǡ���W�H�,j^8��1ݾV��9rs?�����&qsH-�z|N���a֐� ��
��v� ��Sz5L+_}g���0��Ќj��]*?#-$'R���)}�p�5���3�~���d��HmL�0����u�-ё���U%�����5���媘B�I�7��>�G�m�O�@�|�&	�����ӝ��%���H��ʀY����SISQ��=�v��<rN�|�M���Id� U�t�Q��čS��/Vw\�m㢻)i���:�O�h��Y��v=�F���� ���պ������(9��Nys�CfZ_K��8��]z�����T`�5k�a�q�Ҳ�*^i�Q:����)~t���I�����}���q��h�f���h>����M_-�xb��-�h#a�D�;,��n��z��Mr��=�.j{�ȶQ����m�����t�n<!����($�+y#2cv���N
)�|��Dt�� g�"�E�ل�4�Гj�|M��%	|-IR�U���C�9��ݻ�r�#��#o��h�b}�b����{z�'W�>W(�~W����V�t�����_�l��[�L�Ŀ7��޸�L�����,��[��G��]��n�A�Y�iM��h�Z��8��kz�ك}"��	:4ZU���\W@��<��p���F��ߖ����`��Y t���k98����?�#��޺�+�n}�٧B���O]���*��zpx*f%��gY��.G�y��9���jhG%�(�tq��IA�XN"	X�!������I�B:ħ{�^����¸��47��tEB�����Z�~ù"���G�s�5��)�)2�5K�r�k׍+�+v��Ób��C���d����Nv�	9��c'2yh/=�fU��ڰ6*�@��j�C&=7��
{�C2�<���,y��;g�O�oy�}a'ۙ^�H#wQ����	���Q��9R����ũɁ��߆�#�� u��\��.��8�U�	i�����&x��&���������k� ���D�~$J'�jw�d��HBE%�Ҧh���ơ����`��n �@��1�0^�/��?��=h�&8&'�ج���}�9��ݻ	9��D%��+'����C�y>��[����@�Z�Q���l�a�᠊�N��a�����Ϗ4�X�I;s1J!����E�h�q6�E���N�q4m��.P+��L'����L�����yDo�
۷��*��{�ͺ���~������o+�m���O:$9'�,~�Z��Q��C��O`y����~�!�þ�t�B?!MA�G�  d��u���f��re<\�1�>��N�yn� [hN���6d�Ĳ碠�$��Gi����p�&�`(��Fu��~�I^u�щ�9fk'S�9��װ��}�.�l��������8#������K�ρ��/�5�������ؠL�E�[�=h�Ŕ�"8=Ţn��P�}��z,'�P�IUR�b)zu�Aр�-��\�8 �')t�A�e
$Σ��mU\h��JT����/v����Ⱎo9.�W]K$�Z��0���#��`D�0�w�u�c�05lab�q�DP�E��İ�t�x�0'sޑ��0��N�<�6��R��u�FeN�^�O�ψ�(G'�D`U��v?���������F ʁz��ɠ�������=2M��!��~��]x�TJAm��
ֽ�y�e^d��:�	�"�m�,���N�_�6M��J#X
j�:&�o0�]^�����Z�|L�t�gN(^ �Q]o;���Ǡ�#:@/��@ �К�������}_�}НMI|�����P�9�4���q�_Ѿ \mey��&�yVn���]t�{PS1�.��,�O�_9/S?AK�쵦GH��j������Ct��E�M����Uj���*<~�/]�4�j���:��$�Z����;���bN���PYC&��{&��M=Ӟ��r-x�`j���++��Eۼ�U�Ug!u�Ѫ��_������A�aF.0n���M��g��U���S���O� �7�qP������2���!�c�����@��ҧ-��Gfw�-���s޸�����R�H@��"��Rm�w|2A��{�b�i�m�n(!���H����,
��	���9��k��B9��+.�?���%e8�&��t�J��'��^֗�T�������O`�v��q����Z�S:��ʔ�%��q�w~�f:�	(U������������9��y�ѽ��E���� '�q6��[�Wi s�"�s��a�# �D�,(C�ݞ��D�)������.��
U$���RPk��޷�,��-���������c�u9�ٝ�k��"4���F����g�ޣX?� D�K�/J���-Q�D�Z
�*(I3�.#�
6?ބ��\�?绞)��p6(�q6�/���6�疸���{�t�x=�]RP�$�*�?���[0��Y�W�����0���&�p������Ȳ��k�B>���x=V
�4�A�w�9��l����ݥ$�t[/s�񱕄� g����m�աF<M�w�V�4�eȢ��3�XO-���-�p�M=�s���U�#���}lg.�Bˢ�o�6�G.񂩗��-�L�Ez�]vf�6��֝�H�,v�iN�E];�{^��~W"YJ��A��lY��"��	��e�CO��#�)D�C���TZ�9P�.��t�.ڗ҅�(NKM���R�LIo�<1�H(�F����#�G+�]�]"��n5_m+m�[�� �t�s��NwyM b���c\[`�������݇j�Zl��d�L��/-���e`�a�3<�bm�8(�C��5�o�Om����������V�����魨*Kv�Q�����8~���?��:�3^&2zS��}��G1f(L�O$y^��EɑY�.1̴�Ƈg�=��UF%I����%c����Z/�v�!�eH��,+It�b���d��3��5e��ɵ��~ԉi�LH�U���h�zn6)�/�ßW`{�ɡg�\�bQQ�b�8_�fg�{w�sI/]�Gֶ���Eƿ"q.���w�s������sp����^�/|A�����	^*��G�֢T�vw5j��󰃇��@o�.UHE�<�,�H)��-���s�6�pc%�p�u�N
O�E�T5���=%�+Zܤ?E��.H�0���i��0�rk>�c5�e ���5E������&���"v�����gs
�����l.��%� *�\^�9f�a��G�v�Ǵ����PN���э(�a*W��c��@�8��;�O��+8�u��h<-����6���<��q�N��L���`�رD!Ԋk�@B���+ٲ_�
K�j��=h�q!]�.i��o��	\����Q���9<���@���L�<axp�qAn���H(�Gd|Pd$�j�L�z��������!�DP�KriO�1�N��c}4f���jr�yc��?S�1��s�"r����_2��!\n��/��C��yIeT7�ġI�=����cNA�g��3��C>�4���:>�Q����cUl���DӼ�Ù?D���7S�V7�A����4W��Y�?Vl�ɏ�g��;�P{��8�E��2H2?���Y\Y�i�I�_{$�
bM���*�qɳ^��^ƨ������E�maA�4C��j­y[�4"�P8$�H��/h��r:�9����t�֘��p�!!L5��6���4-�q	�ꆐ6��^E������b��� 5�j	�m�<�r�Y.*}�D�`� *��6��������{��)�9�D~�Z�$[�:��{��֑��i� �1 ��cAr?��|'��x�Ӥvڤ7[��`�'{���хÇ ��ؤyqqH2p`���9��P���N��>7�������.[��p�,4̝��B�|�KY"P��)\�_t�r�U��Xv�NJ�Wȅ1&�$�%.0�c��o#)���
p!ěi�f�T��%�8��������'~*��>`����[�O�A���ζ8�(�8��E�T�����a2�Æ ͒|%=�߱> ��2�o(�������dC�Ų�	�9Q˓>� �׭-Mv�@V�q ����J�vRA����h{O
�c�(��=.c%����
ԯR�a��dF}	�K�Q�5q��>��w�gKV�5��xȯׁ/��X��[94��*̶�&���M=T�O��8iV��0���`���B�s| �,˼c�{�x���v�6�rpC����80����Q8�¼���gh!$����qT.�D�L �h/�$���w���Z�(�:7�lO�Y��2��1��]��c�(��F��ʰ~l��������'E�$oH�/F�ȸ_ؽ�����Y<0���$�^������-d�6t�$�~�I��׀DD��v͜�<�P4j[���aA���mlQ3&�ǅ�x°'@�O8n�G����6�q�i�O���B��7�A�y�	��-���8
�,c�����2��w��y;9��cGf��E���4�ذ�̙�X}~���;���<�!��gw1e}�	s����"|������<ț� @�?J��+�ኲ�iWr��Ҭ����S���(�[�j�����m_�Zl&�lw���V�2f�k�]Sl|ˈ�"�8�W�8wR��-����{k�'�ȧ���_`��W\�����G��5��WB2_��>2��9/�'Z{]$��t>z�_Zm_氩+Ÿ�FW��zM�[Sܹ���k���w?�Z���ܘ~��ф@j�^m�����_������:�	[#ۺ�M�9<���#c1��(�g��ǫ��3v�� mnO��6�9a����b��fd�v`T���g F|�����w����2֣"��J�YI=�?�uD�*��y��jW��c�
[�|���x
����ɾ�\A�ߵyZ�`��x��+��.4�y��D�dez������^�w�Z�:/�`i� �v�+�w���Q6�Ђ�&�&��f���XU��b��&�m�M,�)���upk�t�)4�\k�T�Z�D+�B�<>�5�]𧐌XM?~��<~ͷiUMP�4���c�B�iӝ4XڭEKs��w��px�r��n�V�T4�c�Y,��QR~�ȼ(�'[��B���⶟l��������P+mP'4��ʓ��3��_�͏:}=Pe�W��:E��i�K�|s���å2��e&��ZP�L�G��E�u��/V�P��(���ƤӮ�5�X*V0���v��kؤ������y�-���.��*򰼲�7j'��y~amz��Thb%���?�A��9��.J��@BP?B��/Ff�<c��:;� N�g�ˇ������_f���V�H&�� �h$�z_�yd7��7�����M�A[����D��d��ׄG&�O&��5wv&��`]���o��9�I�� o�=y+���/�Q�dI��U��|�{X���cX��j�c�,1�EM:B��(:�F�v���}NL�,h9���p��L�9I��e��Pg�y���C��|72�A��0���3���ZT�Kɂ�5��#�?�����0���Y�S|�������LHGd�L����vp��"�X:�Lȓ���?�8����_4�t|��v��Ou1(�
ΐb�a��:���t6H�)�%��FT'g)�Zq���l%g��!u/����?]@�ћE$���jf� n��fy�$+���c��`M���O�ŧJ�7~��t��}�lhR�g����Fxaٷߴn��*�U�Ķ���bD���5j�# h/E�C(��m�rd��gE�X���/��ژ����{LJ;
�8�Qߤ>��C��Y'4�g�A(��'[�䛁��4ԃ�Q���6�a ��p%	t�sN���No'���NtPEf����D�����]��l�)>�nY�TS�1YBݻ>�C�B���u.P�$�2��8�A\���{�O~J��>��4
?AteMde��u��D��b���V��Q'�P� a�g{��m�:#��l�u���cظ/� ��=� �v��x��w)��������[\���q�v�C�N�y�v�O��z,���{I)��0��z<
�9���Dh���1���cB��W�ز�'O�l�q�)�n��C_��~��S>߅�}SM�A"o�It^����(
C,�7����e69�!���ݝj3�Ҏu�dw����ss����.�]��@c�L��=`�G���sO���� 8L�ޠz���Rݣ����WpKa��ZMW@�5�^�N��"�����֋u6�N��L�j9h	�;n'N<b�n���t=�q�Ba{�t���$ӣ����돜�l}"�m��t����dU\���9_��|�ۀ9�:t�B��${��a�]S�O��(�K�>�U�P���$�*Κ������иz٦�p���n�X����Iw�����}��u0�|o�e#��<-��Y�'O����:8�8�"��Tg���;����U(�)�qbz���ʭ��|�E�8{�J��U���)�=Z�6���E��������F�M'�r�w2C(v�
��&�^,7�\�}]c��f�ceq��y�MӉ���
5��H�	\�������g	�F�}>�����)���g.^�:>]��!�>e�hoԣt�7�`@o(���ʻ��3Bi�lN�ߺ2����q��[݅h	Xd�G�}�بD�4�W���A?ln,��O�M��(Q`5
P��	��F����x�
$9VYy*C4o˙n��s3�����$�Z;o��s敲��}[Y� �>�_�}klx0r�]��CӨ��Ͷ�!9�+aS��p��Q"<�,zQI��������X���?/�e�5����5��� �/��o�o�owS<e�8}��^Z�Z�#������ׄfX
;�/��?�]a\i�ߠuv}*V"r��b��k�o"�A�:�	B.�������{l�.�����Ұ�ӴU���y�toH;˫=`�!PsL�=��G�ߡ���5E^3SR�����U_��ą���掃߬�m�=t��Ã���z�8F�����O5v�g��g*pf�ݷv�SYmCm$N��V�R��x�R,�\�# ]��&t�Wc�<��}!�Զ�T��'0�+�Y��'�o�V��ᯂ��X�ݐϟ!�t��zysb���I�?�����l]u���CHW�#k�-����[���s��>b�R0��&�*�ąyaT���9y�t�1��1!��3�Bz�]t�,f���Q�ŵK��9%=Eo�r'P#�7�P������3�(dL{��]�]U�H7�h��šk~@t\��AZ��Q�['���g�s1��zVpşGy��,1.=
�'#S�� �@��Ń�~����5�c�WAQ�s���T`�~�eS��b0	N�������ݭ��˜I��:bB�R1�
A��9��6kS����t��G�_3٫D`�ӑ��5y��<�y��a;�H9��1�����*^^�i�c7�R�"�S�(\�+��/���U�@�eՈ�=hp�4����t�-����;��A[�w��gOg�R*��)���[�?w����1.�ƴ�P𦋇�.=F#�YTSv����{D��ڻ�]#Yr	Ζ�z�[[��Тf������8��Kq���Ge>�`�w���L*���ܵ�DQ��<�V�sP>���gH+)�4����<���v ��y)���͖uB��4O&�@w��Bv�HN0 �`LS�
�8+���0u ��Z�=ϭ�����@�G����
i[T�n�Y�Ũ������>=vă:�x�kXY*��GD�ɦ�X<ݐz^�O��q�f3V���?F�Y���3B��惍'�{ ֨�4�U��s�����O�4��>}����	2c�@?0�.���"kW�����SxLZb�oǞ��ϔ�v�[8
>V1Y%Փˢ%Z}�j����
;[i�f��ᶆ��T �w�3���0K�4-�]��,_PU�V�?��VHl�U�õ����-���?h�W�sz��mlfoj�[f�?��È4QgXCcr-�xGM�>�]g��0�����o�~�h�����K�ϟ�RP�5���������u����p�B��W�����/˹��2(�+.j�&��A#�"�y]�T�oY�"���^�	���u�#��Ů�����T���D�׎����[lz}i�LĴ�m]3m���.��H�4m��m��K�qTy^ˣьV��=���Z)�vM1ufdO��� ;��k�6g|�/b�8X*�
���:)b��x�nHA�G֠(�-
V�|����҂������P��$T\�ұ0�:z�Γ�Γ������g�@�����<B�����1�69m>/��.׼��_풔F2ul3����i�i��W >�s:Ձ�	ٺ��Y3�F�
��L���)���ʥ� ��P����YfU#���-a�n>���	�a�K������@�DkVa��i��������\��Y�U� ��o�]t�9����@�XA��o��0oa6��s�v��]���!��d|��H&���E�=�[����C5��ߜ�=���Ҕ��e�W�׸����l���H��TK���46=��������
W�K#f*v��a�� ��"�� �dkt�����RQ�37{���.,��<��>��6]���'Mj�����D�M����,��c�䐼 2�%!�����ͻ���"f*��!*������Y���B�#����cx{���N�>M�X:�;����i뢓s��j�����W.7V�8�KȾM�v�
�� �I�'�&BWB�Њ�[���e��х�a^0%����b��߉Z��w����Rv͑?3@}��{�@�=�cw���B���a=�+>R���s;u����`B`�F������9g����9�Dy������_�ⷐ�$v	=� T�#��=5#[' ���ө��߭�R��(��}��g�J��� 
yċ7�7l��IVs�xY}Ut�֋�jI�Kl�%0�^���g�L��󚬝�v�\����%t��,n��]�p��T��> ����fى�AFM5L<�_�7���԰�K�p4���,��	�k9��D�]1����G�	둍ZmҬ� /sC�3׈;��*2L�R�m[��1r�@ .�H�uG�(֓��⋉��鄉l�f���8�$�������x�h��R�t91��$b2p���"�s9hk`���CDj���x��1��4[�6�!r�v�4]Y�f��ɢ��j�E�`Z6Ăx0g5bq���⏏Z��	"�J|������)Z]�_��������U˄� ��8��pm�Qš��y[��+JEX{�h���<�x�<9�ȻC{��:Z���V��{�O^��-.�2!�\;��R2���-E�L��d�T�^��p�bںEZ�l��6��6��TL}J" sG�SQ�xS�X�3���h��o_wxt~�.��7��7�� 