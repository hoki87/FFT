��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#���������l��U�~�׏O����j9�PY���`T���x���s����uí������P��"��b%>�1eτy�<�gܰ�N�Y�	� {��I�ɍL�ݫ�G�R�k��Q�!E	�5E��.��:�͂2��y�m�-�.E��i�����YS�
��@�H�ۼ��nD��Y�l"BU�.TԊ�=�-�����q���Ǹ��j��ԋ����tr�a�ٵ�]�b	��%�ɔe�)rYOjX5;V��R�������M\�	D��ҏ����9c=�Vͼu��Ro�P�Jf�tRvsY��c�"n�XO��	3g���Q���^�Bʹ�7gQ+Г���$�-��t�8�����A���<����l-��*�|d�n����j��z�l�|Bq�¢:<�)���B�v|R~����gVn���J�i�����n���1��x�	�#r�����J���p��v�j�y������lfW'9��ˠ}J���t��;m�փm��/�4����=me�Y����8Ť�Z��0q.{��KH�6Ը
�v����EW?�Lg�p���/_(y�g>��j#����Z|<d����|�fT�v��])X*��uN$�dG�������F�� ��[`gx��	r���0<�(��3�'s-��m�Q�Ñ�T��&i�㰢�fϤ`u�8���?T���%�������\����ן�����R��#�'F�|��g"���(��5ѨO���C��j�κ��.)�8�����'�zm�UW0	*���?�B�d�={��8F-E�:/?���$�����Rz��[J��{�W>3Db�Ţ�N��^'_�  ���ɹ�ꜳ�[>��a��4N� J\�sKBW�p0��x��� Z'��B>��r���+	$�;pB���:q`��剻�gԵJ��oR5��V��^UrX&d<������S2ǀ5��f\ӡ�Kѭ"F���U%E]ޭ�����{fH���a�a�T�k6i�&Tf
�FE � C�5@D�n<���6s���*�� Ҍ���J��g��B�>?m]��醙h�y��Z�m������ױ����b�W]����G_3q7D��H%�P�T�g�fQ��c����!x<a+���3��` Τau="�^�;�7G��be+9��O&	&��Τ���UH/��a2��e����-ǲ�C��B��9�W��+��S�r�<��ED0����|�$�LW	��0�%�&���肅1�	�"���<�ߖD蝒-���l��V�! /�)80̻$wH_ıPƣ��G���JY�w�#��]��pK��6 ��7/�����b�L�D=����G�q���~��$���3����� 
0�mk��/�ĤaE�ߣ4T
6�������Ki���/(�0��7�`A�7{qKE�w1Wڍ�B��+��uJ��j��E���i3A�U���@7/��QI�4&"%��x:G�{ڻe���h`���mԽߖo���<i�	,�&����a�d����+(�> ���S����2����}(�䁟�y8���K��,B�{gX����*�ʕB��V�/03v�-�i��Z�_z�vBx�}�⽂/ٟ,oBh�\����9����"�Tyl,�r�vU�:A�������ߨ�x���MS��!������0HJ6�VV^����'�z)Dt+�88�w��������\	#�.�3?�G�Y��74E�3cr�g�ܚ����Eaii)(�ȶP�i� ���D)��8��ձH� v%bs�bͦt�l��Y��$��/���H�|-_���E�F�������C�ת��8���VĚ��ı<���~;��={�b�
8;+hU�U�+L�;��S��V�U�f#�s��<լ��ʬ\����$����:++��K��3m%w��O�'�����lh�D ��D���ŏ	��wx�S"A7���h[w��I����m��/2�_�R��Uz1�a(�wl_���	DQ3���ۖ�>Y�������d�y�[H`���2yH k�܈�1�����6�Y�Q����<��E�6$�75�uoy,q�q��n:��F������������U�G�4�2gw�m������>8L�;��\���J�f�F�y��yQ�s8;O��7��Ui�eT�~8��^<�JS��߿���R,;c�Z'\��#�ݠ$L�NC��d���[����sf=˩-߱��˟�V0��-��zcXx�XT�\|�eHA�����4��ڑ1��-�
я��.�+jw��T��/h�xwT����=��R�Z��^
�A�H�*�ѳ��
M%�Kz$���ф�Y��9x�l�XVKd�E�t������o;���S�Z�+}���*�����K��I=`�N����d��ѐN�-]�fX`?�lNg���D4��B~uؓ!�OpS"��ټ�Y*�3�)sS!�)�B�(��L ��#WS���;�f#�U�����E�H/0����b#��s,�G���Ȣ:D�~��/�?x3z�����V��i,�_ ����q�1n�U�B9a?�b"�e;���t0�W`e�H:���4o�Ϝ�}��f$D M"V��5^�G�svM�~(��%i����v*p�3�xX(����Y�<e�
��I���剧(A���مe�t�k�#5�����Obk��g>�J��r ֲ҇A��
�MC}�Ws���ꎗ�ܸi���>��3����ߘYЃFL�\����[�-�c��xy���i��@<��9���q�3(L;o��5��ۓݫ�2��j��|�`4��"h�M���}��A�俵=&��7g1j�Uʮ�M�����ٵ4��)�n鮤�#����D�v��ۇm,e<A���������UB�Q��Dp���0
����F6����:h������\�N_ڣD��1�83h�R8�@O,��C_t�"qC��F�z���@�^t�hr.�G散��c�^�h��bdn��[j�g�F�+�2�AB5����4 �{˨����Ʈ�g|#�P��W�H�_�m2,��4%���>�H��AG��b6��Y��iRI�7<�L4��q��Б���ټ�[�V�? �,�s�R��Q $�����o�����-4R�<���Q�?v�֒���{/.Wb��GD����C��W��zg�|L�M�U�=��p {q^)�5���O	)lC����+��YE��}�'pN�M:��������7Ĝd%�aw�����q�4 �R|1�+��ۨ�%o���>�`��gX*0=j�~�� p^O����2�!�O�Vb;t����*��6#S*����^��tV�T������i���������	)��y�3~�� �N,ф	ֻzZ�v��:Q1�Ab���$����K�1k��KeY�#��k`cO��
�|��$j��K5�x����c��F��6��!W��4ܳ�����;&����j��䕐�ӏ�4�L�ۇ��J��KRaw�!b���!�#+6MI�v(Y�`m{�h���i~��@��y/X	�j�Ja HXZmPQ����f'� �F!w����ॶU�,Y}�t�)|�9���vq���Y�^%���P�/�X��+����V��j�o<c_�ۂV�j)�I��{�N�0	J�vs�u��<�e��N�F�Y�_K�|�;#�����A��*��?�TzO�ڼW��y�G�eo]u�L}R\?X��X��$��n/��(-� �^��^	��*�"D���f��[挅����"��n��}5��?��+ �EV�r��g�&�9�ɠ{&Koƥ���ׇ5�W���_G���&j���K�XJ����+[���8_0ϰƒ�����!�������K#�m:8�������4��N���ܫH,x���
u�Sk���YEK����c���mf�3T���A�U�A
���pH�ay�sӫ���A�N?Ifz|c��C+Mb`�$�{�l���/�d�0P�5s8��T������G͑�������jS�P��b �q�� K���� �6ϑ\���;fմ������0V���^a��JX$FKN1e���1�QQe̪̓�m��s�[6tń����!��W膀S��N(�6��=�8��G����8.'�B���r�SlO։��%��`���� =uC��س�	��ڟ�w#}s�z��;�c�����?��ؖ�]�(�Se:����%3����&�{�5�6D�!�<��1���&y���:�Do#��C,�&G��Z���=��hbv�$?�oNu�����a�F�?}�0��*�@K�~�,�҅%�~dxF��j��"��ԌKn <�Y�z�"D2v4�J?�f����k�X�f��������D�#?�&F_{,�;�I��G��a^>㵋����R����H��U��7K���_QK�����fiP,�ĸw���!�!ױv?>����d-�/��E8�E�9s]�&\��L��W���B)�y
��\��Ŭ����*B� �Z4N@�z�EJ�9�pY\?oy�o�U%�{c�5�{D0ud�`��p�L��_��#Wy/������?CsP�k5��F�_��(�}ϜL�y�b~ERv~,�NM��L�k}b�"�XܚJ���5�6��%�"��ȽxO����_aC��E�fe������srvt����)8�}4���|�Sh�����cM��?�?��S���+Q������� ,��׍@�֫;=�׻�c8���r�R,���)h��=]�)���U��B�*��_ɖ�C���b�Jau�2Qׁ��{H[׽y����~HR��cr.<�H�$SHe��4�O��i�#�RS_\�`�
���i�nu�Q �a���������G�wX��Tg�kE%x��F���?�d��j���5r_S-_HZ�c]q�>u�#�������Jb�{@Ӽ>���
�Ԓ��1��t�;߄zI�Ժ���š�b�,�Ǒ�MF���$�p@�@���
Z,��l���~mM�{��J�T�h�@8��<�a'��1��sz��~�/	��h ��`\1��J��OP�ۯ�=1Vkܫ��J��DB{{5�@���bv��K:μ��@G��H/��q��0��ք��hnF����E���$E��4����D���@�;u��X��4 ��by�f־#��@�i1�X�O%_�{��1��L՜���;�n6�Dp�/�fH~}��9���,�fb��d,���Xp�}��ck�n��*~B1=)L��$6�s4j�"`}&�b��"��Vz �Ѥ��']��Y��P�`�>���]��͉�'O�Y�9 M��Nt�Q���ݍ�Մ�9F�"h�� �Œ�ʌ׍H��AM%����(�Tު�a���#�4'��Gt�5��ol:��c�LC�>��Oj�uS�`��	J�=�яC����gկ\�ɕ<�|�dLȧ0��x�a�-�WUu�wkRB�/���y�Y��6����+��t�Ź+�b}R9U��p8|�����E�[2+���tL�� ���t�8��ܺ�p" �>�@���gF)^Hl�\<j�'"��*�#o��_Fib�_w�j�P*)7�o������5���ݑ�v�0,���������ٚ�6��̆yx�	]��S�(�W�<��bq��H�D2.B�'���n��t���v7⥹j��Al�1(������|��H��%�e�Zy����~z���n�L4�غ��6Z�L��Peq/�ʅ�ZE<�wR[@i�^��tSIi�dԚgQ^��U�Tm��.�G7��H�Y�/�3��N&���3�2��T������I�69}����Xw�$� ��0�?O����U�����.��Tt2��4M���P�K	���h�L�Qf��y�+�j�9Uf���,!�*\U�֙�\�����K;o%���hP�X��2k�G�I�(L&��A5HḐ��H�`Tg�.�`�Ƃ�D���+�y�%T,����i30��^� ���v�9��Y���a2�V�R���Kwo@�	ͳ��g�S�0���8p� �T,�ZB��{Qv���۴�vÔ�s����cI􈠛��Fg�L)�Ip�%�{�jhCf�V.��F��r6�&� �G�h���d�H�Ѓ�oxǹ��nz�;)��>����X &��My��nu5!Y�Ys��Di�S����L��o~���2�����w��;]w��S~k�}S=?�?T�ނa�\4K?2��z�mq�5p�&�5s�0��@|S
B<BU<C�qj��!��}n�mb�*	�8Zc�g3˜~A�� ��������u`\�S0yv�T�Y�yC��Y��a�aW�ƕ,����o͢}�,@ m)|^Hl�_C�KE�a���q������{�F�n��~�|���fW��1|��E[�-i�h��*��.�*��5�叞g8��Oo3G�ɷ!��UB��	k��b4�9�W�+ ���{��-.�v ��/���:�捏�f���r����Tq��n�dK�!�p?ej���V���1	}��)`�)����5#��Y�8�V������8FD:�y�4����V��{���s�s��|���뮷���mB�@��1��3�ɡ�TB��(:���lș���)L�QՍ���M�²_gl5���ɞ�ޙa��^�ә�"�{��ԗ�<�ѹ�yg��j� x@F���z<c"$���[:�BV�^Nn��!�3{$Ϲ��F�� �O�~��k��	[�����Z���mEk2)F��lى��
3E��`
�#4��;����:�uY�5�N<ٴ%/�58=�X^����V�ʣ
ڪs�ڦ>iFe������ˉ̏�P�g����x�pݎ5.�]V(�w���w�`�]ؓTL�џ�sƍek+��6��i�̱��y��T�ľ���e2��}
3%nۅR�����q�\�F���V��0U	�]ʂ�t��Yc �?u4��/.p�:�f��T0$�1J����|�X�6JK��˵Bv�r&�ۧ�r='dm ����MbRt�A��sm�|%���pя�Z��5�oQ-�a�b�����?Ʌ?�Un\8�>h/�=??U�W���^}��������Y���DS{�Y���AjԄ�p!����D+�����wuq�Ki>C����W��0��Z;BӚ?�%��9����+��y�E��~J�\ȕ���3Rf0�av��\q1�K:�������j�N<��]й��!��t���.sm�����&�բ("x[�֓��_5_a`���o^~v�D'E��@�?��/�m�I�\�xm�Pd�,��J�W�8ԓF>* <(��M�:*I�:0I���2#ȵ�b��k�6��(N%n-���$D��{P�Km?VE�n���!�|���c��μ���p�朥�.�mCM�ӹ����DF�:��pu� ��ژ�r/v��0�|l=%&�{�@s����?�ﮎCL�jV��Ч�S��y4���@�d��*ۣ'�TP���T��^��J��b.v�TP76�\��ݥ��om��@��5��<Ӱ������� �dPT��W+U���k��\��ܵ���َ^��6����3v�p����3��L�%.���k�LL��`�	���x�t�`)Bx�l����k*��nn����r[�,��,6͐vb�T<6V���q��OU4�s��^xi��Y/b y��X�L�w������+�ΟT�k�=k�g.����e""����ljI�v�l���J���?���F"�I�P����Ű�чG��I�Lӱ�Rd�_�-D��_.���8��bT˿ϯ=9E�'�Q�B��<�)1C��K�۝J6^���4������4��z/R��3&��c�@�o/�m]��89�է�� Y���qB��S��'���\^m���&s�E�g�s�g)٦��-�r�[y����B3l� Ws�$#\^��\��`3�s\,�ɖG�}��t������t���K!t�ąў���eXa��5S��9 
�t�h�Cg�Qو����B��G�[W�e�0'����{[�3���,)��K��Q�K-p�NjAg0��R�i��o:��:	��R�pO2��~��6|���T��}�S

���c��t��!��9�{e? eJ�wuB���(���7��	'ni�?P&�;6�l*��[8�#Zg8b��W��K^�ũ��������M�y?(��(�.'�p}P��Q��l^������ϣ�W�8�K �b3A̎+4a 1-�v����8"v� �芈�,2'� ��Ȳ�ju.�A���`��&I�i�_s'E$y�ְ<J�9rˏ�#%�sv=�f:!�qX��r����ޛ��jZ#��-�
�yf�����0����@ٯ<�3��ս5-����Bߩ������ 1t;/�Uy�]6�	\M/�{	���Ю��{e�� �[��DQ���;��J�6��n�HƧ|�L��d����4sw�;�e��*�|��9�S����FP�Ʈ�U�0+'�Oe]����QvP����\��R�z�SoX�Q����c���4�Or�n�ӛ�S7X	�Z�}���]���ʧ��=��r|PT]�����S�>��
<yQ!����M��*l����t�^����'����cy��'!~��)S?�$���������2D`W|Rg@�ʵ�_�_/d���<�|?����R��,�)"G6���9���>^�A�Sk�A�.�ҿ�B�׽�:?�dt�aPa�7�!ה��ݸ-���T>�"?&�p�ʌ������bOJ��l���G�#ϥ���9��p�A�;�E.Ꞡ��?�⊰��z!������=�p�GX���h����:�<{h<yT^��{P9��+�m�Iue<N��(ĵ�7��[gm\�HE���ߋ~@a.���F6�`h������
����Y*�^�q:��6<�g�0���w�Z�sk�:� {]���� ���m�~3�0DF&P�3:ȶr�X�x�"�q����A�_!&���y��?��B*�y�'$�da��f�,fs"ʿ�0R��'����/�Z7�G����C����A�P���g�I�^ ��%yN�N�o=���\�sQ�U~�T��t�-���N�AU�Y(�b�-$���jƝ�p�L��|-.\?#��Y�an`�dI7����� �&^����jY!j/jЕ��!܆J�z󎝸���n�	[�O��oI��+w�-i�-@�O�Y� �����E���yA�J�O�q�=���#h�`h)�bp� '-<e���`FT����+��r���<�B6I��V���AQ�ǲ��x%�{�#���lG)^�$hT�r�zSL�$w�@<4b"��I��C���y���/�"� ���!�{o��*h����	��U�S��G��0G��S�.��6��
:^�v<\./�2�h�ϡx��0Qؼ�tC&[.�
�m�C�-�AJp��� �����������7��j���ՖG��(^xP^�jU�����"f ��@�F�����}c+�w��	����r�ǻ�iu@�,�js��n1$��O�a�z�E��bV���E�w���9��.��ӎ�;
���`�%������?%G�%I[���I��a�'��+x�X��]��B��<A3��S8��r�
�SH$��W
16d���;q��C����A�N�;�-s�,c|��}����nY�F�4��n��ie!W�S���k�1U)b������3�O=ᗤ� ���Q�N��o����ᔖ��~�w�P>A
��c�����<��?�TR�e����p?��,��=%��ZN�)g/�E�7E�+!�WY�or�y�������5 N�S��&�bъaB�����:��X�,$!�|��CH�eO�g���z7@@��Al��6+:���SWv�����.��I�
�K�G��`�h�3�T8D�C�Ȫ1��Bwo���d��?��sH����3t��d8;M��1H�tSd�T��̒(��*�Ϟ��9Ux��x|�*�sh�Z���jI��Sw{:U;c��+��w���SD��l5/��%Z&�u��1�7�"�j��[Rģ����'�dR�2 �R  �v`˒۹�����c���c������.��'�

%v�Bȩ���E!;?	3�Q!�� oXn�&Q�K4��g� z/��j�#szlMb��$t�M�h�v%	r9z"p�d�9�FEP(�S\�P�#+ÿ�!�Q4>���6H�k�%|�O	��I�>!x״LP�6DFc}�g�y��)1u��6������u�
��4��г�
�7�L�V�H*hk�����&����� F)����Z���g�YN�8U�)�U�Pe&at��L����o��q�=!%�{�P�T~DBT����.�v��%�Tx�rqt��k��}�4%AN�p�ƴBɻ�"�Rѡa�u<H{X}�D�Ky!����%J��%�Ԩ���Y;�'*��&0`�9d �=n"���0	��=�x6%��6	!h�1�#�Fd���j�#�������^�w[�:�]\vr%���.+_�n������qJԎ��$�q�� ��Lx��]�3�trFζ�|�k��$`�t�o?�2�gq ��E��5����J���o�`@����JZu	���%N����&4x�Nʔ�P�i�o�$�y�lW�8��1�K�qg�l{kيP��lN��j��Sl;rEk�n-���&�N���â����7��QH<a"�h=#D�7��eͷ�%lD~y[�;���fI��1�͓k�5�U�:⧪K��+p �c������b[NM�NA�-¸�s�!�Ҝ���l�}5���������:�o�0��e h��c�{�ͅ�d����TM�����yL=� ��3�pԻ&|�t�^�"q֌V��B/#e��Ml͂�_OY�8����a��oA)sg�c!�}��.a%�
�X���L?�U��W�"��j�V �7�]Es�,s�m�-��Ȕ�Ի7�O99c��YT�}\6�~��S��W�;����I��X�1�D��d��O�&C�>	j�WT^G:���^��ZA���D�ZnCV�W5��a�߫Bs�!��7�\^�iq�p�KS[�8�Ϙ̶@��ś��t(p�p��`�MA'eSH�9UwZ�t��	%{^P4�"�mK��/c�ˤ#��������9lR�{Y�@��,ÐE�Q���)x?T�9N�ot������q#�� Oa�n�[��V'*L�=j������~�}Qz��DT4�#i0�>Q��\����[�vK�A�H�z�d�s0�=����T���t΃IsYC~|�����j�,�M0�N�{BӉ@ty�%��&�2�og�����T�vϣ�7D�F*������d�-T)�5�#��~ɖZ��$e��麘��5nբ�W��~��Zǹ��V=��s�(��'�<�e$��")3�m���ג���S_
w�5�S�$�-4> ~Ѓ楍i �&(Pd���Yi����Z-�U=#�$�o����SXy�[���ڶa�w�B@w��z(!����Fh��WU<o�tF<��X����-����!�@R� �T�B�bk)Ѝ~N�1�_��z�+{�3���Ԥ_�ƣ:�ihU��إ������+��͝c&�9��|/��6�^�p]�$�DV!�6IX>�r�٣�a*���H<���*��_��)�/V�����B_[�l�ɗ'=��j���B�,���|��r��s�n�����<�ӽ���H�:�ٵ<�W��<
$� ���[�e�����+V�X�>��ʹ�g���f,�e�$M�5 ��[�����h��OWe���;����$�-}O�>�T>i�(� _����g�O�6�װ� +��(��}-U���l�Mx+^l.@��j�����b:߉��	d�[��3�:���Y7ӓ*�^�W�y�6��	�d��'G�n�atr��@���C�5p��P������r��p37������~K~۠va����An��v<��^>��⾥+�Q�>0�?氧q�����G���D���v�9�@�F����W���[���b����.��T�A��W���J<��{Ұ�G7(H�d��]]ל&����q�~`
�*�Gy�u��/u�hs��ED���|�#^wܒ�N��(�^��8�ףH���F����7�3�8�*��~X�-��!�e�
KK��`�yˉ�W\���e�0y�W�:%[V�#2�.����?�|���IZ�`�3����ϓr��5�sO��[�[��k�ܴ�0-��`��$��J����@8m[�,�$^��ô��ͺ@���,�C�K7vW:�k%a��j?:��ۢF��CT$�~��@b�5*�P�Y< ��I+���C�fU����+(�g��K$=��T� �d��;
�5���i<��+�&�� B+�#-�3~|xV߀�IQ7�c>�$Y�Lg��#��v.���Ϊ�z��?dr$���)�f�d�%u����%K���Jk�߽z�M�+�������O�Z39S�r���J�ڪ��M�>�7
�IQ*ĝ.�r2&c�<$��%�m6���1߹;,E�L-���!�l1�T'Ǻ��}Ҵ��/��dBꈵw����?�e>�Z�M��p"�j~*���܌��M��4�[�/$S�����)]lIR#�P���C�X#���t�?{C���nǽYw�X
(�j���kDke�K���ai��I�a�oVk9ѐ��x6�Z��t�} �W7�9����ƨ��]�
�ws)�c!�@�CWB�%���4]�j
��㠋)��/�)$�d��Ѯ��J/[�|�:B]�^��q;�e�v�:h��e�h���Y�䝝c��x��P�:ʭ���d�;E��f2�T�.eܽ&xV䦛�i8����� '�� ���7�6J�ji�p)U��W/�j`��&��EC{������r�����J@;?���,�d�֤�	��om=�M�wx��a���C6]��'LK��gV�M��w��FZΙo��օ�D|�u��L�
�&OY����V2"]�h��;��=$\��v�3��>��,�B���%iC�Kl��R<�)���1����ؾ4o*H�k�!���f�v2��cg���5�9���I����I���?��;n?.d�������9�ı�G� G��,fXY�d�4���&���#eM��?k3���v���v�crN�䌆-#A�I�����dҼ�Ⱥ��ckz�1�͈xJ�դ_�}�F|�(%�C���k�i��՟�4ݲ�|��}��ʝ9�<�5`�ȫ���d!�Zц�'o�Za�������
\v��k��l��T@��˞c�Xw�ߙ� ���uI�Ċ���Kq���/Rx���y��Oa�$�S���&�S�D�	ې@>�����8B�̂�&E�#s0�O���ϔz�G�U�Fj�M$�������N�O��`�k�i�,1��v��|�2��#P���}TE�kqT��0N�tt�&��R*r�3�(&�D.Ѕ��6�>����ȩz�5�&��I `3�F`�	Z��kTM'�%��?o����C�g�@����s�w��q��j��)qޙ��bb�`�U�������1
ߥ7e�>e=ʬ/kϷ�p��3�xm�@�%lTZԶ!@�?�Z�(E�?��M�Fh�yr�4��p6��q����/e�����a�;C�M�~s�ӏ�\`(�qm��q��6�1+L�#R{*���(dV���7��&Hx�sG|�����Lb�q�R�n�na��1��b��-S���ir릈���gZ"��қ���E���S�A>i!&��5�1l��5G;���U��mܡ�>�]���X��*�I+zy��y8>*`(�;.gp�ۢ䰤�f�V?��H׫g��Y��E	��Ɖ)�g�ƽo��S����׷Q���:���T�Z+n��j
�K)��\wb��/���B�kE]�<�����S\��"����K�C��J]��s����70��@%&iw�;@�
�q� ���4���E�Fn��>V2z�Rl����˝{��󑖳���BM���!i4�T,����3��3����G�Ϫ!���~����8�6S�@]��\I�
2B��P3�Ɖ��Uc�����'���_0�c��@��l0�'[��b��3��t�/��������5�����P��q�jmpI�}u��,�h�3},��Ro{,~��N���$�̨�G0����uf��(��]�����!�����bS
@���/�
���䦆|�̎`�>į���1j^�@��L��G�MCެ�K�}�<���^G��/��L��uC�ܩ���Tǭ�PQ(>(���%*�
��\�<�λ���,L�4�`Ar׍КG���t\�
�"����Ȼ��bEp��"ɳ���[�J�Q��zԳ���b#�n4?�	�W��T} ��{�1x�\�,$�=8�*?3�i!c^ж�wI���:%��|�K��0_:�h�e>s�\_�ZC��1VЇ���:��o���6V�͆Hyy�9 ���x��3�r_P1���o�qo���p�:�	w�rT�q����Np�;I&�NJ�B�Gr������c���N���yW�cU�
��)�*���,fGwt�+�	������ۂ_&Ȕ8�z���E7�g��N]�K��9p]> ���+�sO�Ԓ�҉���g/:;
��N���5�ߢ�N�5���UF�t��k0T���ٺI=	�	|ڵ���N�ȷ??q��|�e�C��H�i�|�S�� @�c!`�+���i`�?��>upEq6&���9��p���a��^bj.
��n���>|.�k����)!�J)�Z7O:<�d&����&P���J��`�&�m��
�������H0m㒩FJס�9����t����%�/�pS�JlS�ŵ�ԯ&��g�r���)#�M�����u&{�7	�Xq���c�T"��b��|SXV�ʇ�����������/�W��6s���F�\)�"�5F�,!��k��g����K~rZs�pW{1�U!F ��z.������ ȗ��|��ޭ<���P��2��U��e�879��:�16���vt�,��e����(u�a`6dl�"�M� 0_��i��&�U��P:Re�Slx+ƪ�
��P=dh�FH��K0^}�)�	[�d�Kz*R�2˦%�P�6�p<$���n1�)̓mJ��$٘��ʀfL���#s�v�^1��Za�v\�#����a�S3r}jW�z?n�=��%E��xF󓆖\�`����6���H�2��@��1��I]�	M���vEY�N.��������s��(��p�K��nA�j&�1Ri�ac�:���퇤f|Ƌp�(�94�����l㇒�������������`0��,�o�D��l���;����Z4�%�u[�ڹ����z)�6샀>C��$q�0%L�{�8묟���
�{ܺih�μ�#���~��x�z:Q���R����N%M������@�������֜[6Nγr�& �ڽ�RS%�=��!7/������/�g�i'�Q���}�����Qӯ��_>��o9�6���t�\�7�������g��s�&!�|VaC���,�(R�n��IRSH��zi�")_$r��?=Nx�`��:�_��J�������-�o����~2"R��ʦ������VH.�Ƚ}q"%���58L��u}��W.�r�u�gy��#��=)�\�@U}�X���<돜c3�}��.��|�:�o��.�A��j?���v����R�]\&�ݐPc�N�nʉxlD�L?����WDj��ȴtFk��[�O�|D1����8��}��
s�Lp���]J�"��ѯ,��ؐfI1
v��q��8�k'Z�x8�0|�F�>�A!;���t��+hܝ���X�5�4�_�H.�lw�ͦ*���[;����j)��W�a��6�����ycCHݳ���<���f��w����嫗B��a�=^�Xߞ��maq���dT�D�R�˧w���7�نh�?���8���O$W�{�6��6T��<;o����`�ڬ����?��d��*{�,��B!B��@fh�=���7���$l�A��F�$X��i9�O���\�P�����#�č��z�3�D�
����uť�Pڷ�/�Q�����������(D�^\���Y�Om�1�a.���&7eJ5F�t�H�:#���|
�@�wa�3ػ�'���f�j���a@r�N��Q�~&�6�s`$X����Y}f|w(��;�O)f@�иm�����Ck��2v��s^͋�� ��ń������߮�tal��J����\�y��^���D��	.���gAR�Z��A��/��`���r޵qrN6�j�"���a<�����8��=k>��iS˒h�D(v�N�ʉ��A���^?c���gQ�h�[��U�zhn�Us[l��ɚ&X}��?�񠲤�"��=��K"%�fR��h��/0jV�߻��t$㷦^���ƾ#��|&ԀUeD�T[1K�׹�K���5*R'k�B���L�֣��1 ����3�Gx�T-k���%��&[�W����ٓ�F>�z鵽��M̏�C$+jK���`G�ĤAy栟���BA
�P��ԍr�9��[Y��� y�f�s��a�4���D�R)Af�΋^	�7t�{�ga�����=�1�#ι�Nu��E���]|3���0;�U�|�5���FB�I�����s�I([�߸F�2/�:�fd�'7�����Nl^*mm�^0v"�w���v/�S�V!N�&B���k�?�����3�|�i]*.�ؙ���m3����#���)m#��6�,��i���f���I0	����8�[<l�RR�mhk������*&;����el	s
��޿O��s��ݘ-Z��Ű�]M�����H�(0�J�3CE�sm�W������Syb�U �'�^�9a 0	�|6���Ǒ��������W!�]���}3��Y��Z��Ot"[��<��#��ݑ� �X���)��L��˗j6\A�@�CRF.	�%{3\��2�������{�:�;��#���0�a����@��9�_LY�jwM�ED���K�F�Z�L��w���Ĺdv�c1� ��A�\��e�h�!&��3����O�@�r�<���=Ϣɨ������g�Z#"� �=��@���.o�k>?��zy�O���K�=l�r�Ĉ�t�W��F��tm�D?�D��HV����]��y�}�L�º1c�5�N��9U�<=�*�yj`�p���?Wr�Ӭ $)�����JԊ�c�m�[�\�wzf�oR�-@t22��:�E��O�oJ�n<'�G6j�!�Wv���h1�({�Dx�]ۀ.���WՁ|18H���h��^���U�|��k�X�L�@��d�53��\��gf����*̅����R�/�T�+�,���o�V�:	p�#9�:c�R��=��f]9i���5��V"�e��*M�`��}"��BX�vPu&8�8!Wνw`�.É͟�����ҳO�ɞ��η��b>��ȉ�z_�V��*������mP��f�_f{�O��B��Lv	dM$��- Sd���+�d���<���P.�-�Xc2g�o���zߣrY�!��R���g4����g������lh��l4�L��S\ޗ4�
p�W�S*��"R�<R��<W���R��0��Y1N�t���/�77�$'�n����:�ڪ�j����Uٯm�G��R9�>C����*m��5t�����Gį��$��o�";h�o�r5Bg,��W�qfN�lO9���V��3�!��m�*ID5�㴜сX�9Vy%!��.�b���֘��u��յ��,1r/��<Vpz�5�MvNǳQ�5-��o����oӨ�l�����y�ӽ� ��т�D3^�}��
�y��.HYPpLb�à��ks������<8�픛C�z8�,>��i�؊�j��`�i&�4W2n�����1\���M֊�y70[�u���^^���#����*�9Z-*<�lΡg&k�=����~A������Vp�vID��㝻�*�TK[�,z@�V��9��h��W�%>��0h�����}����';a�a��`^���虵�w���(o��`Q^I˄��̸J��WZ���_c4���~F7.��fϦ,�`�C��c�߼'a"B�ֹ���t�$��`:%��B�#�s��v�˼V�#��+��4���)�c��{�W{�~t��RZ�.�DrS�E2܄�p3��p|��)"kH�x�Cv`m�Sem��܇ěw��J��z�a�l��y�I�}3������ZD8�Vbsf��R;K�P�}>GzA�\J�
�DL3�Ű�	������Dĺ��t����d�ŗ�m���7[v��f9�����4>b*%�Ws"X
�3��n���&�����2�c���9�� ؠ���H���A5w� O�v���T��v*�>��J�M<��U{A:���hp�"��\P�_�톻*w>i{&�""o��y�K��ƞ1���Dc?�x���"�����N�Xjn|D}�YI �4"K��C�c�\�"e[%]��d|��}zgZZ��&ج9��5x'�����@%>o�k�i;5�fB���K��v��m�g���B��Ī��]ʾ���^D����LJ�`<+��I��B�^S�,��~)�%o~�G��.Ι=����W��N��L����z�9n��t�x�$�l� ��KM�Rd?�t�gB��jԍ���	��vq��ӻ"�N��80r	'���'D�C��
 ���Rg�o��/��rw��RE�Aö�$�l4nY)�NNx���GIJ/m��}qN|�mG�6�� ��HϽ�3>��D��.�e�v��'�%0��ݏFJ	�29/?��J�i�I���ms�����o6]��r7nWQ�'2�"r3[��7���Z��;f��Q�͚�+�}���P˭��ر�Vf�C�o;��i�G,Z�+�T��B�X�P<ZzB%m�X��Xl�.����鑘_^:ȡ��E�=�]��0���o�W��7���+���H��ը�^s�A�@�WIfI�6���I�9���ӻ<�TN�hw��vg4w��ߖ9� ����[��� rtb���PE�d*��&  f��eIO?���_
z�-�]Qw}[���BbIX[��@��(�+�=\{d�A����}�{\Ŵݐ�_)DmdV��w*���`�g֭p^�~[DEϢH��_>y!(���&�}��֘�$*�[\Uϡ�d�9E)4M1K�A�6\ꠐl-���v��x���� ڕ�
y	g�-4�k��]�/��:l�>:كِL�
ާ�O:�j�Q$��\�����>q
B�0F��JRy\Gzw���ɗ��۰K�"`���m�S 3a�.�Iw%���^������f�#2����]��Lb�����n���������ǜs������uvVUP�2g]��Su���c��nv�#�Ú��
9����Q��!]�މꅯ���H�t��65�v���J�fwG�'@�م�����)��f�z��c�o�p,��	6�z���W��F����8)[ӓ�^��~թ��J��.���t�G��%����V Z�!n��_'����<��_RֳT�;B�/�_G׎.��-�܆�(��*���.1O`���g�(�xy��(Ňi�q�E�^�q�����7��|-�)�I��p�|�g���o�ya�!O�+6��%�r�^�ueѕ�:|h�@����Dm2`3r�}�on��@�����B� �J������b�.�{�*�n�@qL��x�nx������*v�6�6U>��lgd�k�/�Ձ_4�F���?�',��T�u��K6�1k�ma�)MS�<V��EE=�����8���P�JGV2�&p�<nD��Բl#��@���(������67��4���S"�u���KF����p������<�+���1��~%� �+h��KH��̑LAVڢ�����3Lu�^������+[N�J�{�`�
�'�$Y�Z��`�#��E�Ϝ1��ݐ�3�����}��J��>.3�g�cD�v��� Ã���s�T��}W�H��S��F����,a�;�,]���!�9ұ
_�I�BSa��.F@�R��o���W�_[� ��c#}�����_0���������p�J&w7�
��}��[P�Њ	�h/:����Z����ks�2$��Y�ǿ�N}�8E>�Ɓ�41Lƫ\�ۅA��H{��jء�@���4xp���A���e8�"���ԡ	��CS�	����;%�i���9�i���������. �^G�q�=%��c;)WF�jc�<\��p&�����# hɅ%s�v3נ��4���ԙ��0��6"�4�i؜�i�E���(n����;�'�y�-������Q�BH�L#i���k����A���
�V5/�A"<h���f��{��P�m�v;��@%_�e<27��&�W�+L�7P��I�f�d���g�7�	i�.m��?w�"������dk���~����@|j�RY+!���Y��S��b�*v���^�ģ-����D~�)�3��7KC�a#b񶌖Dѱr������K&��3��}��S�EC�Ʃ�dz��� �i�Z ���f9��o�kqJ�QPH *Dx���}����u���ak�>�:�->�9C���B�-��߼���c����'⤎h���D������\�2�D<b�QeQ׳����k{ۭC�Z(b �)���!m�[���K�td�&�$A�j�5T%��ԂW�4E���"�0�����W��v������?F��k~�׻.��>�v"-T�ryq�7��C�G28	�^-������:�c�/�.r&Dt�ӵ���Mk]�	Γ)�hӢX?t�f\k��V�B����kqPcDKD��b�9��T���ɂ���2��Hd�Y�8b��RD;���$l��-F��
�<1m�M����{�6�~�L��͒��7,�P��a8�����윫L"�l�f�PQN
`�GU��&�eAw۬���继5��j��������R�{s��$8��?�ל~�@p̔�����7�^�l6������莡�B#�;+�˔㼷 �R׊]�;dQn~k���h*s�Z��m��g��/3r#�(�9#���lTg�c/�N��n�=IU2(M�Ӊ�?e ��tV8{�9��O���Ae�]�[V�؊1�Ǟ�m���J1X���n����UC⒓zx�5��g6q��e��h���(d;���۽��oj[fp�J�ߤ\�C���G�@Y&��å���g��N�Ng�����BWP�{�U��\�9x���</ٛ���^�!���7�-��3���%rp%�6(�D�q�{�D/��!l�~��ferj�ˡ�$ykl5A�2\���Ӛ����E��9Q`Ek���o�zBӾ3M�q����G�vؐ򒶝�6�y�2㪻{�jn���=��7CmK��&�5 ����7���ũ$��*���݃#yej;il���6(Gw+Ä��|�~��Yl�c���rѤ�k+�0*�F� ˮl3^-ė`3;<�k��eSX��Z�֝($_�;��ɩ>
8B��о�l����$iT1�K��:ib�t6 ���Ǘ��Z�	�,��
M6P��p6�;�y펈&8�'ء2_�Xw����8��D��� �P�%U�Bc��s;����H/�>�s���e͆���9[B�:��Fխ�{.^$�r��"��e�	CRuMz�ekC�¤��ysY�o|]���3S�>�]���Nu|J�	knt��G#��cK;Xe휾I�m~&�f}^_�F	&�\~��iK�����P�ِ초ي���ibh$z߸VHm8��P�WƔ:'/ڔ�eO�^�K��oVf!Ş����JliS��/�J-�h�Ѯ�k����5�eN	��r	��3�X36x�j!����^�{��f����'���N?f��Ďi��YSdrV����q�ۊܼ��φ������v�ǒ7�J5����ur�q���Q^EÛVf��LeBJ�F(I�>P�!�A��,=�Q��ȗ��reP�z3үvl���ڌ�𵑣m\�Օ�q���S�b�½:��p�m�p��A��}�oj��Y�f2��u�da��Q$�"Ir>fJl&��T��$n�$��tE�{�zw/������{Z@�Q�o���V��E�00r��yN��%�r����M��q�7c��d�>��t�[��������馹��T���G��8'��K��>/���0�%�G�.�F&�Ͳ��N�1K�x{�Z�j���t�n|�z����ɔ"�[��	��Ą^ȍq�w��AH%8j�8r}Ϯ�+�ug�3��I��&K����ܣ�\an�u��J��T5ao���S��^����ta���������,`u�mE�R"?���W���*x�"�8S��R5@ۘ]�:X��\"�E��k�H!P~����@
��%"�55׮�X'�[�_��4qW��7�|V�9KR<S�'j����0v��gT�O3,���J#�}��>���
&�{ͫo_n���8�_cu��/��33fz�ѿH1��i��mP�G�Ysn�|���V5mX|4F��=:^���ee����N?_��4��[�1;�M=�Au�����-�%߈�F�|�'��ܘ���"d�ZĪ�O�d�*N2�oS� �]�H��E6�9��p�M7��������QK�� 2
ձ��|6��)4݁�bLS့͘}�����4�����i&�0��cDZ�6�g֍�&8&�S�,��䆀���ʌ!�X�� }�6��U�;��E�Й�A"��\^��Z�i���|���P��O{>6���Wf��hFԯ����$��Rp�I��q�T���T�d(!w��Zr��-�Q$�?�,���oKqP<۠PT���{j6`�fZ=�)P�U`�S���d��[�w�4�I�p��V���ku�`�=kײ7�<$�Q�������Z�&^��>%�oZ����wP5,�}~���?���k�x�ӁeC,���	�	_m.��m	͚�
��;yl*N�0�n��?��u:$�&�������o~�:_W��<����[5
��5��VLCN�"�/p-���� �_#$��u�H9�3�;x���:F�@m�2����у��>��u�m	˛��ǥ?d��(���MvLy�_n\Tb4�0�	�Ép��K9��������(�P%�V%�Z.ӽ�[���vG2פ���ӳ�@-%��B��a�*�lp;wJ���1���!�q
���U�VZ�/P�YH�v�k� 뉵O��:�$�
�-�0��hogP��Z��x<�n_��ԙ0�2#@ǊZ�U�#k?-�e32��29�xC� RAJ8e�H;��b?�$��n�yi܇/
/:�5��>-����a�g��(|�
���qC�� �������(V�����+�
Ԭ�G=�+)5��S�¿t�G�im�yGAk%T��IVbV� l���t�y&j�.�_ȧC`����f�2��v9�a�N�-%�m@\��@C������l�Q��
�#�upr!�ߚ6�$ꑄtXR��:��FK�)6����*���hu��F��0�,x���~yu�y<�{A��"�����4b�� ��PW�$��أ�����-Ax��W��8�~*�J ���aӆ��𠇍��s���8_�h�;vr(�V~N���h��?�H�,P��(k�P#�~[�N峼YD7.a+ר�~n��%^ �wfx��wm�&
�ڷ�a�,�>�zZ���M�|��㸊�.�������Bvf�G����]��ԮV�);[���j-��7��<t�g;h�>������"�_��������K���a[%�O�`&%�k���� �U�T�,��m��=ڊ�X�$�*G���A��q$d��7X����6��B�2OM����MO�P4�������5�^T$�wF4�m� ��N8�Z��+mU|�[�0�G�W �	d?_��L{�rR����CG��������Ao���5m�#�x5�%'#�7FuD�i��@ٌ���!$5�.��
W �=H}�x����I���+�ú)�3�R����|�n�փw�7뱲��s�Ck��g�2�&�`3��߂K�`{k[�B%�5�=(g�>d0w�.�� IW�.V�tBhh�`����	y0c��)�c:b��������]��&��A-=s|�OXZ��Î�����(F}iUW��?f�����6Z�޻�����@q��;��,���e����y|I���q͐�&�h�{����`��(y8/���j+�����M��z���c��'�G���)7�x������Vz�
�3|6m�}�
�����/K$?�.S�(�Rׅ�J��2>�0�B퀯	Wq�j��9M�k�����{���R}���d���0IXdX��a�G�5c�#�!��!2��jTW���`+G
Tj�o�%2�G�1q `J��:V���5]M�e�9��{���z!&�`�w��X�X'�D�EY����[��?�O�7�?��^�T�C�@k ?x�kMq�)4��׵BF�0�����G#ƛ��&���^H`9��T�&LןJn��H�.��D��������7���ʺ;:�EDtמ��R�	�C9R[*�@i�e����-�2;&e"�j��5���-��6��6�E�6��Q٤w�ifˮ�<_z�e"� �,�X��KU.��I��Q����K�����f�D���͡~�yGLǗ��ز�����☺Y<ȋ:�yL��Mu�l�[�j{����<��7B$'V��fO��'z@����vGV$����y~q0��'���m�w�5	W=�6�p'�5a�8&JU�D���96��*8PȰ���݇{wu�ݚb9��$o{?�Oc���-� 4�$�U�є��@��}nfd�Z��aO�0c��n�<u����P��P����y^b�Ö��%����QM;$u�i�~䢪��O1����yǛ�yh�����u;��0�-�.���j��r�[iNe褽S������j�4�x�Ww��|W��D5V�r� R�|yA�鲝b�0�3��.���u�Lz��)���4�[o��tװ,��H��
'��b���6s�p)�?��z�n��k���?�G�^-�x���C��$x�����Pnޜ�1�ր- H��A�t���9N�5��Q	���=��H\����YS9�X�W�"��yG>Ɠ��^��Ƒ��1VR�-�KX��rj�׈z�:SWO�g�+@�xG����P��ݏ�/撄����t���w|�d���+�V�Kj0�f�$�.�s}xFx�NNV\��^�FG��n>���/R-��&Ip�4@BJ�	W�\�"�`���6U%��'ڥ����#����	����g��ijė���@�Y���mr�*����o��0y'	�hS6:K��T� ��� 9r$�XG1�˾1�]�Zö���\��DVm]�h, �,Q$U{� �? ,�S��@YU�U���1��/5e8�3Ŷ�><��հ9�[�p��w-=U��"�Pgآ%�N���>/l�*�� �Yk�A�X�����Ք� Cp�8��TS|�\PQ��XxcN�9?QPt��؝ѯ� B�EZ���m���w��0�i�"cl6���u�%49������p�����d���WW`לS#���ǜ�(�@���k�;`�����h����4~"�zNͯ�,h���NS���Q�s�*�3�	���h!(�������xR<�3�IM�NM��]炢fGJ1`���m�>M^n�~#-ܢ��[��uR��!�Ĕ.(n]�r	E��Rn`nп�@�x �!�@�6��F�B/�%3�#M���D=P�� �n�ҭ�E�K�:�]�V�ue�;R-�d�A���h�J�H"%c6���3G�jF�p��I����2(�vh�6�F��:E���b�r�%~q��"L/�C,1���Q�b��P��\�@ÒC"��g5 �|O��N��S@t}*p0��6�����5�@4}����gt��v>����m���o�d�X��2]��2�Ѹ-v�t��-='�#r@K������(�����Y� �l+v��Ċ�@ĥ;@}�K9�so~)��H�@�5�\F�x]�hb(�+{%��/T�BF�_�D��on�Ѣ0��	�2���g��q�`Bw�� `��e�$��c��,���x=4�.������	Xbt���[��#p�A,��8^�5?�� �o��Od����A����ió�W{�|Y�	�<�b7 (;�ٯ�"��V-�I��r��R«NcQ�u��uà`&�]U-��ksk=O�ޯgb�V�$Ҫ�;?7@
+2bp;�t��b_E�I��Np0Tq����Xi��������<�`��c��:ZK��Lx���CǕZ�qJ�{�!���>|`�)tc�2ʳ�(<�ȋ����׆��"�K<D�z����Ft��^���+K���*�[p����o���3
����Ⱥ��9T��@� }6�W鴢�V�>�j#4�8o"���`f�2��.�I���6,��H����D�g�b �R�J�^#T��G��#I�X�&�0W��5�c��B|��7���|�rr���8i�����j�F��D����ƕ'�~�R�CG�xu�"1L���}ς<h�	�|�Ͱ��v��2�?U�dr����#,�t}W������dV���|Mhj5
J�<�6%'��r$Qq�p$�S��~��ӟJ��r�iKU;��$���Ru���=W���߫jY����v��.��7�(�UM,jo���ɯ�@@d�����z<%u�4�,O��ٻ{�c~��I0򴛷����ӿ����פ���p��y��+�G���@
�<txL�^KHَ��0�	�>��Ðpf�AU٠��������T�iD�eD��+���#���/qP�}(�i�
�k��ּV]��F�J���qߗ�AӦ֢�1��g�&�y� ��39
zI����c[�;���}�*zp#��r[��tY��F�2ۄ����üO�b5�"��Z�;�幓;zk�91��-o�*[wڈZ�WwE���2]����-����?�y��e+��˱�n���(��Ut[�r��~_�w�if���������iV��tP��tcj����_��$��[-ԕd��7�;D�էժ�2���+��a�NE�͔ə'Np��u?&����=.�%��%���ń�	r��4'Ѷ6��R�$a���G��!ߊr\w9�D�-&
��u��쀡^n �g#WF�S����T��?���*���D�RW�8,HoT��$-�/`�}1��UTZ�Lv�f`���? 2�4�%[����(�k�~� �1�0<��6��^�Bw%�P���E�98&��V�P8�L0��x�̇WJ`��2��V���<G���;��! `��#�+RQ}kQo�T�s$d����`?������~��aE�Ke�ۗ5LW)��BJ�o)�K�p��N���9rQOCb}M�CW�?�A Kc�UXU  �Rn4�O�n�J`�&��R��{9�px����k؈t;iHu���S����:��%mGE�ע=-�!�F�����'�*��T9h���*t�������]� �"�k[���UT�S�~�Ia��z��"ԑ����#bɵm�4M��3rsО1s4���=J���S'�B=f�ζ���P�OhLHt�S^�>,6���H�O�fFL�"�K��u���2V�Z���� �����㦩S�_{�;�πD#���j�RT���BӠ��qo�Vn�TQ=��:F�(h|�O1�G�Xw0d���iR�L��m��ղ�f�li8"!dSڑF���￐�R�EiiO����U.T�lώvk«q#�)�l�2�Ƽ�����q����������y� <��T4Z��}�o�ԭ�  G �����,�E��>�j��_�C���վ���k~���K:���j.\�󴿾<!8H�W2�
2���'�$Ձ�Ӳ:��jR���^B{u1�[���%�$�e�X"���S����4� {�"�I���N�����l�ɍ>X�b���f�t��A��n�ZՇ�7+c��]��{/Mxj����;�N�c
}�g��}������2��,� !ҥ�~=�`�V�3�����5����nbe'D�9�l.���:�f#]�CQL�y���c��R b�~����ŪR���ߴ�'���c癘�5��}B8k#� ��>�Y��2,�Iuj.�j�;*���3����v�����2q ����RC�Z�t�w��uǯ��� ��G��fBA��7�`��@�44�qM6����������,�t�>lL�\�K�����٥��mk�AɄ�c6��	�9F����ʋ�1�!��K��142�s�<znTְ�1�ב�߸6�JLx��?ns��:ı�ＢS�%��vC��+f��sE���`w��A��j�� �.З�8^u��-�*�>�t"-ϴ8t��ٷʏ�%�WX~P=��'=�Ø���Ѹ3'a�m��
擅�'��0Ű�\�/�΃=eQ-Fy+z�n��d|3?+�j����5�h!��AF���`�X9�M�?����>y2��Ӳ2��\��m�����~���:=�m`���V|A�ow����WYKd���.�D��.����fZ��U�S���W�]�h�Mia5��pӺ��FL��aT.Fu�Y"&���H^{�'���!���ߴ� B�.�jI�Bc=�Pտ;֋�NV���=M��%p[즼�i}�û-��낮~65����� �]�i`L��]JqF�Z6�}���9U�$Fd	�(��B�����2=K/Q�MA�Q���������M�`<N�T�1d|�v��x�����Tt��UT��՞�;d���94Q3�8zc"ț*�f�C"p/�.�l4J�yG����l��׎�HW����B�T[�qiQ�I�C4Q�4��@K��؅�s�J8��=��
��Ȕ��}��m�/��!��r޿�x��~�xA����2��"X���daC/N#��%
��յ�/�=��Kl���$��R:���y�J*�+�1�%�n��@;}����)����dO���Z�L��:�,-f�+烱��D�ד�.���;� 7�.�/�/�BX<���m~A1{$�20.!�ϖ85q -'��ϧ�����Ô�,��7һau��+�CzTD[��ϭ��d=Ң�m���1""w��x��an�o��K����^�y���Q�M���~5Z>�]�,�j<%f�x�a�/)#`7+C{���^��N�����Qp� �3� Ýؠ"[�B�h�-s0��fj�F��A9�'�0Wv1���j-�_&�S�s���!pO�����.�3 �i�P�&�1��߁�l��^}}�%±1��Ty�Ti05i���8�MT/����k�[a\��&K��ܵ��]r�5�x
��>�o��ɉ(��u�Fv��/���#ղ8��Ց���&J3�c�pkI�ͬY|�����nyK�`�!�D�_�[�<P+�ѽ7l�Z3���]����uD�s���>oז�<��[6M����$;k �yN<�\9�?���~[,]�6y�)���P�Q�1���0h��sz?���|Fߴà�I�V�"�V��6����!O�4:�n�����
�z�Q�}s�� ��dKx�#Q<b~3�&���/X��0H�l���$߆�0T�Q�"X���'�p��5�|U_�4;w�nNrV�m�~�_p�\���g&��jTEI�7H��GW�\p�_ b��2��J^1�o��쑥�8i|�"nX�f�O癚�I�d��v[�oK�g�3~�o�1iæ��e�K;� V�����/�b�ݿb���F�`�J�Ҕae*��ē-q��-�M�d�:d�F�)+���Vr0�w�o-���՗ +13����h�7���!:Ew+�11�v�'#zv�-N��]��q�I�L�à��=����J�F�%��Ģ�:�]��Ŝ��,����U��a�B��R�r	��@�G����ϯ����B�,ͲB���N#z��1�:Xz �A��m���h�����L�?%�s�����Z$��ɡ�q%r�?A�i��� �	�._����L�~[�g:���?�����Q9ϵ=� �h�����oR}�{�3FL�-��C�P�Y�[O4|U����no ��vXQ�����֝���J9�nF䬮��{����-���<-6�b.���H�l��aT��	�
;��N�+R���b��T"�Ph�Z�Ƒ��S��}�5+�6$O��`��ɉ�cL�ݹ��=�JQ;8b4�Hv���/N���S� �R�1��+O>C;R}���>�%!�L�v���s2>.j�;�)V��&���Wd�qR�&�5{�K�����پh*�}�P�MXN�V�u�l���q�'8[-����9�,��i�.�(Ԕ��"�he�;�|��!~��!�n6m5%ax�Iz��T���q$*�����C{ӕ�H�y_�B�(���N3�ߥ#�=�:��9]��/s�͊�AY��jg��d➋���]�'�M�T_N����/���-�.@��TpmZ#��7��rܲ�"������G��U/~����v�E�,��1w���x�۽~M��Oq�x�b��6u|o��E?���؅/"��=�som@
E�l���RL ��е1��:PO�C'a�Ň�ǜ�1lq+�iȥ맆����ձY(ͭ|�L��¨Fr�K��q�UM�J�� 0P��>sw �>h�<l�O��t�:c�9���IĘ8�ㄼ�
~�*�1jOo��E`��xO��=����:�ӿCTWo����2�׉cx��	2�UGs?P�W��q�|�)](�m�3�����SJ�J�� �,g9��:ɾ�01%Mbѝ�:��|Mfɕ�,�0�,Pd�ߋ�EEs]!���B��H�_��2���&Ք�i9DM���1�t�ȷ�Q!t��#:�8�rZ��y|۩��2��p�K��1�o`�d��
������,(�k|��J����MĲ#��l�Q�h��0l�G[�0��Fi�G���<�
%^>�Q�`CW�P��X�@(�-�ز��ث�Y<8���O���P�]�y��sð�ק�n=�;c��@��W�9�H���s�T�C��-�Kz��=�b��n	�P�˕	eÂ�9m�+#P�ʌ\?�tiȏC��6�/@�������y���~듍�k�K`�gx� ���/:���+�L��As�VuБ3�j�k&���)+��&�C"B&�B~b)��	9��y���_�:�ի�~�x��N��r$�9���Gh�/��Jn�c������~< I��8�	˧n��H����e�xx�h�fؖ��+ެ��Ff�G �h90�{�,"iO�B�_��1��̮g�b�)8��e��s�_��A!�'���#܃Vyk���G:Wf�H}_j����$��q.��zŨ� ��-9��������wT�W��7��`L��BIJۜO��ǫ�&]�E�
� <i��c�RNS���r	B�������s2gct�c���FC^d�jg�!��ˇ0$��Qn�LlI]���3X��]�hӐԪ�y�o�0���orc:f�i��|�>:-~�Pa{��:����	=��Gۼ�˄\�2�	! &�T{%�Jn�T��JNL�X!����F�Y�ӆ���c�:H1m�F.?����*`QO����̠��)sۆ�{¤HW��I����m�d���z�A�@?b�H��T�n�C�ȴ�.�o~�ĳ&0��I|}T��H,t���ѓ��	v΃jV�;r�L,��u*]@|a6"�ݘ�ۏо�A:���1O��Q��/�[�-?����c�a����VV��g�mJ�a�=��#� ��=�g.�mI�*�v�;@���&�\�;�B�A�_�v�7��I{�}kA=2R�X����͂�5�zlʖ
*i�s󪹡E��42E���������*n�@�>\�m�s�g�O�/pU?[4h�c�a���@�V�Kb��&�h5CBR��Mj[�܏��Ol�0�Fp�C�l�@����n5y�^)T�1�4���Q��O�F��7���~>��:U9�e�����n��k�q�\_�A����?h���/�:Ѿ!@�(���+��D`2�Zwڵꨊ��g}���~��Ѹ�������N��-�.�3�"XM8Qg�E��d�Yl%w�%�t e��y��{U5jV,D��d�]!�`#��=Q]R��Uw�*�j�I��嫊�ހ7�����,/�%�W�BýS=�ڿ3����������d$e�� ����R�݌nB���_C_ЄJ&r�{����p�5�\2���.2>�F��.�i�+�j��p���cB��mF�ÒT+��ZL ��)��{���_�d>�������9m���^QW5@�Z�����1��㦢�r�S�x��i�E�x���^����ܨ��sk5)�����DrI `�X��=����y�2�_�u�Y��
���L[�����$���Λ��,}(�k�.�Z|<���T�(`�ivo�o�����si�h����adķ7ꓻ��Q�;vH��F��:�d���Kz��ݴ�Dl�{U��{R�]�8K�:N�@EȤ��T�:��D�����z����heeG���#�~�#x��jK��b�m���!�ɴ_���N�=  7f�9EVt�d�����z��Ӷc��;�u�o����1�1��ˋ�J�a�mA���w��wy���3 d���G͠� oVg�:&�@:Tq��g�n�4�7�4Y~\j����
|���T��mA�3M���m��h�����B�k<��@OV���b��A�ܱ:�l�΀�d��{��ȸ����ɮ�2ΞWw��ϥ�=��K�Tbs�-�k�Ҳ�����H��מ��(]�A�V@p��P�Ǎ4��:Ϝ,������PN�qv�$m͝��Ve�Mjk(1���_}�B�i���<j�Nj2É&� aCͺ��`�#k�͐0ΞD,��I|���o��h&?@lA��;�`R�(@x	\��ש�̃�_9�bǍbc�{l�����$�ۏ� �Vx1ЮVVQ�+jATFa+2Y��$�V	w�D2m��O����FOV$)r�Μ�/+t<f���97�6�=�n�s���{��iR�xpTO�h/�K�c�����c���p�w-~�$�d����	f�^���ٽUJ[�vm��浑��x������B��SƖ"�~:���"���ww7�57g��K�2�� ���ǁ���y�O���f��'4;�,�';iy��k=*u��2��</7	O��t[9�u�*���t�`�~pG��L��.e���ґ���]������={�9�mx0�F��_��1/��x,����`�}��Zuw�� �6��Q����*�!F,�k,�Y�Ls�1�8a��[M�o5w	6Md��P���X�A�����W�R�b+�y��gL E:�����R��������W=�p��߫��C�u�lI���ЀK�.륃�|D4Q�	kLV�#+*2r't����gY,����E1u�
�B*�����W��~��������	�0a��~���	T׎���U@�����j�J�/`x1�ŅD
/��-��5ߖ+�`�{\�g_b�����@�j�sj��� �~���aY���� ,	ML�s�Z�ٛ`�aZ�W��6J���d������ ��yך��w�^O��%-(ORihrӀ��U^)~&vQw׿2S˳tt���݉2�beO	�/#�^ف~+�eڒT1���wn�/:��[_���fO�Lk�^�A��"nQa�p����+�:����Q����诤��M3����F��R[5RP�������j0\��|���0ػT���}�8t�q�%�R�	��Dsc���j��l[�}���?����F��Q��� Q�]ΉH婽x��&��I��r�d���}��.Z�����������\~�'jU��1�����%g �ӯ�c����WO1��__�d������p�z��7�@^��Ô='
O��ĉ*��<���U��pB��@A�Ef���n��a�41 �PUGx�e����w-X���u{[l&�e���N����*�뭼(Gz�Ƿh�i�q���/�B���3	H4�R��S!W¨l��e�$~�o|���� 4��c_
�ŠO2`IH~zc��9�~y�h>2��$g�������o�	���J��m�z�����K�}��$gz�N_���G_�a%O�hZW�&i�}�-$]�/����9��&���6�'Y�<��F{҅�\�̼V�$Y��:FZ���ׁ�pi�-��`��KXk���Qqv�X�%|f��*Ο����\E�:p���(�DDg�%W����#4���>@$�Jۂqf������˧nܟJ��m�g��	`ME�8���	 K��=4׈rkZ:��
�8�36���U:��9�)9��g�<���Y߽G.��x&�P�U��W�ĩ0h���˱lK���BF���{,�v��~m2gW��=��<�ޮ����1})�����h�U�]}KU�h��}���'o��>k�~bL�W�h����,W)x���$Y�L��e�-�#S�]������`~Z]2�!P�ʁ�ie��b5��\�/q
OI����˳�o-o��D���Ղ�/�:�nԾ���!����@>�<�/mp3�t(�V�T��?���⁇��M��H��5W^�g�!�ٞ��B�w;nn�"��Vt7;�z� T��֍�!Eo���_�R���Sf���.��r����b)���.�(�qj{���[���K�Z�C���EiUT'?儫�w�jQٯM-�w\�zw���=�j_:�~J��h���m�m�L������55�
b��-m(A��V�؆���%eI+���-Z��6�bL�2��u��D[�����:���u��� �&Ȉa+����w�˻�Ew��g��-�V	��#7SL��VAk�����UFµ �Y�6�y��?�2cX�O¾��W��
�
�1��%��3�(�I��1�@��'���2���Sv��7k�2
�'y�D��`���5��Z�1Ƹ��%��>�|�OZ`q����N�U��:f_���3�	�kg�?�R��ܟ�ڠ��ؔ�bh6+]tE d�='+�����cN|A��"�Ow��wF@D��׮�r����pM�=\F�����z�^d*)�!W�#)�JQ� ЇO���4x9T/��\E8�?3S@)��ͪ ��3E�q�IÁ���Ө��F4�]�L���(g�*��9�}H��A�>���f�� �t��Վ�tLpM� �nq���Dw���-� s�8��&��b��4�NU�����#F���^K������a�aʑ).��!6�FS�m~.3<�3�P|b���]`�f���u1���~/:�^���8c����I��]�w��ר�R��@�^㖯®��m�!O*���#�mi�#�?����2����]�e�#� BaeA��}�G�\��MZ+B� 6Zi<�ĺ-8����5�� �<�k& �U�Xs`rN�r
����N�­��,p���Y����/�Ь���N�=&'�+��](�B�� �%oo\(Ww�����K��nq�D�8afZ�>ؐ~�+$͚�=��_X=��=���*aU��3��XEL]9�5p(>F!�h��Ob�EEˇ�.d�<J�3T5:n0\�5=-O����?{�̚}��8F�P�n[�q���r�`[��BcQ�B��\I��"y������(�_zE���et�E�1e:���z8e�fp��T����$��]UB���.6s��z�`��p0���s�� 	�ß%�����+	����|z�D\���._v��/OA�<�n�>I!Ӷ��H3  ;����q��Q	�.�8C����e�qG��0��$�j~�F?�X�\H���;���s����$�X c�4�27���-���>�y���O.�Ӏ��@#;2MZ���uZ�j�	�%��C(	�V�ǎGއN�����q}m��EݿCD�@j���aG�����osֿ騬fv���:�6��AkH'�yJ{�vB]<���o�j��?=�6VdkD�fo0�&*�{#X�p��\��BV1�?>�1H��V`�[��Żk;�-�?�4��EZe��!�H��i�3	��DQ���hR��޻.�,�u=���a�x���o{� H����&�Կ<}\ �4]s��Ä���x
�o.uZ�0:{A��v}��%>��j��+s�~�* nͭy�<0m�(���|����B|Xjpk^$�"JC/XĈU*��ƨ���Tֶ�=��fE��͍V?y�0��]|gOKE�`���UQ-�Z������j��7��= y",$��\u��ҖS'Cb�H�<:�j���3�I�% ?Ǫ�íy�m����>�BiQk�� ���.�E�e��<�X}��)&�q��5d��� o�S���6� ��fJ���P��֐ |�9Sq��
���{[�ps���#�=�����`��J��m"K����3-E�K��n=U�Pb��D���Ϊ"�ӧ��g�@��c�
��`���(z�O��4;h�н乙��_�kz/nӝ+X�0uW���$���=� �ym�$D����T��,Dy�Ɛ$����R(�ЈT+`�:���L~�#�z�%�/N4��M�	���ܣ4] _T��<rv:;�b���Lx<Ȫ���H~B�ts(܍B����v�[p��5�1�F�M����LI��}�}��]@/�
��-�aãPn6��ٞ�;'��wx�0�,e�c�`\,60��X��#��E��S�F�OuO��E��wJ�M����L14����﬚
�ǝ�����|f����tӤk�+�M�vWz��,��&޽N�wY�۾�*�Rw�'��}�mD�+�>xh����c��+)�ȡ�c��-��	�/�
"�^�����	:v)��_����ۦy���z
�H}ߟ��,B�$�׭��������/I1SY�q�J@I*�&�a>e����������z�D��f�%g�����U�X�Ȏ3}k:m\�|��>����_�X��7ő0��8u6�(�B"jغ��BQ�w�0(�:.ӭ�C[��LQ�.� 3\'�ShhqV$6��	��ד
ݞ�G��uc)�N�|�۔�/�4�R>��l��a�ᾤ�c��6I�zn���R��vю>���������Z�8|�,�vE�	���2ΫJ��_��[N�HA�OxDBP��`䩤z���v.�G��Pt��u����~�g�Tڪb�����}��aˋ'�����T����>���'�<]���ǈτAuKGOw0�H�7f��� %]7e�G�3�|!f�q��k��,����:�xF6w��t�-dޭ��ᡑ�+�:N�|�Ө�l��ѧA)��]��?��^Ǻ�q��[hX������GB�Ё^ V�i\�r����Rf�Ɖ7s��I�c��Kӫ�-ކ�6>�M�^?i`��1-%��R)E�����U8C=�I�ux �諈GTk��܈��M�)�6����ou��+�������ޥ���m�u���Y�בׁ"�:�@|��h��{t����%�b։?~nMI��ݒ?H�T�i�&��CCXCW��}�e6n"�����/�H�����7IlS����l��|:3w��?G�,I��D��.kSi"���r��;�G�x� �<a��2���^~�u���H�2�����bۘu�3���Q��J�����>�6F�{���a]~��L�c`���D���?�,� ��/�+ �`خ��V�L��%al7��R�ܞ�6܇�N)�����å�w��Z�韢<��CKe�WXbΉiQD�d�Fr�*$0Mm|��-��z��걱]xX?���/���_>��|5FzI�^M�_�p��9�_�	�ru�k�
w��
q��|)1u�7��N<�PI�]28�$�jg�������c������6�ج����0i�ݛ��!/�千g�r�փO`[�q��`�Ę;�{����К�
i�n��<����=��� `*"w@o�c'�d��W�Z�P��|g����g���V%桯�U )�*C��C�j�C��5��Q۝�L�_��Ŀ5�n�jJ���#v�n�*= ���tP5/|DE	Җ��&7��O��ı����a�c�j�KF%��501L=H_�'^~�h��� KW�d��Ji���.����qB��`k3��m��0��2�&���Y�{�*6o��(��qb��'�` ���o�g(	qo�!}p�0�K�K���
T"G��V��Xg��z"�D���w�N1��:a��Nk��U���`���=�����nU1Ɔ��p����4�(��#FuC<U�z��s�p3@O���`�ID����}���k�c�'��䶾��=J�	f��l�ԑ�j��鮌д��9��hdm5u��<ߦO#B}�c?{�+��������\n��y	P��6/��{J"AVpl�/N��ׄ#=M_k,Wڬj-}�5恜]ز�OT9mfp} �^��E�s;�Iy�@`n�]�S�o�!�`Mh�Օ��y.��2��U��)d<L��?tF�p;L�!��";���c.�2�=U�Y[M^���¼�b�g=�!p�&jN�>�y��V|?<B�d���{��!e�����[��Fb���`����D�ۃ16��@��A�(v�69x�ol�V �� D��|O�=�����%ۣ#g��_��_=���r�@��L��:��S�R��w���B/��ǽ��)j�oW�v�S<�$�5�j]����צ�Z4�@��ۑ.�-��
.�E�Us0��C�6]�����4��2�.^�����+��G��G�s��"������Ι��� r��`E�r��
�
��
4&����C���J�n��"���R!_K���l�js����d�>�$B{������;��%���]<Bo�G��r��:�{\J���V�&��>4G�RBU�;�0�;JX�9?:�0
A>��U�s�;�-ȣ*
X��a����>ZԨ˅Ϝޛ�}�:�5�[�)�AuX�vi� ����Y�N��W��c��;�J=�-��+�����`Ï�����K����vx��F]��Ֆ�����BY^#��%}�������Y��׍7tW-C�դ$o�ż�@��s�� ]���5�%-����JݜK�;=j��['F�!�C:����_�7�`����m$�48H��B���/�g�A��p��4%�u�G�Z(�e9��/'��ec��� �±��#7�Z�:�B��`�^��_x�^[�Pf�}Ftg�$
\B?P`*M,�Q�^	�ӡ
��b�����0]���,�x
Uʆę@�%Z��M9�b|�q��?�5����T��,H�%t%|�\a>�raz:�J}�8�Ó�0Ci�n0����m�`J@�h�Z�r��`X�"B�O��3o�{�6�M��@��]c��ǔ�l�J�����K�q��)0�Q���C��`��>�!�tH�Y^{�hQC�I���2�*��
N0��0�x�T�E���Z�y��Wf����Œ�>\A�$A�``!#G�D!;9�` )�i��D�<�#�5qj�&���Q1?W���2Р�����ˊ�Pן�5IESE5U@����]��}[��j�y���7�|~����J�@�y]�,c����M�v�/������	"�\��߷A�.�`V�f��z��p�p��#$�� B������z�'�_Z��	V>M�xȡx����Z>k`�u%�'%D�@}�ќ1��P_k��;ԁ�M(��F�V����� ��-�(z7	�س&ÄK�~9�#9��C]��4��paf}���Э�=�dã�̯�LĜ�9c1k��2���p9>��-�4�TRV����9l�n���I�Y
+���}�A��T�B���v11�)m������^����߾MҚ��7/�%��I�
H�lA�k�3ј:�o��M��K� �`/LL�� �@�BR�(�s��9
ǆ��zj5,��PD��a�E��@�Z�֊��V�;�"mT�1/O�n��9�m���$r����w#�d��Fex��H)��{�5��J���h�����&��Dҟ3�T���ΡP�lL�]R�&����n�=r+�:���m�-~�K���Dh��#�U�QT҅ {��b��Tj������{h��o&��Gj��-�&�On�d�MS'J�`���>�����y�q�p�\+��uF�5J��̬�qyt]Dp���w�U;�Z���c% �?�Fv��%��iе�>�8�3�U�K
�X�,��rI�=�c`���~c�!�_�Xօ�<ߧ�t�T�Z�i��Qؠ�̈(�;�:��W--��.��䎕MW��A(�ŗ6�޸o̅�.�+����`���6� ����;;�E��<����+�ÿP{%�y�XkqV(�ۓ| hG��X���+����Ě�����'��ĊgX!'$s�0	i��+��A� M"|�J���;�+!>���ґ�3sp"�H��mX�������*����~�I.�:O�����92�.�FM�dē��� {�	{4ؘ�`��]�oʍ1
E&�=����a��H���NhP�!�O*��/�Xb�Y�������/9`;�,��SC��j��
�4�	�n5��+H�_'�YƁIlO(���Q�G��Fs���fJA��V��3�����Eү[��0tQY��=dWGf^��w9	H���1�Dv@��~���&�96�x ����~��_B�Ic��J:�	��=��⇘�2on��Z�9h�H�Zw��#�u�Bs3*!%��E�E O�"���&�F���CY[�1\���X��9��-EF�;R�En�2j�0��l3�%���A'�"����1��E�x�G�<� �Z�Q��Pn��4zlz��o���ki�t��I�ȉ��H�vX�J��}i��e���$���q��U��4+[��<btd��L���0bC3�(K��}��PEE=ο��
�PD-,����3��;�!�����	G�GpG�%#�<*��7��Mr��a[�3����wOc%Ҿ���Qq�:s�L�e9��.ƸJF�KbDTZ��dEꊨ��X�dPdz+�������;���!G��(��t�h(�=�.�a�5h����m�a\�%�.��"T��"5f(@z�ğ�~ �EZ�����M���AH6���i��̿�S�e��'}��)f}R��"�YG�����J�G�XнZU\�?W�>4�xaGKs�?c�i�!1�̨J	�`��\J�X:J�oi��ж�x���3O��Z�5b�=�Ͼ6�w�e�8�N>��h��=	��MY�ٜQSS�"�cˡ��I�8��P(y(�2nF��"�T3?��h������w�3Qu��I#���jdf�<�>A�Rm`��'Z/��rk��q`��D��
���
(L�'Pu�Ȅ�fn�)z�pW&�v�f�H�Ĳ�/D5YQ�ڣZk:<l�w�s�]�S� <�� >_{�,t�4�U�w���j)�ڵ���q>s ;N"]O�K|-ŐW�_�c�R��c�s��w5ܵ� �R���RdՌ&2������$�'�N'����AW�m�nn5��Az�ҟġW��d��23���'���pm�|]Y[9��5�ӄ�5�q}֛1�pл/�٣���ʰ�=4BD��G�o���0�-^93��m���]���Ȏ�y_;����r�SЏ�?�i�'�H��lH��1U�N�F�f�R�П)�zJ��3��(���rQ����z�!}uΚ�A�ol�Z�9�TfF��!����}�](:�I�Vh���p��"xtP5��5��Y��.cЃnȟ	ӂ/��O�g��a�Ɣ�b�gw��v��������U��TV����q�F�s+����9�Ra9��´e���Z��L���n֩ۤeHlBH�ƂC��۵��ӓ!�.�"�ޏ���ph+����j\m�snt�p�/ �U��*���g�#������=3Zg|�e~�3x\���-��˯��.m�����,�A���3W��Ө�1���i�ҍ�-����A�Z�p��_����(:� �ݛ@@��!��	�e����<Q�8%�I�H�p/���(W�}!�ۑM+T�2u.��_�#ܴo�h )�B�l��Ȱ�xCUx�}�(��䜁i��"�K9�,q�HB�y)z��7����9�����ߘ��O�MMG��^��U���C�i���w1�da��_��5	���W�0��+e8� z��{J5��H7N��M��=l['Kd��H�0b�C��D�Y-��]i��*�C?E+��Ę�ia�tڨ�~V�ChVP�Ee�#����K.lm'��b�w�qd_��� (���d2��Rxt�؏A=3/�y D}ن�_A��_�.�)&U,��g�F'di� t��;V0�P_��'te�uw0B��~�F~ϝD�_z����W�u(���pv�c��uq��|Eb��՛ܓ20[���҂qDi��;aN=;�I��zۇ�>����7�-Z���*�w
k @�p�y�Xӧ�A m�a�Eܶ`���n�XN���Z��G�B��MS�߲G�y!��Nv�	E}���<�xL��6U��HP$C)�t�k���L<O���	�w��NB]ܳs0���IR�]��ڙ��-Iw��& Y����+�J<�*g���%[W��}1���~(��SO�f�{��w� דuvLp�]��eI�elS�Q����32�fף�y�d�8`y'2�O*�5Q3�d����b�l�2��M�;�&�O
PeF�8��ࡼ3�1?�dY'��1e��6�������QZ��O���؎P��=��׸�yj�� �<w%�_�Z��qB��肊��)�/�aD[����H~џG�/�q�c�;���"y��^��q����2[�����ͪGr���H3y�^��lۏ��.:��<B��K�e��2�B�ڝ�N�G�g�S��ciF���jw�Kɏu���"7ֲt<!wo Հ8��@�4��~wo��	�2N0шh��#�7k�K�ê)�m�J\�(\<"���&�GƉd�6]�Ey�M+�`�MC�`�7C���Kh4�|F�f	0���l���0E��\�(NʮS��s`g�U<��G�Or�c/��TB]#�����$�$�v�`�[�P��#dNn2�u3�V����ɹ�QT�c���-����It��7wh�1�� �?J��g�}�U=�a/u4s0i쭫u��:�����7�pm��:z�1L�%���ד�{|Y�V=�>l�	���;�,;~�G�8���L�o:��J��N�"�8�d��H��lz\	Ϥg�udh�[t�U���B�)-}^Z|�~����%��ɔo7��0����y�p֬���h�
��}?��62إ������P���$�0��-�2���/Np�	��Kp����a�k{;q/�����ɽÄ����r�!j�;cy�ø�_n�ȑp9m�qF۞������9Lh���aI���!!��%lb/���-9%��F gO=[w�>GF��1��ԛ8�ڟ��ζ�8��6��.Ƴ��>5�-�������8�_��^f��%V��T���%�$}%蔓#�j[�Q	�޼�"^�qsu��M�.�7�;9Y�o�ß�:�S�@c.�=}�k#yy|b�Yq�U�]�1������عq��Ⱦ/Zt����	�	?�#�ee��$�DTh�-��}0z��?��&�)��A��6o��d�0�i}3j�M��B;FSL��0�1��u�&Ƕ�����rKP��3���7@s[����5o��C�Q�M�Khozt7���n�汇j�1N<Qc>� ��6�]3�c�a��N�ZNx��L�~���
u_'����y\����1�"��z,�=%�
��V6/�D�(e�'B�$��~GT�j�1����ȥ��c����k&�FG_y�-�#����2�3nUnԭ=�e-��˖�&����)�Ue�������������3��\�<I���r�|�SHjBmraK봝���e�{���Ϡ B��k�:���Ʃd�o�-�̦[�V�D�P"���F):������.�ÓD�]�j��O�WVC�wi�QtS¡��[��N���t�(�ż��6	b=�ͥ�X`��#ꢇ��0�뗒v�l�K�e�8�HZ��H����ۺpȹ�z�X���b>;@lM/�G�f��s���w�vr96���_\����zgW�8=�	����2$��� }�`�,>���)����)�^|��U��ƺ?�.�I�CC'3���̄�X� ����������:ahkz�!̏����g*��r��%~(iC�$����m���a�=�lE�6�^��v�k� �����4ik��Z����;m����7���B�J�� )��+ °�5�|?���ڭ�`�:H���B�^�K���s.�Ǌ
\o��jb۝Wy�p���S�0���~��_=��v���a�W�l7��}�f�W����e��U����5:��7���s�����9!3���nhSsy	�B��+t�ɮWa:�8�����%�Nܷ��a5��O���|	˴_��4�x��Wy�B�a&�����n�~�J��A�O�/��)�Ha�t��
����z@�1#�{��m2R1���"f讖F�$0)</Z�0	poؙ��7��.�f4�iM!?F���Q��#�r?A\��D�cD�5Oqk�2�y͊���Ȋ�O��C�����r�xɬ]���Q����U�=�:Z�I�f
[����_WV�?��ٜ�V�DX��s&��~d�R'O��͛iC��Ҭ�_�}ku�w��G0� ����^�O�6��J�!U���YsX���s�V^}��p)b��Q��<������s
�t/���`-��h�b���'�n�M�f�E������U�e��6p���'[Y��B� �Ȓ)�[4��]�ds�f�{�f�����~��CJ3�.��Nb�D�$�<P�	r�52��lp����e��o`T0<(g�����GL>.$!�ft�gGd�z	��A	>�1)w���K�m���Y�i�%b��Uѳ_��+��d?�'�^&  8u����w/�]G�
s�����Qg��<�ׇ�G�Ll�xB�{;�	B�0��ՙ��2�	�_������B�7��bo��$�VRp�e�tL�����;g�R�`�y��1����t�n�]6љ1s�?���R��bA��}���f'#`g�U�+?�P<����>��LȺ�]w��?O�w���5�0�-���}�Ҍ�G.8m�o��3Ti*���d�'p�m�v��qlF� �#�K�������nS}�mlR>a�ǂ��$���h�)����5�Ǌ}�Kg��^	6�I�6�e�Q��n�k���I-�_)_d�����V]�m�%s��2�6�s��� ��8�n+���'*L^̈�*��R��,�w��h���U04}�O�X6\�V5���ZFL�.	�3�c9���L'�J!
z�1b�4���Ci�/������!LM7e��,H�S�m�~��`j ��Y|k�L��	���\�0��ґG��X���J��z�t��m�(E�zs۴mc)ԯ���O��`:ޙm]@e�c��_�2=�����<������D��#Dr0=T�7�1O�KK�1��殘3�}R��P�з��޻s�X�'7$h�� �uj�u��.��2r���5kh���45@�E���+~�'f�j|GB"��GQ @p|�̈́x.�c$�:��k��.�Ƈ~�;6�=����������e�?�ֳ��i��o?�+u�[��A��p/��#�*�0��	�%S�� �j��فL l�E���"=�(L8H�Y�&�p�3ӈ��6�L�r��!�J���lϟϾv@�Z��6_&�έ����2AA�W�~�ql�vS�Q&�����!;+)7D��6!�G{��hR��&\�W}�S��.�,F����9!��4A�ݯ�\\z ��=�k^�=ԔgOi�r�S�����H�`��T-�͞�F(�)a�!*��1���H^��+�5�D'XS����ǅ�~A.�Of3�#������z�匪d.r�僢R )l?����������Q�n;��"@�bfҿJ�ٽ�2�#?�e	�G�#*�c��i�p��*�_���9�>9��=Q�yҕʊG!�Iā��dy��������d̿G�<VL�+Q���g/eJ�J�/�nr8�0�(b��V2�CJ֏i�a{G�x�9�&�BDŲ�L���9Y��n���xg���vJ,�s+M!��g^D�S�*�u�#2�1�<p/4A�y�ܠ8EP^�p���4���x@��q�CmT�Z���b��`��S������'?���zjr�W%}�w��!���)~�M��%��GU�~��D�[[b�ֳ�lr40{���0��S��Qz�vW	��b�̒C�F��>��Ϊ�Jr�s��MȔǮ���:��� ��t���s���[��"	���eƱ�fHq�V֡���*@=X���m�G�#!��vwj|��K6!;[��_�PJ�3��{�6	#��;_��V8���7��_���\#��_�SNC"���.�+�ҷ��WB쏀�e3���%r�c�A$o�SAT�-v(���^�]RA�����c��I7��FcV�T�G����iˁL��,���D!/]��ʅw�q����X����ie���E������� m%���[!��=�'�K�O��#�R�\3�.Ymf:�x~�8��F&�]��,�q��
�}������E�����H��ᇱ����%a��VI%�Q~�>"���n��s\ o�N2���>�����6����˃���U?�M�ʈ �BHJN�Dt�hZ��P�/�V}�)�Xtݥ�^���,��}�n��a�.$�Ծ�5kb��w�21_/H~���)�+��r/��Ch�U~A
nG��G�"��S�ϷQ�|������O���[�
՝��(:"�A��(
A���D-��,��|v���:�$U1:����d��t��{[��k�F= Uo�ʹٚ�z�c�괸�fl&�OJ8�V�`P�ou��(VjԨix����1�t�`U�C���0q���,�ዪ��~m]�ꈁrR�U��/en��dJ�NF��&��������Dz�� �APQe�7^��]�nhp�z}�B[�8��;� �bJ��L��C��șg���D�t�c �9ұ�`-��O��f-0~ZY��Qze�ބ<i��N��i��G��ײX���dO��(��j�IV�����}(�.<?�e,��=�n=�¥eL�����l�6�;�vR��g�W�Bl���@ȸp���P_�s��]@��!��]7��U8	�9�S�N�����G����j�>9�i#�ܚaάn�;)b}h1gF�je���u������ɽ�ƞ	�\9�J�d�?oM
�Фx#���F���zqY7"����Ğ`=���q�Vݶ�~O��]cZtDj6���?w��V�?�.��c,ďB'���c�I@��7��[ ��I��C[]����2�}��3%��F�E���^���&��毘�'��؝� Q4�i	R��3�J������\��
�־9�.�t��o�nVp�)u,ʗ-�̦e1Q]H|�ڑ���cc-��V]��h]T�ѯ�O")@�>2�C��=�`L�p���TME�>Y;��E������ .O.����D��lYQeP�Y�'>���2k�Y:�A.��ѕ�J�{�.޸e�(���;�(u��o!6���ܘe�1ۏ�ZLʐL&CƇ,+�[���b�;>��]���hehA����;}�j�6�\ʶ�+g?ʉ���e2�E2���>�E@�n~��QZ�8f����]����]�6��������H������,�#CF��g/��4ƄXB�����a��eo#ݜ���u���Qٗ<	e®OB����$��b�Q��[���G�wwp5f�W�+弃n5�-�������_ń��~R�|]�`H}�
ۗ ҥ�&�[��Cy��k���$�,����Έ˶|L���F켕q��+�Ű�::��#������0 �bz��$���mQ9*甯� �ڎ{l2~����Y�J���kx��}�k��U�V"�H���הxk��5p�o���d�Bjs^F�H׊��p)���NӔ ip\=��RA���/�eB�������y�6��E��a~�壉��Ue@J]D����lg�UEq���>:N�"΂�ɘײ�O	��A< ���ǍDH�fXo�`Fș��*� �d�����pb7H�(`1�����Sճ�2�7�X޼0xV�%O���R�RSP��'e~u�| ۸t��5�6�G���'�*��%GZu#�g)���i�l���PD�_�.u݁��M�*T��8����i+cq�Ok�%1�7�.�y���AZY��6���c��5l�ۣ���`\-r��}�-�=L)�H���h@LVz�ꍭx�??�Cd�W��ڳo�����V!�Ӄ�T����ʻ��Ό�W����&�p�$J�3����bJ����q�.�f�Rj�R��3�<�G���
iy�<�n�,*�	��r]3A^�4��sXB�K
F���/�f�{�NՇ�Aӌ�D`���o�r �it*��:�;��z�� +'r�/#�{Y�֥[Gѹ@yɖi�:8���9�����!Q�۴�i���].t�7��
��ح��|����}��3��l�̖����v��T��kL�셵 ��4�}<��F'4($�U���OE��#��vQ�P�a�"k^�LwUbNhf�YR*����f>�p�e���ZȪ�狮�oK~���ڶ̝�V�]�C�d��������V��������:NkQ��C�\r��o���J��q[J� ��>��r]��Ư_�UO�k)+3�i(½��.^|!�1�,�!�Օ�Ҕf~o��v��`2�:�Y2T�i�0�r.-�������B�Ą`�[��F��ՙ
��1)�ǭ�]-�=�UuXx������� �0��������"�%�Z��1]d��d*6�.`d&���=�M(ߩ�9Y�&��Eb�Y��k$jsAh/��K1	1�J���*�x��u}��4qqwH.a�����Q�7��v���a��/Uo���]���q���M����~�!�R�Q�F�sf%Dբ��+�����ג�0yv�u��ɪ`�kPg`��@��M|i�"D������D>��&�}R��X�wv�'V��
���������8i�)��F����l��jx��r8a|��)�����8P�"���,��T$���Dd�\��9�D�;��&�04�֞�/v8�D3�2Zra0�f�OԄ�� 0����(����7���.�r�\T����|7saҫ�&تNO��;�yQ4P��-Q�2N㮆}#%�'BFtW���9`�	��5�H��7H1�|���Vs�TW��:�s!��e-�l�Aa�U�nN���z<�&{�˱�Acz�a�0ٙ�����:?���(r�t�32Z���j���ҐYG g�Þ�Gd�7�&������o��*���u���/�O,�6������p��6"�����7F�遖N6Oy��[�ɋ�����P��(x��R��ڣ��,�+�k)+0J�
l���>�#� ?���j`�L����l-�+1�V<J�w	��,�!����y�6����&�v�CW�D���)kY�@r��^�jjL�Q�&{�|����V4�8X�jCx�m�r�ՙB1��0u�̢K��s�@Y-�%t��o���-XL�l���A1�������ޕ�K�3��h�����&I�B��O��W�d�	o�;d��ڼm��g)᳨�k{g;��F�o&����$�|���mo[�X/�OT�[��P$x$[p���Q�����Wc��/���������2��FU@P�c��u��|C��S6t@�:���?.x�3������W��}�ah�c�G"n�C�o����fQ!�������5$	���R�]F���A�R5��Ļ���Z!�������ݢ���'>/\l=l�Dtr�/K�{����T�]���o���螟[謌[jB��1��~P�|�o�	�1㫃i��]
��m�S-�_Y7����l���!Y�j�+ç�L�������=���r<�徼4�pEр��s�L;��G�{Z�Ƃ�%/����S�v�Z4b���
���2vB�z����H�;Pd��a�ϡ��@�=AŽ�S����������{w��m�y������C��dR-�E��N��Z�ik��-��u�\�q��9߬��cT��簸���>�Hexx�:�jF��w�������]\�2�_h.��+P
nZ~��շ���j�	Ľ�o����rBJ��P��j/h�Mr�����*�]0�����J 7�P�kk�O��I�Lݡ$j	�L��д�D�$q��X�H��,@��v>
���R��Q�ѭ��U���]�]r��h���C9����*��)+i�����"��D[O�eg�o�U���~~�ЯH������bG�KS8\�mf�T�����올�����r��|���F\�?���Z��z}�76U `�)k�W����3�6|G-c�������ҕ`�����xC��(�ėA^�9!�}����]�f�hϪ��4�Ը�=���g�)+���!��{3�y��X���%؂<7$��)g�Ӽ���[͹�?ƑG��=�ް ��cy�?�Ū(���ZXs~ �^�.�Lu�xvվ��t U�ʗ�DIx�L=O�?�xLA�0�*�J`����3v��?{I,l��-�+���K���~�?[Z�\Cv!Ѩ ݣu�t�6AF�l�>�n;�3NNQb_݄~���=l^ƦT1-��*J�F^'a��%"���x�{��.g�2�~6J�w�gF��4�g����@كa3V�����ccO���ę�򄴛���ݺ����瑩_*��țڜu��;.�G����O-�zC&x,\C~S~u��*�WTŏ����F�޴̚UuN&=!1s�BG� 6�P�)c�n�bf��˩�pf{��$E��)O����r�'��k�s��_	>�n	vS�'~o��l#4�#4N�:7����y��o��i�i@��BS�m�`�pR�����f�_bq��s���u��������Pَ��������O��9�Z7�Oxdg��/|\�.��{ �R�.6Lq����؀��+Hj�����@ʪ��'��3�Pض�[��>V:��e�"9(k`�
cb����RIt��A&�9I�#q� �eW!����WKb����m�8�9�/3[o25�]���y?��a$v𳗑U�!`�-��6��Z0�Z��S�b��w��K�jЭ�u�k��(°��&��.a!�8��8t���hr�E�˽/���&���g��V֖^�,�o4������VVA������83⎜�F��NI��~�R�,��ƍӴ8�;�S����Y���Τ���v�L�!�I�?F�Q��K��&��J�Qea��!��Fމ�mJ%���u�#���KQk;�lX�(Ѻ�<�(�G�~�~�P
�v�B/�v�q������jr۱�iD�	*n��?n߆A��\��ٸ+�
�<
w��A��fn��k�a����]�{��R�J�*�4˧��M�0�ʰ�&����ʼ����c�Z�A+@�{��c�YJ9n���w����Jtv(;��{s�0	95��(�\q&��io��{���z�b�����bB~���׷@���;��S�3:Є�LP�1"�C��
X��l��IWt�r���f�b����r`����D�w ����W�5�+�TN4��p��4y���zTļ+� L����ݟ���tz|��٦�u�=T?��P��Ջi��f�槦@,Z���R���2��!Jq��A��|a�u���aiMdc�t�o'����y7�Ʀ�;�M�s$�T����ᓨ"Hy��r{��ý�K�aO
9#G�-�Z1eFоƝ�C۽l�U��[(a,Yo�����;���+������S�a1'��3��UCgox�k4{����bp����p'l���W���\�x
��>QC
_D�+���j��>��-���?s��1#�^/b����}��Zj�$-x�S:~�F9"�QB����F��QZ"&Y�D0�� ȸ�����\bf��E�1n����Y�]���7�#��bE�!`_Ӗ�%����y�9���`���,��έ:�䨒�Аp,��fk���F!�v��c$�ğ�wwR>���� vS��UN�W?���9(���Իʄ���~��*�g�q����"�K��}��������e���p�N�jr�&r��9��L�׽�9"-���$�>w��! ~tKb�bj�m�W�H���ј����ԘN�$�df��9}��Ü�!=���3lűF����� 8�����k��1@QĬ��H��C\Re&�s�!�Ό�������ŷE[�0U�4�z�?����6P��xt�?�B��0���ay�Ad� �Q��L�/�F7o)~�A���0�����[�����`ƌ��d��������_Q��#�G��&�Uʯ��s�O��<�`�-1�#�NL��H4/��g����TH��Ú8��!-�$b��`�g,nF(=�a*xM�?K�DB��r':���աlu$�!/L���dK�w|���%�N���E�Q2���ͳ��r\�o~\˄]'��<%-N	���3�BK�ʚ�
�?/�1���W܈V�3&�->��+��71�̋^k���N��G��^~:��R����-;y �p� }FG���p��]ѿ�b��Ġ&B��N�7�����a<YeAs�'��K9�;��Q!�Ǯ�CcԭマT��G'u$���<���y���	68KL�2\}Ki���p�K�����6�m��e'E�f^s7��`!�K�ۃ�:C	��n�P>�vW�jQ�:#�%�E�ϥ_�j�q��)}�4�H�Wj�T�4��RP2^�l����G�Ĭ�:}���7����,+�;��F!֒��?���kh�Uv:-& �J�8�h� �.g�>{x��V�8��r��-y�}�
�8Y��'�Њ�f�1L�����`˛#��7��
��/j>뭎�&�-�X�mf��_�Au�f@"�1^�� �b�ǎGs���Y�F!2��ʺnm�L3lz,bm���~��]����g�(�go3@:�6���]P4?M��\������f&;�Q̔�ߘ�]o<�sC���)�A�%5n(�0���P��Ю|"@e	�L�� z��b�t��R�"8O��tr ǌ~u-�#��6�=׈ۃ/9��4�ۨ��Fx��$6��ƥ� p���!��ģ���s_Q�荙�Xp]�H�,Apd�Z���/�i�l�Aq&�$�4T~̍0r�����1��߮W�#�W�����^B~����b���ٟT�11�l��1t���8-�3t!H��C�F���]�<	qf�}tTd��l;���%��D�����Ae���s9�/��Mp�'Ⱥ�`�e�Ϣ�Y�e'�����o�]�Z�N�4�B�֮�ؑ�s����6}`�]���
LM-��%=���Ӽ���qDɳ��*
Bh_>�I�l4�,��ɰ:�ݿxk�#>L\��&$�A9 ��	K�a6UxWon��|a<�>�+˸"��ҼF��Lż���nl�O<%A}[e>`�(%���^ B@����U'ա��>�Z���Y���(���TσP)?�22li2x�bd�)��f+Л�}�l�ٗ�+@�����T�� �d�ٜ:1�Ѡ)�(���D�ٞ��*?�]x����I顭a�ݻ�Њ� =I����ŧ/��3XA�P[ܺ�Wn� �F�̐���U{��E#�Y���:<[_&S���s�ʬ���c�"��*�Zy�
{S��Z;��������y��V�5�'?m�`��FBiD�h�̡#��5������r4@�2�	´���hQy����o����a���u����Yq捭�*^+ݚ˴����|�ċT^��������1�T��]L��-�R�y4�27w���$gɹ���4�M"�Ӣ�j:T�_AR�+�amN��w�����t��"b7�xU�)~|���f�b<!���!\�ons&{T���7Gˈ\>�����c�6��{�)�Y� oՂg��'�ɢ�ړ�Ѱ�T��Q��a��e�YR��Fl�=v��&ox�>:t��ۅ_9��������T�9���/y����l�R�g׹�F�R���/D�Nc5 ���Y�iJ�8�B� ��[^a�7*���.�m��9tgcTB��/'8�i�"7/�!~2�J��J�_Kl_B���{�m����y�u1�G� M��.�*��PE'��ȠI^)9��a��I*	���d��@�L�E�.M����{"ѹ%f�<&SiW4J�t��)J?�4\��N�I7BF��!�NN�yF�xRΜM� ��;u�<@&_����b�cW�֨������������w}(/~CSUfi�?�7	��Pc0���p.�8�pA-�� ]���b1y�6���5Ů?KUS���g��ȋ��O68O�7��^-'��4����A��+<*��g��등�Jm3k��A���Ww�����9T�zp��,2])f�}/��[�Ǟ�D�>��-=�R4X�\�Gzy�.�Rd����=6\��Td����^%3�l�3�,eA�{�QT/k��͚K��o�d�1�f�;�g�C�{����#��.�������]vd���c�(���x&�O��YŠ��aYn�mJu�/T��㬂t�"�+k���yx�Ki���vC,���b��Q�
E0����ĪȦ�7��/Õ���y��T�u}	�]�U�
G�"c� 5�qn��la\��0Tse����CLJ�z�1g�����"�����ob�m�5���k���`�ph(�T��L���~�gԏ?×Hr���:�'l�����y�ӷ��`�0�M���)���L�d6U�0`}Ӗ������&�(��<Q��2I3[�u�H[Ax͖��~",�����^q����G4�Lǎ���.�� �u�z����T)��k}���x~_^�S��� m�r���iF߯�3�7-�%v4d!��O�vv�N�k����x��%L�B���������:����{)�(l��rd~4��i1"'\�lN N�tḻiYe���'Ѯ��b�?�걪�[*q�w�4D���0��,��=� ����_?O���$_��l6�{���3��k*I�$
ރ���)�ă�$�x�k>�1˓��P��]d.
`�7�Y"I\�.��`.��q�H:��_�]�+�h%w�ҩ����L�]o�^�"�F��������x}�V;�TZY�)$�U�z�S?gf�2�Z�Z�~�?���l\�����~=I!����
W�H��'D{J�̄~�JYK�N�EJ�{�����!�W����1C�b�Xo6t�L�e��Z�F ���^]�+�
��g:��[rR�v����t�!K�5Sr��,�c���c	��5Wü�f�ފs�6�2�@�?O3�M���Ԣ$U��	t:��wB�&���^�m�i�!���T�F>
Gb�Xk��Q�"X{ .����>�U��O��oL��a>�R�+Ǚ�V뽼[ΨT��v��и��T�d�)��8N�N����5���ݼ���
�gssFkL8���[®#�H�_=F�.Nl<L��?5-{&G���8�)���#� JB�.����*�}��{������Ҷ�@ �G������T�+����B���9�|�(~:}��.%��"�Rk�~����o5�k��zh����[AtqM��x-�U�C64y����A�
';�h��L�R{����f��ƧK��Q���Y��e��J��N��P��b�'W(���S��f�ir��g�Za�����C՚�a6?7	X������w!��\N�G�ӡ-j)q<�˔�@9��x��n@���Kg[c���6�����_9`��_��!���ҝ6^�(3�ޟ$��^���� \����s`������	Љ�ż������NFg��j�F��������'3���!�H,�WA �;"�ҹ� ;ɗ�m�-Y�S(���R�}T�by��a���Ct��K^Jy%�Ĉ�:؜B�Z��3�q�3ڄ��8m�q97��ș՞�>f��<9�NϜ�"�.�W��vj�6,\�6�D���E�bt:w��/;sC���=�&���3>�BB>��F����h ML���`�����G0��4N��>o�S'��2���.	��3"���a
�}�͜-ԡ�I����N�%)S�bsv�����'�N�yd�?;G��(��#�H�m�g���=�����ԘW$� ��&f3�R�)�������cO����x�ة�;NFw�C⻽lNr�_�ؒ��9}$.\rU��� ԍP�6j�w�����>�$�^���R��H��cp0'�2XR�@d�'��ﮭ.+T�P&�gE�C�� �F����&����+2��Cb������u�1�9wM�m��Z����.�T��R*]��u[�i�U_r_XR����N��0�5� ��¼�9ǜ]�6>��+����3W�I�v�4���Ll�R��<?�������Kǧ��k�U��Y��ݘ	c�����	�VI��D��i���N>7[��'�������s~{�󛃫F!y��R�q̫��h�l�"R���A�1�O؄H|68,/�5��Ì�i���Wu�>e��|�?-,�Wr.:�/��-��޷F��oY�ߎK���?+�=G�i�s\����(}�.�]��B�Zn��xb�R�n�ea��Q��\�����|��hB
��l	��͝ �]:qd��=*0G���CwmN��B\���s��/����j����|��v��N���ۏ9���\��\lR�b3������j{J}����Q�iX� 6H�*V�6,�

;�!���#����+1�>3xD<bn��Tză��mvdJ�Dh�M��!�)+.�01����Ae��{�8�1�8���	P	<�E�{���X�+����&��k^u+Z�G)�O�a5ot�Vݓ-A|�c���R�X�rh���9�� uKM�f;>brK釶w��&	%����������1*L��S��^-�7p�iK�
�#;���S�0+�5'O���\�l��MyT~�mt\��imlCЃ��Qb����OP���u�A�����.���,��4��T�hl7OY��a�#Ĵ7@����I^+M��0D_K�YC����~�p1�����D`
��ͺ�-|(��d�)C>~��w�=Lm
�o���+�1��N�e%c]Ӝ*i	�s��=m���δ�998Ѱ��qXj:w��+ד�B��s�h'B���	�Φ2ʪ�Ho^�����K��i6?Hy��D#h}���p"Ϟ���jA�?Tp� ��z�fN7��u�q��o	g:GHh*c������U�ɕ; �X�Z�)r�43�l�R��&L�a�
������`]A����T�w/�TTC�q
[T&ۚL�-W��<��m�Dѫi{1뻏a���Y�K\j�^喲�)�,���Fsg�c9���xhjšåD#]U
���%qs�����7��-���Ns˵<����z����?��+��JE֮SF�5����d������ź��S!e�C�7Z��J7D(VR*m�3��Uζ`�>��'�~@�����N&�o1q�'V�A_�j"�<�Z�(��>���
�Փ����j�e��`2;���v�(���W�c�0�a��/J~�H�s�hnxE�O�_�Bd['gwy�N���y�6M|e��J-"������4���ͺ����]�.<�!�?�*H�gT��A�_��M���8��c�h'�����w�Xi��݊��S���#~��X� D����!��[�8�Q.�w� +��N~7�p�s�2�z���4|&�ַXcVژ��>���?`՗!hC&̔^[8�Z�)�<��0~�;�D�^�4��}-���k��Sn2�j�+\���x�TWxgE���U��^��wj�����0�+I{?y����>R��E��X༓�Ĝ�{��N�Ok�!˶A�&)?�v�����)4�*�́��&��0>	����i�9.\Y6f�ݲ#Q�'���Ҿ PT��Cf�P���7)��A��EB��a��꾄uP%k0��� fV1��V�:�,�пnEE��n6�r{�v>�xa&�����W��_�@�ڈG-`��sNNc+����1���$>[i��7�����3$װ���4 �Eut�6��$fk��h���Tvb�c��;)d£�|o9��������y�Y��^�E*�$�ע�ס<��c��fè�[�G�G&�tEYxDɤ�&Q'FC�Lm�F�� h��<�)ƚ�a�v�ﮃU�� g�/�h�Z��0�4B�~ǒ�|w��v��7�G�3Z��ٶ�Sbu�6��%�q#�7� te�.�H,�b�IN
��J&���=*����L<��˿���9
I���\d���>��;���|�A���ɟQ9Lύ�]��a"����Ż��aZ{��u7�[�7�`b޾���Gʗe�I��m>n�m����Z��U�W����y��*"{V�0&����Ó����Ҧt���kÙݦ�@�����~=�V�oկ����i|��)hb�+z_Ku ��^d\W��L��BEG�*�$���4[�̸����P�W^����-w���d����?7���3zk�E��5�T���..���cӌ��S<@��54��CID^w,���ϩ�[�6�[S��G�6Ol]���tc��^�B���>��K]��)@�� �~�U�ِ��ݛ��1:���$U&��R�F�q{@I"Yg���}6D�rǠuL�,xs�=ۣˬa����b�7�c�9�9ȈT(�Ms��`u��� Y�ReH��2jbKTNu�^z$��-�.<������qv�Jv���c�<9���W#XeI�-�˓
�}�g"Z���)�eл �S���Rr��s���a"�)ݘG�d�榠����\�Ȇ���f�&�]��Y#�*O������s�
�R [Nںw��
t����j��\p|��B1�igb�LJ�g��w��%y.�N{-Z�˜������,���d��s\���*�Dk?A  ����<��9{���Cpƶ*G�t���!0�����85��d�
ǫ\`=ϓ������I��w��8�eΐ|�P�u;�K���^iஸ�_x (ǘ�K<Lo�2�!��5�-�!���`��J�OF�ds,�$:������#\�n �L+$>�U����M�|�����)�IǕqi���Ҧ�O��3��_�Y�l��x��������vFP���j
�4ɺ,�8�a�6�>������𖀥��际c��#1J��y���X
���x�+["7][rfr�����Q�ܺ��m'خ��12u>hus��{�O�k8��B�|���w�e�t7���s�U=�T����Z�iU	eC��cM�t�z����)G��'���%Nd%ҷX��l	�������c�m�(W����~��C�O�\9"%�w�iD�=*����>��T�V�^^����/����Ƿ������-R�g����ِ���1N
��-�V��CD�1w���㺈��{Ͽ��飍j!�: hE/B�� �"U������3����a�Z�9K��q�?BV���7��p/�}^�V����� O޼�"��Ι�/X�bm��u<T��/|�;�w^��L�:Ro�3X�����m �;.V�9j�/� ��	*��O�zgc���
�en��������ex�4�!Ǘ��~�c�.t�9�$��:K4Cp�#=��T]G��%�
d܈?���Y�C>�t��:D�SM����=AlYXx�J}�s!=�9��6<$H�hd_��-a:E��X㨽��tT�(��O��#�lܗԃ�ʊz3�P��G�,�L�d�K�M��u~����`�Z ́��ұ�_��@C�����m߂�������!�d*�ܠ���ۢ'8V�m-�����'V�4l��P��0���<���@AO��#��"^p�gV'�!��u�֮�f�(�J\v��PWa�g�M��8�M�!dv�vzO�&������}�4�^==��趭Á�%w]��$1FN���,�q�n߀��������S}y�G���ߙ�������k�C��ҷ�.�f�a���d2wH`H��f�e�G��K�ޒƆ����/��{�������	 ��������0h���u����0\i���%��m<�v��W�B� A�V[7��l�F&��F32��H<��H��e[�vr6��SC9�My������a��3�2��6&֪9OTڭ���SJ):�i�uL!`�BaL�b��5{o�u1�x�&%�Ufy��twÑ�o��+��fsE_���y���.�|�1�	����3����ө�������Dg/j5~.WL�O�=DI������ҕ|��y�&Ë�" |�em<��#A����Gr�|5V��Gz�`��<9�1訲�u�"�e�b���J�s�y�Tyx����t�"z(du�z?{�djR`��ء\v�|�Ȅ�����H��2'�ĕ�-ْ>Ev0���.���A	�qU�w՚�R�@��{mH�훽Iܖ+��9�Z�̑���8�1`���²�ߓ:vb��]�����\<�T�1�[�1��tY�ߦ�*�51+רF�P����Y�\�g���y����Z��ϖ*q�w��s�j�4�ɱn����4'$�$�h�5��!l�[�~��ޒ�a?!À��{)���x��Y%�Ȟ���=�T�����G���A�Tg���mGa�R�j�^��JJ��h��[?0��kP��c1�ҧ�9�d����֤A�(�^^V�&�7�5ʕk����A��>B��~��1<���̮/�c �h^�Q�m��0Y^QL%K�C8Y��r�S<4�y�;+��<Ų��v����P�T)�@���r�l�3?s���������N�_YOIpQɠJ˺\�S]���Z�3���b��J���Qnq=T=�bN4�O�k5ējF��0�J޵��X�~����ub��V�`دM4�QS[5E�b��0�2�>��O�r�n��;��Pm/5v:���T����mB~��eW��D}~sY��c�n��.����P�a%D�Ou�I��-0�Q��X�Ɯ�oE��T+m���Dx�J�]�{!�/�cT��[K�x��B��~�&(H��	���	�֘����(.��޻f�r�S%�#} u���!�fO�
�<���ȿ��KKp�ax{��>,3��̟[k�`�T���ԫw�-Д�k
Kt��),@x�X�6�\`m~�}{S��2�����R��\C:�����7���V��g��3�"����Rg�=![�wM��?:a���+�������$� ��~�}M�'�0�t�U���Q6�YB���g
0(�P�)�&�!'�P��'�}K��<5·TVA��\|��Tq���?�J��:�k�Z����cIY�C�W���z�i!��$��M# �C#���8e,�i0�7x���f@B�&��y�z�DyB�W`�����x�����
W ��+�䕔��ß; �o��w��%3-Kd���5�&��T�2�#iY�edUbV��w�����j2�v=�+�h[�/f)����]\s�#�K��O��vdw��9+��-7�{�Q*��̯Ç���/Hk��G���ӻC��3����M%�>��D�ұ�;C}�pê�5�)��� ��٧M���/'�F��E����M���~~�+arݭ[rd�	H���vVt���[�Z�|�6�Ƨm5��mZXbczX������5�'��2�E �����<3�'�*���WF}����N�b�����Z�UΜȕ̊P���m3u�vC˫�N�����N����o��R�����y����2����f�$N��9�]�� ��|�?������*&���^�s���wyy7X2�MN�B�]�Y5�u��Mn2�OI5��N1�(�\/b�/�v����nč���LF����ּ�*�d��ӌ#F�J.ЫUt�����MS�Z���o]I��˜�H4a�%/nN,�|��e��b����<Y���z��� r
���ɗ�\��V�h-���n0�K �F��W�d�ù�������P��}vc�����-�K�p��}��l��7z�Tv�A���if���j!(0~��X�	Ǻ� :@#8a<���Eb|#E���I2����R���ɸ빓�$5�����ʛD���xs-Ú�$��ب�lD�^��+�唺tAs&I͠3<�Mm�q��p�K�}���giۿ��dǅ	��5'��u��)���tR���*�Ɣ��/��:��O3+� ���;Zꪻ�R<I��b�ZH`���Bl�߁���]�TT�*4;���*Hx��\�I�c�iҶ�d�g�������w�wP��H����Z�jb��qF,z��Ϳj��������a��5s�+"҂�v�t�9�IqV����S�
�.�*5�N~�]����U&��*�U��=r��-#ͩ���EnV�V;ӫ�?�n`��>~#����4d)wV!✱��{��3w6v���nM��c�e�Z���(K�>�%^��)k�~P���4��;IK�&����U�ϲC�'��Ѧ+5rs�l��E���M��7rK1�Q�
|x���.y�J.Xj�(f��ґ�B;��q��m��a�ڄ�"gf�֕�0������s<`����}���+U��t���zK�*�#g�����̶�������҂FV�e�6�]��t���{��]x�N��O��{q|jH��3ۿ��=�w���D���	wTn9����%���l��mI�考�4�����%ފp/����`cƟ,�R�6�*$`�#~x�dw��b��&�8����n��^�+���{�c��T0¶��V����_jt�DX��}�
�6@��DR�X�L���0�iE�ퟸ�-�>0�,|Jۮa�����f��f�&"1��^h0��9m!�����L��y�_t��<<d�>�'j\~���ݙ�5�ܞ���>8��6�J�oNE~����34eI�%��6`w�( ����Y�<�Ap/gv��Wb��&���6<�B�F.՝G��	��[��i�z�G�X�2jׂ{#�1ṺW�+2(9PbHpLp;���&%�	hnG֪:�_l?�"f"��o_� �xM�44k?��l�1�KK�wT~�Z5yH#�^8X�ŷ�XH�j�\��d�1!a��Y���w<^X�AQ�ʅA%vZ�S_r7���u�h������vÚgFԠ�0��<��&)>��Э[-���k��c�v<�����ݜ��XD2@u@���n�Yp�����ŋ�w���e�*�ƫW���m����W��s�9�đ�Hw�� '$���/J�}�%�/Qh�_h���'!��	z}����\X=G����>6�$��֤�4BbNW�ى�D�n��KP����E�H�eKX4Ϟ�;�b�A$��'Xj4��"����u�"���k�J���w�X�R��ˇ���a��7�'XrA�>"�"��J��{ӶV�1zc}h���ȧ``x�T�p�+e�����`U�	��x�8�<v����F�Łu6Z.�+��O��&W��;�U0D(UB���\ϋr[���E�O,YmlF�g7�g�]� .Y}���,$X ��f���q��yû)���z��l�l���¹p�ｶ�[i������Mƿ5�ɔmu��xݻC>�z��b.Οz��J'��a<�ȭ5�υ���Ȏ�Ȟ%&���`���&�1�5�B�e�XHd�Q]����^��=P�2���c�cQO�������*�T)�c�-���+wO1�2#�LF�"�*���GD��S���A��lwz�ݎE�l83�f�!O�=$i[�sb�Dk�,d]E<@ȣ=�/�
n��k�i�e��P��b��+>�Hn<��@��#`�- c²��iu�B�F�kƳ!g'ŗ�����Mk!�s:Jڔ֝'�(,
�C6��g_�V8ȩ���$⤻�D��6�j|Mo\i�N�/���9q����Պ�`�v�{�Y�;[;J�RoG_OW��>&.wx�����ʷ3y�yRi�+S��;���D&���t��%���;&͚6��\e�}Y�;Zڨ����¿=�����ȿmܾ4zW�wh�/\%n��� 0r}���F��x�\,��ƕQyoϫز��}���R��܈�#�OY�\*蠻	ò�,toDe*�q������e�E,X~�xf"]P��g���-]8+�l�W\�p���0y��Ļ�,�H���;�!��:��/ ;��p��]B&j��O5&Ϻ@f�R]ї6x��i�a?������{?8��$
b��-h�BE�'���UG{ۺ�R_�O���o%��ἭA��-�i@ٛ�/ �
�9��zY�
yK�김�x�?)W����7�C/�o�Է]�m�G���q-3.W	]�HM0����c�p��t!`m��P��g����=�+24`Q��^�ءP���=�4 ��|��SS��\��sa~6e�Y��(u%�ܚ��(���̋�*�Ω>OP�����R���T�V�uڬ��Q¸�e�h���H�lJc"f,B���)S.1���IbƼ(H�{}��^��]��f��6K����ƌ���p|���id'/���H���p��m"�磺��*W �d�9������U2iC�N�5i%�8���$�8D۸3<$�2O��ew<����0`~�j��U�4K��I�"(W�9$�~ymmT�`�������+���)b@v���Mp] 0t�=±�t������*俖��}�$\z��V��z=x�
����_�[/m�r��X�? ���#��s5��#�,��@�?R?���Z��#�L���\[��Jߤ����_�����f�i���� �����ae?rL	1��YZ�E��*ݪ��*6��&�~6J`S�K�Kn%��1�*����q��v�B�R�	�� �#��)�B���POe��GgJ�H{��7*N�%OM
}���ߊ�Q],�?`���B�I}�f\m'�_��q�;���ϡ��. �-�FM���b�ש5��g�� %���F+'�J滿r�p=;t�~�Z����{���M���2#�B�ȎG!��Aͯ:����WV)�DS��?d8qs��1�nޅn�dF�Τ�ߣGՂ�o?�`w����r0ajs����q��w�}��M��#_*Z���gW��k$��1�y�Zzį��(x�e8d�fn�����<���=��\L��ƭ� 6�5�)�B�$�����]f�$0,j���b>�~�AjU����7�c����cx��ii�.L �HV��X6	�r��U
'��){Ze|��pZ��������������〼�p��*$�чDI��� .����7�C��dh�Ծ��R0���JxX!���L۷��-�`­[U�V30j�<�G,���h-����V{��4��YvҐ<$��j@�X��o��x�ҎgR��ƀG�K�J#Y����ɦ�!(1N�� w {n9E��^c�Ū&̍�"39�W"��rsQS{��儋%� A�g��)uɐ�Vx�k�q��3�E}nWI�.�fv��
BvO�����>-��G෻���*�V~�	G�v7�_�����r�1Yy�p�f�^�!�'�B���[�EH�1�H�C�J=�#a��|��LE
��ZH��S0�ԁ ��y�&�!GPݣJ�N�e�|A�����)�����S 4�jz�7�"���,�hy�G��p��妣YWLs[M�j7�]��Ũ�txdӧ�?���> /�$�@��y���f�Y���L�e��oQ�a<2��!���O��2S��p�?���������;��m�R\���^�h=_�:�M�zH�$\W�%a:>�4��g'7a�ϕ�ur��x%�6=�3���F5��m�0����%�lB�Բ`���͘I�!�����I�X�O��Iw]r���@W��l\�.'�Z/د^�Q'�Ҹ�*b=�"�B��|;�u�i�n>�1��:3��3�o�[��}�1cH%6"���=��'M������Cb�!Ғ�p���%PBX�xW�Ah<he�P���E��2��t�9�}E����H��Q��w�K�����*��-#O�Ò��mo���H|�iέA�.\��ϧ4���X_^���?Ğj�FI�t�xnG��Rҥ)�����1kq���\z�P`�0��z4��@��ױ��QN��lj<��':�iK�� �x?��ļ�I�ep{Z���/,��"�b���~Yyg�HɎD�L��ޏ"���W�3�?�6�ڝH��oS���������J5L{C��)��������f:`�2�x_4�/4���
Om��]�8�&�qlߍ'+���̝��|6�QL�S��eT'S��s-Pl%���w�n�����1��;t�[�U��9��^5�.T6,6�к*�W� �mx�!��}A�kw�]qDÇ	��J�� _�
BT�B@,�X��hx�$w)��ֽ�����`��&4�3�����S�d�=u��KKP6Z���flhL��JK�!nB.�UV��響���e�bڛ�I\ꖣuk��U���uI���p�v�v}Zv)q���@�i?������������5)ӚD������P�upe�H��T�9p�C]4�\y&.E�3n�ZP@�\������N>b��*?��U��جd����#}:�*<��+u#]��@jB�W��pc{BW�8�d/Y~�ᏺF�k��bs�\#��+p41�f�Z�tZ�?�+c�Ә֗#��k��3�]��s��K�S�s���y<&�ǖ	��ȕ�A33�S����=�J��0c!,w��qb�N�2T4�yp47沉l�$��[��z���6 q:�PF
߶���|�����N ">��	
�e�*��jΘ��֣֜�WA�#o�6�1����W�����q�X�R���9`d+Vw��!S
Ǝn��M}�v�ȇ>:X��JhS��br��K �Ѳ�<�T���R�i�+?P��k	��Oe[I�P�Nr��T�)%�v�s��c��~���K�ү�_���zs�G	j=�	�G��S�Sw�eG�."^z�:n{@��E�W"��Ӂ�41�ev��@~|�ߗ�4���.�a�x|��%S��mD� �m��(���R
�K:�ۼ��-��*#5 ���a��_�d2|��:lU�kp�hp
5�C ��-�,�|e�WNy�s˖0'�6�`����i�L�q��_v����$��V�q?�S G���4�'��z0�ng�A��M&1�F����]�����E�(ۢhT�.�*t<�B�����u/��rR�W�,r��(��l�
3���7D����-��n��4gl�ֆ��n�]٠��rB�[�1,�ￛ).�N������Ϗ��IZ�� __{�6��/����11�d�m�n��hM^k��*ݘ�[C�
������������`�*V�V�뭑��a�vg̞x9\>۳����!8<�4I�^	g' )j�:N*B|�6b�^��|�;�@�4�o���n����E���("Km ��/O��_)��HK�T���Ɛ���SG:I �$��!	��uy	ܠ3f�� ~�E#,Ht@���ߟ��e�S��v@;&�z���s�b W�jR{2�%Jv�E�l���}��v�j�a��̏8�Vdn��k�MjX5�s��RV�C�-��-U.�𘣧3�$$ 8��P��܁�d��b�hRJ������-�d�(r�Z�̥�os?ʱ��̼�}����������.3�Mq��ǂ�ag�Z}��`��rg��Y�87�|��<�2�	�> DYS�C�r	����@	zҪ@�qʢ���d�΅��ߔЕYˣ�߄�j�V�fe9%�ݪ�8��Ǻ
@(��U?L*�|F��F���s���J��7a�I$9��y��W|pHzs� ��_%K�dU��}�1L�fT�����.Q =����U�K�ϲ�7a�FS�>?_|��4��[�1���M s�D8�>���G�W`�-'M�I�(F�����DąٛT)��������K���>G��O"�3�lI�K��ԡ-�@��1N=l�2���ňW~M�	L�OT� ��i��nmjR�+���eԵ�c��G���^���b/p�w~k�b��U�,š[�3'�C����$��z���$m͈�G����}4j[��M�W�	�i�Y~��e�r՛1b�X�C���P>9�0l�n�	F,��ħz���zed�5DTZy���uxov�`����}�΋�.�������f�����%f�<��J���8W�3�T�J�_o~��0l�c-��E#�g�/�T��o�s~��u�&҂K����P��O��~6�����f�Ǥ�yO��M�ĈL~ʇs!��ً
��z�ό����bT/�6��fZ��K��N��K&>2<���p��3�T7�Q]j ��Hh�����F�kV�)�iQ�i�~��P����%��<Dco<��3�O��E�,'.J,�e4T�D��j���]ĵƳ����u׳π
��!�p�M���r&��� li�!����+�D_.+���!��������'4L���Q���r�A��Sa�p�Wb��c�c�4����Cr�
.�*���,�,�p7�P����~ �i���ݲ'ˢ�v��ځV��2&7�J���R󗶛$��'�*#�!=9���8^W���FL�Ĳ����S�M3@m�e/����ue��j����]��	]�@	`s�B"��#?��v:��������^�8.Z���b�A���,�O�eh~��i"�aV��X�2�?!ǗS�ƀ�uV�Qi�73��c��H��!v*'&���W�z�>�(MZ����\;�$�vr*"A��#�}�G�p����2��k���|Z�s	 b�Ӛ��.A#����=e�8���$��x��l�-�p*�F���Ҽ߮pR�� ̔W��,d���^C!���	���;d��,����N���yq	��>1�3<�w`oD��*M���N�:������ޟ�	(7�^���qn�����v_���P�iи�fKz���̕��KR]�vc�&k��KNc}i��L��P����M>��A��cpҝi�p�?����\�3�\�6�F�<����>7I�&������K��}�/�"7�����i����1vE
�d��eo� (�k5Մh뀽��
�M|0�^����ޮ�a( ���	3Ϣ6�LR����@��C}����uڞ�F�c+�[�}�Q/��o8�c�'Ѥ��8�?]ûcL���H� �b�<#9\+B�k�zT�Y�q�j��kԕ�"4�(����|�����Iƕ����ᪧ�~�o���ֱ�b5��j9W"�9��,~:Y��<�-�e��<RP>P�_��&@L�Vl����7
�9w�5������#5b���EN8�F��t.�b�����f#�1S�v�Ӣ��P]����QY�(t29�eC~�m\D���4�l�-a�w,��3��u�Ġ�vE���2c�� F�9�D��Ag����ꪽ+�G%|M̙V�#�t�d�PL��-�L��!d���}��� ��8�sTǳ��H�$��M�ݕ0���.{~��W�O���.���ߓ5(|���OT��(	N�ڵ�-���1a�����"�/���=�P��ƙ^ZF�r�b��O��0O2(S��E܊���Ib ���pd@�	s��=��%�0F޺�[n�N2d)��3���m���ktP_H������Ĭ	xDck|tK���8��=?�v�H�[�}W�	�[��CcA�ӗ�:u͟x����(sa�;�=V_-*�-,��N�$��Nn��,����U�r�-fH�c[���J���pz�M�*a���K�j�(�߇�p��j���_7Y�%Y��q�_�8�i�e3�)�ݍ4 �(�d�ǒ{q�h����N;��g>ٗk��6� �<1J���Ẅ��aFS�q�H9d-c�����ª,#)*�E_Q�x���pn{�<{���.>�v!C�W_�g!tH�p��H�,�O'��wQ&3��Ѭ�1g.���挃#�Xv=��̳u(��������h��Un��V��O�T�v�ړ���8듎шoG�RV
��A!Oө�sHM@|�z���|J�wꑢ�IߺiV*��鸲c;t��\�C�/!vK-М��'�������ue#>Ok��MI�e�i�h��}ě@h�軾����H��Z&j�V�UN��I�@g<P�0>o��kdX��ʛ'�s�v�|��b�����p��	%i�5HyKI�5b-�	�Kc�|dKj{k� |���cj�m��U�b���6���ot��=K���/��&��974BN$ԡ����`��ƚo��)!�`�����"���i?�%��R�;��N坳H2AF5��1�@��Î ��sĽ���.nN��:5#��G_h(�no�pz�1J3����G�j}��t6����7�jx[�L�Z�,�V���s��LŪ#a]p��e<`ߋe0�������2~��9������"=�4,CiIa�TH�^I�k�8w�x�����K�<!���}�ʂ��l��إ��d�Q�MV�7��8v� �ׅ=�kNJ�,�H?�݊���׵:@U���G�X�VD�����s��G���d$��<����1f ��Q��(HQ�O�C>�-Y��:7J�����5m��fg�v�,�Y��_�b�ID��L�dM��N��p%���7V����P����},��=��������Z��J1��w,*lz={�bc��=��L(�L�͢�9�5@�F��a���%��W{�~>�l�f�vT�����=�2kY�Xe7��9���p��sg4��4���̍��}��e����+�wyi��{���{���~�Kr��v8GY��'���KoId[�).�I2�T�=W��A������n=F���Ʋ��g��2b������]d�����8O���g�^Y����֊*��_���pd1�������TI�ô���I6�����x�֫~������H�)�"B��W�IN�!Y�}�P�?���R�-���x��QC����{�o;{���S��Q��>+�=�{u��	�m�l�S�F���m����+]`�{~g��?����"����h���k(3�G�	b�\%QV&#�t5`T�V�P�ΰ���=��Z���}o�KN/����ro���'��x����hu����z0,�#��r��|�i�SĄ��-�G�^ش��[��tw���d�7����߫������ڔo)6�f*���m�����m~�=Vh���a��G�꽰���z�"kAj��.L��r\�iVr��K\�p��ɶghۍ3n�t0XG5��Y�^u[�UU���%)���ԗ�>�gqКi����Eo�h�l��!j#�%��~�Hh
����V�NkCF�C� E���!C��׮��*t��\P���Jq8��$��u-�9�8�=�$���0��#�I�*�SB��Wl�[S}�Jx��G�9Ê��p��Վƨ&���{�u��RE�JM0HOٛ�,UY)� �/�9>p���L(�Q�a�v�P��g�kV�.7�Nd?ښ�Jv1��-t�#�;bȰQq�+���pe����Y��A~�RcޅM���.�̣Om5���m���&�p�� �(J��6�3	FI �(�\{������*�Dk^0�5��nǿm�÷�j�Ur"MҊa�����NX|O9<�aj4p����`E�~W6�;h�^���DN�k~>Cc\���&_���V�OӺ*�}��+d#��=g҅��Qc�����i�l{���b�����J�����O���~�y��"�,����e�&̓�ƑV㻱�KL��qQ ��ш4y��~�$��"�-�!���6�S|�n5�&���~8�N�]��1��
M��n�O���qt|���X����2�|���S�\��-۸�;��
G�P-����P�ޏ��a%٣)GiE9P��ձ�>����d�(!��/�[�)���?�y���1i ��u��kK���An��T���f�����^9�!_O7�u��A�����WeW�pr��� 7�{I��?29�4tX|@q��-ٗm�����&NzJ:��f@��mH
�\��Z��)/�{H�>8��g�2�̧����H����}�������l�g<w���-�2�3�<�����e)6 �5�J���~m���*��}|��I)��O��)��?5���%���_��{�+A5zR��g��_��羪�*���O(��AQ2@T��F��{�gD��(��$��]�����}��;��V�SE�Ӝvl�&Q�կs��/�r��Z�S�f��(D����CGU��C_����O^�5.����o�
ݐ>�nx�Z~N�I�"G�`֬UK13"����#U�	EW�>�_��g���T���x�l>���D��-�m�J"�߱�eJh��"jUC�nt���9���d)e7ߊ��6x
�୹����TLB{��Q��1��j2©�C��33~>a/Y�����"���ɣw��H�E�V��^���^�7*]j� ��(��{��ȁ�Dd���|�e6S�b=���x�j,��,�݁��F��+�b���5uy=x��j�IRn�X�1H��i��_/�y 8>��b�e�jU��8e���5��܀����leT�m2h�]��F(z������1z��̢i>�~��?�|�|����S��i�P9TC3��Jmʕ�AZ��@�7l"�q��۷s*��e�d�:2=㸝�AC3����G�9���Rm�P��ી�Kf�o�Uh��M���<�U��� �5*-�C�f��Ð��6��	%��eweƐRo�<�1^���(ֻ3��(>q���i��`����@�$�[��
����=%Kj,�x�%�e_h 8=�2.H9�&7iӾ��|]�)���f���-(:�F�q��G�Q�-�z6�hd�c�Z����T�s�G�hH��k�sYg�<+�s�5D+��8fZc1��ĸ,���}��O�Ʃ�J�[#����G����لE�F�zz8M��^w.�ve)�YH�b�;�0�t�JVq���9k�M2ˈ s����qN������n������BK���X�_b��� ?�"ῌ�^'a#y΋���\B̶8.�H�� sb�:�k��	$"��aT̆���ÍBسnE�a�ډ8�xG�n��ߏ�ޚ2ʕ0����|�Z�b�����C�d�oR�D@�l��}��֓f�!�_�(�ޛ�[~7��z�D�Ag*�y_�����<�5_�OP���L,�e�1eGE�u�Qu���{��A=�c�	1_(4��B~��R���X;s[>B���ȴ��.xe��҄V�T��,���#�sO͙�Z�ۀ�&���������"�S��p���Z|�`�Z_N?�\�^���]�'�%����ɖ�1�>�ÿ�+�mq�?7�������˘ �)ۻ�jz������h�~��@L�
����D��K��-ٽ��@S(�(M��I_G��bfN���@���z��=�Be�O�߼�B���P���i��ȝU��	������L�LCV�2&���cB(��W��|Ӹȣ	7���ŷ9�%l���`WoG��'�A�P����\OҲ���5���Xa�*3.p���� ��G����)�<2���� ���3���-����\�Sf�m@��O�I4�*�Z�ǋ�ƒ�?�ytz���."I�ƀsTk���v~o]S�H�����������hO0٫%u)9�C�</�Z)������D:�c@��vy��\�b�)\�]RF�^vf��̹<�!��c�^.��YuV	�f�̗ �l���4.�ϰv���-��.#���g�e���Ѐޒ-ъ�1�2�d̯�3��^��Z'R�{'�?����ʊ��c
��`���o0r�Η�IV�3c�XZ��^�f
�y����e��߼�\��<+��t}2��C��.8�;���Yz��B�18��.��L�Gʀ���������BĀ6,��j�:3ckr��՜iҧ	���.�����ҟA
����;�h��f�!�wwg�}J%.��M��h��ɲbҙZ`?�c G^e���Ӳ��xK@�S�
�P�<�`��Bظ�E����n!xk� Aѹ�b��WR�8E|��w�YS�,���!��6XE��"�U1~[�#��=֌�>=Z�Ӝ�nnI�\B^��0g�L-��j�Q8z����:<�=�2#�~a�l����ڤ��Ob
[ۊ4�4�z*K��c�8Vk�菙�	��ot�}����5�I%�M��E�,�'�y
��[Ӝ[љV����m�?Ha��B����^����\���7���E`���~������T��;%��lw}j%� f'�WI�\�J?��(���i;c)����N��
M��� "��^��(� H�F;%/[�}O`�˭��Rމ���Zӕ�t&nz���S�%�rB��ލ��Vl9'!������o��8�:3/�6G]�^���ō�j�b@�_��!O��yM�,�C$���h���<K�I,�H��L>l�_`��$���)s�K�ʄ�b{�z0A#���W�M���'�̼�H��I�u�z�?@{�>�<0�|�Ŭ�nˑ���K�$������Ts�c��.Ԯ��W���>b(J���q��Fpk�f% �J#��'+n�1�d_��a���7<��o�<e:㍄��ԗ�͢h7&c���UtF��f��j��s�[���Z3񻍽{,���CЊ.%� Vm�o�X*��j�B����h�m�qB�IL����:D@��K��q�N��p٩��j4Xc[�)��-;�}f�����Zmw��U����~����L�y��Q��z&���T:{MJgA���ڼ��}�]�ц������nR��p�E��!�Ռ�(N�T�*��,�Y���SS�>E:�/�!�E�l�K�5	��_UA�����r7̱qw�N�+��L1�Ͻ,D,��hj�j�Y��=�KIAh�]\�z�U4���.���T~k|"�3R��5���s����#�/O���#���SD��K�����~�F�d�Rt��ȷ�*�J�o�U��ߔF�h4����B^_�P�]ŭx[�ܫp�,()��g���;���|�]�»����8Aܼ�ƅ�E��+�����ӳt�;����������$PϰT�����j�(���{#�#���a㿗�I?$�d`8auS;��e��K��|+�
���\,�:��۠}�BT������@Ա�q�ٷ�&���8q���ٹL�o���9$��!�۬������}�mnNߘ������,ϔ!��p�0��G$�A�`�Η�_!m.��#�Φ�/g�CE!��xמnр�S~�i�\U^���߅�ʨ��c��+S}�E�,3!XgLM�xe����tp%�SK����,E��=cO�j��uY�C��c�x�`�p����+�|��8��"Y��~���'�+��(_�0%3_�Sڃ�����}'�t(�0���ɸ�MkB�}�
jI�]+��)"�K�ן[���S��]{�4)��#�5=��&6{ܫM��VBQ<Q�9�]>��x"-���v����+_���"P}��,e����yB��~֠i�b��Í���?���m�g,I�Nn�;�^���ߪ\7�0��3g��Hmո��8*>��21��]�ߪ���`����=��� �@kk-�d�VRs���}R�"\x��{���?h
{yυi@�Q��t۳x*�M@;yX���=���'���:�
��y鮑�0�ҧrnJ���x�rRTyO��tl;��_�gh�g�p�=�Ka�E�6�V���p�c��^U	�}�׊���/�C�C�_˭��t�g&�J�U��y61�K��Z���4hVu]��ho�=p��M!R�����XG��nYtD��Pp̲Q�������P_Ђ�bD�)�]���J�Q#f�ޱ�Dc�BI���w,0��5 �:\HA.�K ]�JZK�@��.&$�D~�D��l�~��1����PŞ���u�r�V}�V��<Q�N��6�W�[���W� r۠�n�ԤZ�7Ux�S����~&m&��ϊ��9���'�d�_W�[YP�$������	z)��fM�|��d��d��8sM�Nj���״2ڕa!��;��;k���R�R�̃��]�ҿd��yv�	��\WI� ��Q��l�S��D:���`�?w�x��Q��o�0ܰ�l�慹��m[�;�j�n��p��M����Sc�:&~s��ע�U�_��	��m��k��U�;��g��U���=��(N�����5���i�$��S �rLb��3�s���Φ"�u�kY�K����I�431 (�ٝ(�
 7�ށ+x��P`4^m�T�)��;�d攪�X�M3xε�]�2���:��(f$3��f�z�phkE/tB�e�}�p�^�d|vU���z�����������_��S��l���|j5O ����$Y�Ԭ3��<s�1��rx�yN�eϖ\ɘuk�_��=lFM�vh��}{`��E,�#�O[�6/o�P
|���%�I;�����%���5��p�x�P�1����i�?ިS_"!���j��� 0��Mv �Y�e��xd�/9
ɑ(�6��;:��+K��U����1X )�ɪ��ML]����@�0��ߕ1�s��b&��S0D��{ЈĹCJ��3Qp��%���;Z{s���2��j��wͰlE�NW[���Ô{�M��iv�O(Y9�-�����X���s%+[R��g�S��� &6�KM�r����W]Ld�t*Bd�AY4"9�j���a"<����7w�''�����k�.{��5����d���G}�����h�ٴ� �w����dg?Tkq�qC~�F?���뻦��D�y���yt?�o����?NUH�}R��c�F��O�,���0����lY��u���_�p+x�I��>���(B�g���,ӏk$�#L�B������A��8-Mz_��uv��
܀W����<����Jtb}|тh,]�9b���d�r��V
�����X �����ǢRK\�������}�7�gQ����%�*��O�5,�l�H�M�5a(|�1Į,�\�i�I��,�=�7�iB1��@)V�g4��x�%�c��/�^�f{x�T9�IKP��Q�܋eR���m@��� ɧ��OoM�s�O����yQ���Uׇ�Ո�\�,S���!���D_��7M�PGj �,y=>�����U�����|�Վ���8��K"�h6���_�%������s&����� Dw� o%�O����t=Y��Q��o\R�����7���g9;<b�꠲���L�J�b������)���C�� � >wl�x�```ȷ�������"
�<q��qOb^��|� 2���G�GT6�	�S�jNGX�[�B�o�q�1zH�b\��xA��"�I{�Z0�����RQ�	/�-���n�l4�.D��A��п@�Ǯ�YQ�]�2��Y�g|�;�?�+?N��领̕[@���s<����DM0z�P���v(�3�	%p/g2؋��&a+8ʸӦ��@����'1&W�=\���;%��5�H�C?/��X�Hӛ�ܿ �>�/T�T�n�fͷ��Ã���K- 4H)�K�s�Q+!�Ը%4&mt�^�DG�5�ac����8x�U%JHH���	(S��鯧�φJ�+�be���ҍEp9�7�в�ޯRU���#�d ���N}���O�Y
|�A�Ǎ�ѳ��ju�ApA��Oh��m�kXh�$J��#u�ǗP�=@PFb/#�=H��mj:�'�du`��(���j5���������j�X����n�J���3G��N`�̫u���h��W���A^wl��'��F���Vj�(��Ԃ�1�X��[�]��>�Rd�ζ=�)c2	�`7�S���V�B���ç&��}��W�Y�,K)�ݣG�Z+1�z)~�nt��| �d(�{�.N(�����ӣ��겗)	�2Ać#��CH��yP��i0��'&��`�Y�h^c8�T�V	rp��]������̟A��F��Y��X�h)���B^�{�w�%�fy���} ��_Dɓ+��O�W�6��]����g�=��@�Y��]�6uwq��͒���x���­��G��|E�yI>e�	�oc{<�ZV��2�c��EY��)U�Jm.i��"���X},���:�>��(��(-����o:'����n�w�ͺ,���:(�����l7���!|Q�{��nʙ�x�"�t�8��4���@oQZ3�K@Q؃�����!i8Gj�o{џL� 8��"�҉��6h�,��e�0�R�f�� �P��2�_���el.�6��Y�������G*�IEVy��B�Y� K+_�i�ԑ����&�!��I}�������'.6�q��\h�> �E��]�n�9�0
�k��u�"��V�(Hϵ���tl2��,>#ۛ?��h�[���ð9���Z���UJyfyʶ��z�ǋL�>��ތ;��C�-~/n�Q%�K�dS!�S坯_V��+)�x'Z t'�(߸�ܻ6��m2�3*q�Zk��)�Ƭ�*��%�֜�w�@��zUY�`�Q���,�n�1�o��5�K|��A�`-���-��G�è��$͵⍔���$)ӎ0c;�=��f(�b����PuI����$��'�����pWr���`����q�#!��4����Im++n�4Z���PB���#��p��|q�pY��Tf��;��3��!�1r�$|�9�������b��_��:e�1%�?����*�3Ǖ�L��^E��S7\�Ƴ5&�"H]{(X4;z۱�[�;�\�j�S-r�+�y�3��u�r�*��B�A2��K�|2��Q��.�ȫ2c�$�22�w��W�����{���ΧC:��xǭ����	�9��V7��KH����п�]�Y������d1�9æC����yX�R*bS��4��|Uwz�͏�"±'	7X	�A�������~q� �SK�r�Z|�c�b� 5:{��Ӷ�/ P{�����ٸj;�qkF)�Xt҉I����>d�Ra���9�f��)#?�.j#��%��u/�U�%�4�(��nU����������0���`-,DSאyvؘR=p�!Z���	�o�uc8*��=�ja�gmh���Y�)���8�1O4��ϛ�-(���x�ʋ����JX��C/OV�0Q�8�M�	��r-w��`����K��c` R�^�������eJ�|d��k�q ��cb��8!B��t?�����
*�W'��,�լla�P���e�q}ML�1�+���)���_�2%9�C���t�0�BUF��"i᧋��a�jh~�;�؏��n'c'B�imR��97tۨ��)�붑���tR-$A�{�A^�.�X��D���c�; �a�c���&:y<�)YN�(�ip��rjQ9��LKSՁ|�K(o���Qi<�ފ����(>�Co��v�������-��("��݊f��ȭ&RY�̌5N��YM����4x����
P ��-�g��eD�����3�R����ƗҐ���NA.Ip؁=ӓ�!<΍aO����?��K�,�LV���Rb L�^:ҁ�MIy���0n���7:s��p�ڜ�E��8t i����e#y�}�B�5��s�0�/��Z����//f�?�k�#�E���4�W��NjO�)w�5bD� >�J+�CR����ܭ������B�>%:=[�M�%�c�.�3����ټ;y�9����g*��K�[*vh�a@\�Nw�.�k��������g�{H��L/����hV�
4��?F����Di��5	�� ����;��QoUȳzd��UMN��P�1��cT�L�b+�Y[��)wj���0aN�ׅ����\�Ke����[�Y�';�����V�s��KQS�_n]_�k��It��p.!c,��7��F�Y�ڮl-\��Oz��r�(D�''�C��.wicl8Eǈ���В�����I��t��`�v}p.���n
Ap�q	��&����{�*6UR2��P������f�X�7i)nJ�P�fA8�P��T. } ӑ���QY�bT�����4�������V?�[c�"�\���y�e�q5������6�t�{y?�JMT���hG���
z�����-��F��&"�W<����e����VN��߹1�5�'͚Z�!t��BT�qW{r�I�����;}lQw�����
���`�� �~�@R�<�9��[��K��xߺ�G�H�����6��M.���$#,����$w��	lUF:)Kc��t��Cgo�>�������=�����dg���އz#�>��yI5�#��լ����B�t�z[�P�?�K�T�����r�����D����m�Vyɒ\�c�?�Ύ����,�h��8uv	�,�gIZ>��J_�>8�&�w{+ �y���'m�.z� �FAŚ��q�^-[^fd��V`HUL.E�h�Ar�=����f|*O�Ƽh�8�>�+, /=�_�Vb��\�����������l}N�ُ�+"I+�*��t�d���=_��|�q�����*B��Zfj�l��P��
GH��?�~9����Ԣx�۳�v�� k�epl��H�w�Py�Z�ǇO�Q��;22v���	�ES �ג�w [6�IegA�K���r�Ҍa=���nӻ�&�!�|uHo�q0���yj�S�6�����-�"�wzE$��$���Q��T�	���i�%���dJ��?� ESk�^x^I��g�ɤ���5툇������J���j����6Y�{�wm7��Go��?Aou�e1Q�@�Y�w,�n^�zBA%�աuT�N����"ɍ���;FN�X��d�o] "�@I��}���2�(��8��
iY�L�wQ!=�d�h,��]2�I��*�W����'K����9��ꝲ@����@6�1�R�C�Wp+�����p�gI��+��R�^n�Dъ�T4*�`�8�	h��ě���@����0:e���w:A��v+Y|��0�-�-3�Ywe`_�w�'�/.IĘ#8!�s:�o��fnd.��& ��t�S��xD|�/̃Ž[� ��J�KX����1�C;L'8;�;�qS����jNR�|�Z~-��L�D�8���%����R��ܹ>��<�w����)Y�ыl^�^�^�#�H���t�V�����W_x������W[b��j➳�" xi���.�q1��s��v���|���V��b�����-�W�}G�h��`��$�y4��գ���d
��1��cQ�@@��R��h9�a5��)ɏ3d��Y�u��J��ɛ�Fl-�߁����41h)uL��.z�C3��t�8e�cq�slțu�y�
�?��quGԹQ}bp2��1h��/� 	�4h��p�:�>?��ٯ�W���'~,� �^Jסּ����\KU&��hH9�k}��\#�!��k3kmd��W
��ꫜ$�F[)�x��}5T]�N
�3�6�3���-�t�{�E~�9����-���er؋���<�4\|��G�~�9ן�����}�h�l�رp��͉�pƤ�5�E�qA�3�CX��� ܦ�X�!'"���ez�C�v/@�A%�D����=�B�wף>�E�e�OY��I�$I���,X�1]�BU�R�+2�� pK7�NY�-�_��b ��u��5A�����P�m�=�x[8ݬPV��z�����߄��|R�M�(�>�j�k��=�҅a)[��p��*��I���P�*〉[�II�g�b횊th�{j�w��<LRm��f�w�e����Y�&5����Gd[ ���偒L�
���NiS�a���!y�ͱ:mt"+��IC��AJ���ܫ��G(q�dhW�.>����sp����i��5m���Q�o������aD�Ә�Z_��{�	E�! a����(�U��&��x��8'�O23n����r&Y�7�|.'$���@/*:sCG]�l�XG��q� 1����S#��a���m��d0��Ș���"?�i��NqgoC�$�o|�8g����o����է�AR�Oh��0'���5��\���_�Q�Y�p=gq�̈́@���͹ʹc���#wXMm��\�r�/U|��"������K҃mչ��� �9�jc���'ӭ��h�n$��! aH�V�)ޗ�x�����ż4��~9�W%�[�3�򛕏a��K@�y���W��eq��$�d�������^o���B��LU1_�(j�x�B�Uq+ym����^h�m�F�ބ`�9p?H�j�b������F���9k�H�I�$�Y��ރ8E��}��,#��ש^���m��ux|UQB�w~�S���AtYo0�ޅ����o1{�$���\Sjb3�ȽZEg�P�a\��Q]����/=��i�$G5��+�'M�oS2!���ɵ[��p��BШs<�ɓ�0>m����g��_pc�-�`����MSO�O��	B�M1���[��n1��'��F�6(K���vq�:�mfӖ�YK���FS�����	��2:󽿴U�������CN)�96g�i�D������i�lF7�҄j�¿��ɥp� S�Ϟ�9R�D�&<�lU�0�|�ևN҆T������}!Uj�W4��S�m�He��j�h*[{������p�̈́>���M��V�� �Y�fA�81w�,0�e�� ��d���W���7���u�R;���1Py z$b�!�P�m
=H��md��),lƕ}b#0?׸�ڷS9���v����R��k�CZaǻ�R�"���L@�Go5+����ϒ�@V��<�/.�V!�m���.�)���'ojڄ�!���6���a50�i�
n<�J�̯�/P�~ ����Js�o��*�xL�m�*]��e:��-~�D���_:T�;TO�!+&�5�5zL�L���'Z�wO���9���х�]�� ^�rÅ@K��&RWgt����eM\\�ȑ`�T<E�"�����V���xy����Ov]&b(�!ATA	Y��+jx*>.p�Ea��a;�Ʈt�Cy�!�g��0Ԫ׻��C�zӴ�����L��_G-�?�q��"��a��8t;��Ԋ�����lHi,f���z��a��	��9ڼ U���C��)zf�Z��=�;y5�}�3"oi��*y�и��@��4�v;H(3���m�X�Z�������k�����K~Λ�LX`�����>?y�����ߋW�qHm��9�?8�'MP��]% !O�b6���"�6��q�)�����P|������hɂB^6�}������Dꨗӥ�Ԏ�H\�9��Y�c�?�x*�Ӗ��Lc�K���\l �5��8Ͽ *���Ĝ��{���2�6D-��6�����E�b�1 ���vd((٥�2��z� ��*�\�y_����tH�C�=q�S�=�z�,��Ԅ��������Hv�V?%����x0_g3�ȩً��a�3�D�Ð!U�I#	Ǥ����T+I����m��0G�[�QM��	�_ҊK�{yPЦB,�r1߁N�pDI(3Z�e׈����y2��;mS�����L:\7Ύ���G�w���_��,�"Q}��[�f��VC��ES��,�#|��8�u	�}L�e��ͨ�g�(�;>�<"�gI0�móF0�p��x�1�T��i����a���i�s,�zH����s�a�@���a�Zo���s�3q4~�?��?Y�[�����8f���:��gP����m��.	D���kyu�(,��K����a����k�8���־����DV;�w��l�/g�˶u?����$���B���ٖ��E���>E��o�mG�d�	�˿вQ�UkC� ra�8�#�qEy������1�i&'��K颏Te'��#�ƅ~��o]tMe��3�V6�>��voQ����R�q�6�W�)��Z��Oܒ)}�J�"Fn�8�1̨��UD���B+������ӝ�dy���6>.��&O~��Z�k�Z|��D�`b(�U&Ϻ�g��U�@���1{��iyB[�y=N�������L]9��uύ��L,��/�:�j,T�D����?��� 	������#x�"������4M�$�¨�j�2��6�By���� �Ā����gm�(@�4����DU@�:V�=�&!5qׁ�`!6�wQ�1ҥ��/�`���l�4��n��T�-��~7�L�U�>3��b�Dd�����A�W��s�j=�	k��
�����u��И���>5�*��t�N��O�n[ЙWe�=�B@[��V��:���t��?v�#/�+����;-)jx��Jq�)B�''t�\ӓ(��ی\����VĶ��r5�G�򏞲�K�)Fް��˷�B�X/NF�n�gs�1D��v�U�x��j�+��ۆg]�kQ��`��P��*��/�����06&�w�t�n"'�D���f�a�P��69�P��g�[NNG���}���x�����w���-4�3�|?aY�bm
�>��-�m2X�@�@�d"���2پ)m#L�8|I���rs�+:� ֕+5Cz;IR����-��
�"O�b"t #l�;��ou�W�M��_�
ڷ��?��
��	B�VF{�r-�$�f�#3`�q���~X���
/��~p½��w(���;ϰ�R���c�6�.�F)��k\�r<|j,N��d�h�^=�u)�^���z��*l&�+��{*~2���{'�\���>��V���)��Z�,��PJ�}Z�ʾ��<�u�i�ق��|� �a�����6S��(nNwѶ��bwW��˵��mr� ��/�4��ۙ �L��F�{��
�}]`��|S�qx�!��й��:,!$���"�U��k��(�F���<�� �y�SDh�Y��k�����e��7Z��w�����Ә�	Yu�?�h~�����9��*��t�]�A5O �w��%zf�����"nL	~�|���y����	RF�3WG�?���E�>�0؅�oEJo�ᛮ�*��kbR�l���S���[Dͩo�{j�EA�א�NAc-P��ݶ`���\�nΨN���Y��C���a��$��N9G���piG�@W'I��jB���#�i�D@s�������T�j��M�Dp���	��|1#Y��9C�Ҫ�oÀ��I�(�PH9��FC�I`�YP����3��Ҕ]��m��:��s\q��?���(��I�O��[�m�U���Sg���#�2F��+;����	�z��#K�#mCp���>ITiw}�q%jn;�7[ܕw��_��*�a�P�Cڸ���P���!@���
�R'�����XV�χ2����8�J��RB������s��1�<�	�`�{��/M�|l�7��W��QOq�HI;5ur���p����A�9ivS<�G#¸��Wp+��$p�������O���C�2TO����<�8�H1jы<��Q�0<_5�c�Q-N�o/�4|t�&n��.F�
3�Qu��DXfFvD^%k��CM���ރĒe9[��@�2̧�V�&W-�h7�,=��MH�@�D�u�>0��D[��ftO���IZ뚦uI�L��:�1ʋs�P+q��M�;P�_�¸C ���~��%���G����l�:L
L��P�3���R�nr�T��K�� E����_x��ei:
�[E���&��`W	�Bv��ߌ���8��2��?�)�:"���/Z�2��=�+#sy*p����Q(��m���Nl6nr�Z�7<taƽ�%ɛ�k��$�c����n��g�t�+{7ewk�����
��r��P�#'ޭw9L��Ob�bH�;H6�܁�x7���#9�%�`Ԙ�Y}�Q<�NA�(�K�t�J��^�
�>�a�]����D�9�j�l��H�+�K 8´�|2Yp`�@++�p"�����ժ�X�{-�	���/4*���c�獜ɿzRގ�`��㚶��)���e̻�qU90/քR>.x^G=m��Y4�{��Á�ݧ�9��_KZh�P`��w��ѲN��"M�ǰj䗟&D���H�S��~�7��>���՚
k����P��s��_�-����:��a=�_���r���@��y�e�S�W�4�Ƭ�]�������C�nN(�C�m�Ѡ����vy"�:.f�Ǳw�)[�����na�QΉ�.j����O���OIr��z�$d� �o��݈/��l���]k��/�U&��s}۫��7AL�֧��n�3'Z�q���ru�����ϫ�g��w�DK�zz�ğ,;�;Z�%�#�+�#�=|�C/�����!w�JxRv	�/<)N#�Z��7���;��;O x�**̪���6g�3�����lJC���D���`O�|�)s"*�%�l=�P�����2C�ˬ���#�����-���D<���te��BT� }F����ڻ9Y���O�Q̣h�-h�-0�6v��M�בּ���ơĊ�I;��6��y�5 �pK�i����7���:�Ӟ9�ǎ�v�&��.X��+'T�|��8^�QG3�v���=gsyV`=
MO����	���(h�;�U��ͧ[�v-N��-7T��ʋ���c�(���
�)m��꤉�O�j?��"��tد���Og<�� ��=�qc��"Sl�inN�m���%o�B,�G���*�_l¶����c'���������1_�F�~�O�0��c�|����_ӫ%E���ݠ��%NZ�����2B�y��Lا�I��������el�^�ʖǇLO%�'��w���ND5��8��V��fvjE�
2�+]QeQ�E����$�Ҝ.�I�(�i�BX]e�9Hǥ���m�<��>.��Eψ8��Aղ�B���l3{Q���Fi�h��Ty
�Q�6���C/.�<�D�F���>������H�w�Ӏ(��/k���-sEI}�`�v�����FH��b*�r��R��ZƐ g��k�=Ǘ�]�U�8e�D$-'��/))�����K���j�n�<�	���Eث-��?BA��Z.�c"t%ݞ��/
s��Xļެ�qY��'s1��3����*%����P�7���x��C?��=�r�}�H{�-y:��su�y�	�,���*���'�&��w���V�IT�P��G����t��Ƭ�+*�3�D��c5�]W����:�3�`ա�rz�NB~խ��j�h_tؙE\;�q��B�ax4�WZ�BTI�o�F��-����2iYNd��8��nN	�]����*d;������8ifM�?�|28f����#<�mՋ�ƺ<��j����扒��Y-�?��5Hw/��y~Jm	1�!Ϧ���I�`�-�Y������{i�����gl���i=h�z#e�a�EF�`�#���z���������s<9WT����e�X��<�3D�<U;}1�[��H|�@:J��>z��x�$�1�5���ħ6{g>�
���5��Ո���H�u,�(�B����LH�!tՔG8L�����IF�&�$vm=[���Ÿ#	�#"f^�f��_�G�mh߽�h��G%�����{�2C'��X�0��I�x3�� �R�m�n9�����'��D<*��Z���=#t����g�2�����x�1����`��7�E:�8�#Ţ�H��Ռ5�y	�K��1�~Υ�d�Y7��D�5SS5�L�3��Өq�̊͟��'^-������ﮃ�,�2�J^��AO�f�����É�2�)�_��X�Mr+�����s(t���j�n�<!Y\f;L�cDd�zt&�@A�]��Fp�8ʹv���K�����TٌPA3siS��i�{8��vzK� w�s��Ӭ%ɳd��5��	�~ҠL�Ǆ������dNkb�u-)9�t�'����(.�f`�?b��b��N�'��'<�P�X�m�wĚդ�	�wx�Dz��J��q�w t��$aS��K��s��0�U'�e�����[X{*q��:���� �����ͅ�������tq�c�E�"��F�U8N�P�D�]����c$����i[�:g�c4̅��f��u�CX�T6R�')�{Gf��)[���Ck�	������[��!����?fi�#x��S�7���Xy]U%�sl~jǍ��� E2�k��p\>o®3�5�y�1\5r0on<f��If��0���G|��Cy�I؊a"�dR���z�r/��;]�\���#�;wePY�o_�N���+��#;�.���\R��E.����l�H{.�t]N=Dq�S� ����Ť�賶�������)_m2�zP��J0�j��9;�F�anL.��63��L� �t�~Y��(���Dϴ��d�4�=+��ֱX�B&ڶ��;��m����YrZ�n�+{.6��7yDC�ط�9��&����G�l��)��Y���=���%k&�Y�=B�jcq�t�����=,#�Q��O�����CZjw4f��2��/?̼��CK�(�f��A��!�	Va��ߠ�S�^
T`�e~}�L�
��$���vKa�Fr�>�\�-��,�%�F���eOK��M�2T9����?i����S�B T����6�����֫���<t6��e)���o��_�1���i�#ѣ�T��GZ��7V��{s��(t�E��y�����g��ff�2.2eEo�sH��z6�$B��=m�������W�$�OJ�_q�O�}Tu9��*�n����W�z{���'[,F�8{^�4'�?�u.",�#ć?2s���Pj��A������ˀ�`����sḕ|�}h�(,��'��r`_%|�:k?k��s�����g�+D�p�c�.+3{��͢yV��=dvo~��\5!8����,�	���3w'�~��8g)FZ)�4G��q����^j������d�Y��rt	��@&�4�U��G����vM�Z�D����*��f�7�X�xy�)��㗴�I3��^2�k�p�G�<��7ɿA�l����$I�|�������ҩh9"�9)+k��s_��]�?i9?��Dl�9��dd�&6�%���t����8�9��C=W]��/��!q��3�Y����wb&�GkJ�n���u��UH��%j`���RQk�NNI�ʚ̫�v�:��@a�Ɓ�hǎ��Т���%�rc�� S��^��ISK�R��9�$+��$NT�Jlb6�����ν�Ċk�E�c՜\W�}GH�}���>z��6��pTBV�b�띡W�;�]�Ӳ�q���D��b�)jR v>M�D�o��]�Ը-�Wr��8�h��]gfQ��WmDZ7*Ja@3�D�e���C1X��Nk���K����{p�x!>:��x���v�tܒ n�r�j�~9���f)�c��ظ(Q���Ҭ}8��N�?�.�<�$��QɈ`�QgU�.[�LTv3ѷ��i��"- �E���J��VѮ�;���-�԰��ڟD ��Z�Idœ��@%c(��F�l����2�w\o�S ׾�Z}s%
_;c�]yQ�E:fH�B!Y���IR4�_]�Y5:}Ikb��G��To�Ohs���#݈��՝CX�E�^ B�]Y�!�.�.����u�T��	�a_��R��#+���ρ'��.:��s�!*��y��}/���W���s`�������������X}���y�M�7	�X�pA`�y9�pA�#þ��j���hQ�ց��v�N�c9,����=��zEY��g�b��[k!������9V��37�k���' J)��<��T�kd���i"�����4��G$T��w��x�c{�S��3�iE��:��:��]�#�嚗ڄT݊"Zm��A�u��
�qx�A�Q�۪�}�������1�-ŷ	�WmU��Ca� hIX��zį:��\�&uљ�"{`�^�O�;��� 5������˰��LT~F�R�aj��ɢ��r�\��TPT��Yd� _~-��w���b����V�yt<�`�Te����\��7ל??%�H$@޻L���*6i��_Fq'�}f���GN���ۛ�1|ף.a�ˀ��=�����'C�b�����2���NG���)�d���>�T�J/2�'����#�D��qBQm��37KHy,t5.���c���x�z_k�JVs�����Â��Eln�JHm�B���>+������ww�D�E�(�hSA���_��r0��	Y�P"�<a��dC���lQ������TYzf��쑊~%��ڨ��3��J�3E0i�@	[�ov}�}7P��	����d�=�=T�H�Rǵk_��BΊ�����>h�*E����p�od�B�l^��\f���K�E��)�;}P�����T�ܷ<�Lt�X���}�'��p�Z����(�Ώ-���/��8�ǎH���ĲƁ��E=�xյ?�Oi��0D\�����ho�4�a�_�@�j}�R�7�j���3I:[czY�m/Xz�9,T69�+��L.�p�`&��r㣑6�(-�ȒE����{��� $�1�A�s�)��T��2��(����
�I��M�Yq#����N��B�,�2w�!�Q��0��/���C� �{��;������K�P��j�����-�~��X�n"����f��G4u��ɿ"x'�.cmǤ�*�0�p��7l�_P���µ���|�v^�D��Fd��O�E�6�@0b;�<��:��vO_� �QՖ�O�U�)�����\�	��/��<��C�]�쇼����k���NZ�&�j��r���{��8贁 "v��D@3�	�_�AnζPw�����Z{g|y�"l��y�*����f�SL�H�B�lu�}�uZ�7W�Z�E֔pWM´��×����:��W������)qr7�����Y�=�er�ӄ[ʈv}�E��|)aJrE�������2�w[3?�� m�<��t�� )@+��V��L46�*����y8C��5o=5o/j��Ak�Z�c�!g��F0�����>�����h�7��=.�"%��3=h[X[4
 �����	*�����ӛq� ~�wC_���"�W�� 
���7�����Lcw�4�BR���8��}u����+ذ�i��`�Z��A�̪�����$����ڠ1�6�"k�Df��Q����iS�O�
}sW�<L`�}Ky�o�>׌�: f�]GC;~�L�v@U��S%aK�Di]PG7�M*�j_x_׮-n�w��Ƕ����aR�rAƘ|�����@E5�r��kA�|�<���M��� <骇�i��qJ�V��]�>S��|`�����}(z*׭��]�4Ӧ�UU�[ے �H�Sq��b̩#L��,��,I�)�x��c=
k�1�	3�IjM�n�s-�"�u�o�}���
���y�cu�+�/?�
�I���5���<�%Z�R.��@�8qd���x/1�mTKN��"���oU���Wa�d�H�?�\�b��ϣ��
۷�:M�XU�a�\ ٿnCU��G�A�X-�J�X����I��3����:����h�����`��oR���T��Xq�Ȧ�ԬD����RD 9vO!VHE��i-�e�x�J�^v��"�����H�����۰��������d��X��D�o�^�6���=Ҍ���������5�4}G���P�q!�
���xcJmo�V�h �k_d��s�XK�4�Yz���p�cy���iv�J �S �-":�,Dc��IG�RV���K7^I��1��v��V˗�����s���	W<�����(A�1
H��]	b^����~q��s�l�/N�?cx3�e���SQ
\�c�o�K~1gB/P�"���%������~}	=+�B��g:�e��ٸEF�1 F��9e1E�C�템X���鹔�_p�5�O�M��}�-�?jǥ��?�@���2�2͌�j��-���<�H,���Kg�LZ�9���G����q^.,�� �[zU���l���R��B�ٳ�R\���מHg��Nq/���Ұ�a��v<ޢԪiT� �R�W ��8 z%5=�:��Ɖ�|������~��6�c�����d>pʆ��8F�viEA��Jo��o�c�6A�p
��Sch䙩:�U�ଫ�!`�xK`�O���c�h�LS{��N��v1��mֵ��=R8.R����qiaJ%m���P�*�I�8�Cs˃��M{}� �B�\�a1��3ޙ���{�G][���G��w:�T�S����Li]��%��~
��7`��(�J���ǆ�����!<%;քy+9Ҝ0�*��� ��>�FȌ.80��2��N��J�?���X�`E8��A�1�5�N�LGI|&�@���2 .�ʠP�o�A�F���[<�%���0�<�_�,]�xP�(�[���3s��$�Q�L� XFz��"�!ʞ�������=\<9���zٳ"6	�Z�INQ�~��}���y@�:�f:�}���[˥"e4�\��ѹ؉�S���k�0}��qW4*�n3��M���g���BF��� ���#���=�4��	\�F�<�`-����{�P��D�w���^1GV�����Qf�F�����o=�����ɳ	@�X(�[��-�@OX�c�6��h�P�4�������g�t6J�"	\�Q�e���j���ȶ�5����}@�sI*��d3���C�g���tYbFNn8")�&H��s�\/��7��3���x�kx̚ϩ��c�N�~�V���R�~-[��VKٱ|�j�ilJ�ggǗ�gB�U�>�G��}c�'���r\��n���1ܳ�Y�?ꉺ����y{���{����_��nH�#nV�v�
Qb�Ah*�r�'�d��̰��n��[����3�0�k��a+�`�7q�y�JJ/Ko���Rr���E�KҸ$\B���#�i�KY���Ds�Eb�,�)mJ���T�1,I����+� ��A�{~�� ߍ\������B���q�j��s��c�۶���z,c�[����=�"m~��Me(�c��M���J21�Ξ�u�|��,��|M�b/�Z������*��]8��M��"�E�t�\?��F�`ծ�姃t��L�^�O���Ƥ���Y�r��^�7ȟf3��Ĉ�}�|�=�v�k�;�4��
��������,.D����@��C���h�ߢY�8:L������B�{
)�4�#��`��|�G'�	�	0��@�zׁ�.nP���Yƙ�i�׳���p|v.@�X�J�;�	�[���&�ߋ�v��GQ_�{VS��;�
p3AiS|�.��*�-��Y�0+�?��ڬ�$^���>���ސ ��ܠ��H=�#��싫\u�8ߤ �c�4��ͳ�e�~�[�t��J<�Ö[��`vu5���/ �\zr��7"�R߉{��j�Y�~�}Y��¨�kakcR�h��F��P��h`�{���WT;�ٸ&_�:��� p��X�!m���Vf�B|�N��}�?җIx��sL8W�Z�Ƒ� θ�z�Ʀ�̀�����Khr!�{���ZYiH��(�G�T�@�#���"�x`72<%��P�<c��[{�I���w�l<c�����K�.�#2�27#���Ǳ�wH��'kf��A\�3`����G�m��A�@gn�)�E�\-n�xo�:�@b/,����2�8��8����g�<���:L�+�Q�U�]�"h����R�R���l9��_���6rp^��v�L`Ml[�
�s���3��ps�~��1��0�[ivU�O�+�7���KUO"�s�\l��L9w͝ޙ�� �LV���v���ܜ��!-�����R�K�Ef7v_q�4�� 2�Zp�?�xr�'^�w�(Ň"R(���@�5�"��[��<n������Mp��}����Ώm���q1uS�ût��	����: ?��'Q�dՂidH�>�pN��0EM���rC5��,�"�M�n�ݾD�eQ�G��[�ݑ����L�;���͜�Xb�&#���o���GK)��p�<�5|�<pƑ �����ː2~�A�ݍ6�[�].)HS�W��x�ܒ��~&q�[yO_�����W�[������+B����@�8<"�@�f�����I@�V��)���G�tUuL���2�?J�a�
G�9�&N7��KGA���ΐv���BFv�'�������nMMQ������Y�-u�V�#>i!lUO�<��c�wi�P/�r5�����~V��9�xv.��B��>�F'�{{׵7f"XwM-�����f4.�[��tkt��7 ��J5�@-A�a�K�.�SA}���]v�{�R;����b$o�M�z���-���сv��{
�dr�S�C;*~�Z�h�_��ҁ=ՋB�R@�=�"��N����;�sv�UT��u�����oipI���a��,u�`� ���V�_��TM(J�I�@N�:�I\�X�
_�\`�у��� .���LJ�H��q�Iq�?�Bblg�/����^�VDb"��_"����V0�|�R	z��KQq������3 �Cb2�Y�ck��Ԑ��<-U�j�Ns�q�z��rMM4������������А�ƛbR?O�<�L���S-�~��.ʨ}�8��:��}�q�G������At��Y�<�3�W���w4��	�NM��#��� $ktt��h �%��\8��"T��1y|��Av�
;և�U��K�ƚv`z㍘��q�v���Jo0 a;��zW��>��vu��
�x��ˁ��WuI��h��A;������$�ҢA�FyPSS��(OX�n"����QSɔ9 n���~���l��$�3��M���h�L"���=�I�ȱ��uGd�ĚK����r�4W]tg��"�F]��z�[����������v����.�����g����ll�{Zx��\]����4#�n�Y���XP�v��6>#ɗR�c�O���k�Y��a��ͬ��W&��I�f^�4����o���Q[d�2	��䨳-`PV�P��B�5_ȩ���O��7����rj�AϚ��'�� Q��%9/�r�2	~���W����o6���v�䠍��x]&�R�_bLZN��%I�q�;��id/����t�g���΢:Z����wg9^*�|M��z�g�Q�i�\�e�d�C���}t�9��L�D�73q��g��J��x؜YQ�p�B�3�q�N1�0h�
֊/�w���zh�v�I����l�<M��dUc<�88��/�W��(Ly�=�Ʃ>�:���HQ