��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x������jTe�)�D�b���A����1v16�|,J6l��)~�S� �B�`q���(]�s�ˠ%��L@��z^ߴ�E����\>lt܀��|��>Y-��=��v�r@@����Q��2��^ԭ>=h��^$��f]vY� $za��"O� X��R��ȿ�u��v��\@��
��^(9������U�M4�~�&om^���O�|�;��9J0����E�{pY��W��AHgI��o(�s�����SL<�9K�	���-R��_�l�gI��9M>�5��׎m�C����E��V�e�C�FU���n%{��
]�^
;{*�>Ԣ.Q����ǿ��z 0�/��	c�� �(Τ*�?.Sڦ${#f	&��I9�z�u�4[cݻ��l'�W�0,�8#{? ���!6�������B�>%cY6&�o�>��E�aW6�t'b%��>ä.�?�f�p6k)S�\�A����.�ܔ�&�]���N��Mr�*��?�fs�ϫ5���s
�23�#�HW� �F�l�����[���h��u�ӹw�A��}˭ �J\�Ze�2�/$�(̠�tj꓃�fOD�_��)��J��+��MY�aN��Dq?^�u������,X�ěi����6��r�Q�-մx�C�T ��g��-"�{;���+`Y�i$G��t���,}�D���F�B��.wz�!��v\�gn}>�uK�A����}V~���&�;�����K3��9[[�e�e�$\<#t+��~_}�]s���@�EQ��i�R�Iy�:�t��Y�;ͣs1wl�	�l�1}�+�����#?�@Wu����U�	nVչ�����Am�%�����c�E�5��m��Ј�5�֩"xѾ�֣�#�e=�oN��V�"3�`�k���>#H�K|ܠ�]��q�0wq��a�	�q>x��H�e�F��s�**~_w7?���K��*��V2�Cgv����o���7=:������ם�Hȳ��$�i�8�e&��%�=.�ۙ-52�#��ɴ�zE�o��Q�b:]ao"�"g�3�Ac��&�6�+�EC7Ր�C~ml����˙�u�«Ho�I�e����vQ:���c��3ߜw�Hy��$�B�`�WHw��9L�酘�6kn+21�|�50s�^��To��H��t��&�B�J�༴�u�����<�R&X�k��n��J�������G&����/x-��g�q��%���F�zTz��´�0�8Pq!��V�Q�a��p���dşő*�U.��S���%��f\6��;�EA5�r�n.�E�@BZI�
W��0����}!%����`���GkX�������U��'�S��)Ep��-g.��v\!"���k��9�H����e���F�,�I��ׯ|�䪗��EkaM`'R9�7�Q�e������_Z1����өKs�[�e�h���]L����`(x"����	�.{�k�zQ�����]��F]RZ9~�%�IrDo���mP�N�]�ol�'"A����j���A��e��ҁ�А�T��i4i�9���	hL���ţ���g����U\����o���n.��~J<��c���E
DW��.��[�0�����(��.�)��>��5����~�[O�1"�Pw$���欄&��F�DQ?̛�i1{�i�dy����F-IQ-j�.`���	�Ϛ�p.��)�d���<��P_�����.���ߒ�I�~��4.��(9,�v�D�_G��>>��}ͽ2#zhC�܃����R{�|2U�n����˿�uQ�����4l�ӑ�����eZG�仁��}R�HM�l���d�y\�>�@�ܢ�,ڐE��h�ɧ1��?|�<R?r�f胍�!aO�\��S�E��ZeDTU�֩Ptۭ��NIox�-���Ǡ�N�Hd��ꩺ0�v4$Xv��Bp$6�=CX��	+�b3���/�j���g^jv%�I#OS�M��������t.@_La����Ε{>�r�&�$�i�.vYVq���;������a��юe��Z�S�@a!2��n|n;�O/��<��Tp�l^,��e�}��b��}Ia�Ak�Y��@��w-q2��^�E�	�W���MT��%l1+C���>q�u[�<_WqtZ�ǐ9��'���l|㢸Ѥ��㰄Z��bD:f?<��}A������B�ҫ¬�'�����-�Y�|Q�pZ�ŷ�_HỨ��@��=��-�x��tW둝���?����!{}�����cy:���n�(J����X���)�AB.N�Fq��/�sW�^Z��x�A[�����s-�{ԩޔ�҆	������g�
}�"���-����{`&cǖ鹔�=Z~�sn�˵!��p����3�7��7�C%��q�*��A=IȾ6z��!._Ѱ�8�`�N(�뒤�+!�t�iu��.g��>�Z���s���a(	�EO�D>6��͖��΅lP����{�&��aDZ���G�(�Gy���<} >�5���h�"�ӥe�Z�U�N��ͧ˰����3 w�P_�\��+�c"B��=���Ən6m�S�Ղ]=�f�co�%�#W��|�ד�,hD�*jQ���L���G��z��9��Mu"٩�Q�i�XE)V�>N'1�=�V�D^��KP��;�ռ-o��c�Ș�%r=\ۊqE���;���fp�����z��<�eZ�����EM,A/����A%��׃���M�T�?����j/�ӗ���ы�	+l�x]O�@gQcB�a�ğ�@|�����'���ea�o�I�r�Մ��?�r�?ۍ
/�2��(8�fia�r=�Su���*��\;�Ͷ�C&�w"�Vd�6����Y��Dq(�*t��r�-����$�u*��D��\���� �Jj��1�����<�QX ��?�}�MZB��{�u�YX�pM�;!x(�myi�t�3��u���;g7���j�~�1��m��uC_"��_��o�I�\w�T��?���<M��Ϩr�ISe���F�ŝ�l�yCv�7]������)0_���$�[[0�
v06=v���9S5�gԉ��7��q��^�ܢ�]n��u�G�1� �!L��h^)�<Pd����c*2>Ga���(�	�#]s��td�����N�T����K��u����|H��N�?�7:�ɫ�s+����d�������r�It^%.����5���ƍt�W�x�&�-�|�_�`)��8˞NȨT~�6 ���O�{�G��eo�VK����Ӆ�&^t��A�σ�gPhG���v����������6�&޹�J�a]"Mt+���m��LZ7��jgݗ����ѨP�k,�7��L�Z52� f��nW��o~ӥ	8�?K]7?�8�Ґ	:~�<P�,R3����U��#�٘�j/�Sg�b�p�3�M�ݍ�Pi�,�0����Aέ�a1_&$D�lr���R=����ܻ�W��
f;.���U�=='�.���:���<Cö�J�V`�[�ȩ�%��(�9�@��Z!��U1N4FѬ� ���
F��kW���xQv��C���Y�s+��I"�=(�x�'n)�Z��O	�U�f�m��I�Q�AQ�;_֙���At-�z���$Ð{��� z{l�Q�԰h�3�s+�zﳁ��m�f�W>�t�?�my�b��o��"��]��`���`�+PM@;Jdy���;�6�Yf���z��X4#��j��5I�h�Ԣ�p"�6z�)yEݣ���]m��T�H�R�3d�]��x/��9�oXR�Ñ~�u(�r�"�t���:�'ҏ�����K��z���gJ�sytO�zGݝ_�׼{?n[Y����=>=��j�[��Q!7J�!�� Re���`�d�a���$�K}�B0��u�yĖ9��P��#2�ۈb��i����ښ2�w�[$��`�Y+n��>Fڏޞ˦Y~�����Ua�b<���5Wf����A�J�fz��q�����&;>#�1��}��n@�meL�0~6,ma��E!�}�����N�c��_uQ>׀��P����
,oxk��z'}_M���.�j�&��>1S���z�Z�>ɺK��A�-m#���"V�	����.�#?��
u�u"�HH
B��2ԟfc����g���Ƹa=����#����������uA�D� @�3=�4�Aǆ�%?hfC{�Lj���������i���G�Ip�= Kd�1����ϰ��`Dm��`���]�����Ni` {6�V7W��sxo�n#�m�)'�����e�Z��d�L�����#H�k��<����I4���:���5�2����b� |�X�+�� $n�M$v��
��hn B^F��̊�K���<˟�+)7������~F�
�~�~��]O���xպZ�v1�y��é8��Э�`���K�l��*Hz�h6�)#4��DR(��+�����-�w.����eW1_���{P:C`��Dq�t7>��^����}hf?�=��m���꾌x�|�
�@f�q4�ѫQG���3��*q�-dq�㢳.,�ґ�=����ܮ�T�d�;H���|H���=G�����I�&P�QU���2��5&թ�p�y'|���%�aۄ����{��`��ZM�򢾤ۆ�LŢB�"I�NP�r�v9T�5.��2��A[��]�:F|��d𽣻��xd��cQ]�܅�2���B)���Α����ҵ�]�}1��ni��%�D���އ܉����D��:���	�^ބ��Ee\�^ԇ3�S�x�و��U����}�k����\p(|���4��.����/q�9g'�S�4L�6Fl�S6>�����˙�M�@x�h,��'@�?�Eg���)̆%�BPA�ḕ8	�ᾒYQ���#ۓ7�Xp�1��̈́��G���8!'����]�n+�`���$��P�e���"��)�&��.�^0�e��1�C5�|k�N6k���[��������C�ų�zX!@�`���|>냐��qع��W�a�����5��q3�Ӥ�I"�w�\Wm�����1���ŗ�nQ�f��.Mhцe��0N>V+t0�+~R@� �L}�0"��t!Gc�=�����T��`kˈ���!�X`
9���D�Ip��x'҃J���ٟ�!`'�����Z�NQ;n߲䓌=��4O6�&��$�
�澭�r��Blwyp���Ҳ%����]�n��&��q�S��0݆I1Dx���g�s*���C�1l���%Yl������T�a�"�^��Jq	�+����\�L�u�ѣ|�ǉ?E���<oL��(=Y����~&����A����b�b�=:��+���į��
����ڊn>Vw5-����ά�w�E��ގQ|��3���F�N��h�����=74"I9�X?��3������nT��ZJ����NLVD�<I�z���#(�r<o+�4�b�4�?�}��#=��Q�6i5ȸ��A�o��qڣ���� G�兵?>r��2zC�\xלn�O�����8�a=�����輇e����+�.!�#���c"ƴStL�pl����y�U�����/El��f�'pj�&��ϗ��Ⰹ�͸;_�����ǕkD��K��hc�1r���a����������ţc��"M��;!���x�;������L��P !=d�!�b��V����7�KQP�ބE��i/�8�r�8�U����_�Z$�Ey�yYR�p��3H[*�r���70g��om�� <��b<+��1Lg��l�w�³���.��C��a|n���o��Ks�sĥZ[�S*�d,�ď�^n�H;��l9�%��U"^|�s�	�3F�GN%�:⚣ɟ=,�Tm����3\�.�c|��>_.�7��gȆ����!�?��"��0�Vp����(X�V;p��b�R���"rc!о/��'|�}�y��E2�g_Ӆ��4g�e���0���u��wCSy��R��(�g*� ��J���6����y�&L���p
m#�m��P��fm@l�Y�n���^ľf�b���d�g(W˄�i���{#���O.�b�6;��A��B��"�m |��_s������b�$؄�r����G��fܯ뻋A���ëN��c	�)��u�I�s��}W��Ç������F�%c�#7u��K4��y���0�i�a�-��pzs��s��6�=u#�B�ur���r�
�l XH�&}Kj��}��>��!K�4�SK�@һ�z' %�WǪ�nl@vwj��nj�*�0���4�Gp�����G�c����"r�ޠog��@������O��'��`���w����|\av�j�([f[QW��"~ѓ;�}���0�*�n��=���e�Aa�X�==Lzd��9e��3W#�dlQJt�ؼ��O�k~�8X�[��p��"�
M����C�&���.�\~ŭ������藵c;(�;�<���Hjx�H`�ؓ��X���]��O����(���I�	����?�P[ئ�$B7��H�t�v�'|�>��(Agh4ŵ�_�QW�T�ΒrXO��QLﬓ������$)~A_���"Rgh9�x+C��s��:"x'�����y&����Q\:t��<�f������藾�o����C;��N�q���0+n�S���n��Ƭ��&$Hl����*��3ϥ�ģ�D�6�=fH��R��8#����8Oar�7���lj�� �>���w��ONӄ��� �(Hc�J�|���1Y�H��}��6��'�/�j���l���*c�;�����Y&
��_Za^�#�+��ͮSБh��eK��gKWA�&v7ؗ��7d����o0��MT��ʒA�C�7�}p�`�N��r�Rb�z�+#
���A�a�})��2M1[�%����rQ�`X"��#�F�3���Ǳ� �*-�Q��+�)�E��WS<���r������+�l�ُ8��"�~}�]]����@�C�"f��ȫʎW������2����r���[u�5$�]`����0q��e�"� � AJw{�@�b�5xa���n������tϾi�v���Xi�vE*�J>Z�L�4VZeE�`��g�-,�4�i`������X�i��Q�$ǵ��ڂ�_xXQtfLF�ܔ�6r����4"kG��9�;�A�~�ȳ�a֌�kT�/5&�w$|�6�)��+�;��[�l�%{�>P�?��]�����ہ��ӯָ��c�j��r@�ڐ�/֓�}����ؑ��2�p����z�1���o�0_s�d�\�%�n�\RDc���aC��Ό��I�>��庻z�)�9B
�u�P�:�5��J�/ 4X����R��2�D�)�����@��ZhO��c�>1c�9�Z�d���zZ��=e���U:Jb%2������+�b�V��N'�9�!������Ѕ�\!<!�9e��WX�($C��bWpqӞ�9�|[Dx_�Y�����(ۣY�=�Fj�N��:R��D�N��'|��aMI*'V��sD���n����U���\���J=L �<�h��%�gO���Vщ�V�����E�z�s�G`���3d^�x;?Jl��y�*'i��%�D+d$�F�hF,M,��>>��;rk��\���
Қӕ?��Jӂ[�ex/�7-���Us��-�:K1&O&�T9K"�"l{����u��>��VR,ʈ��W��V���7"�O���q�&����^�͎��Dڲlw�6<���I��)�\"C廻�����?N���TY6ٍ�P�>?5p����߻�=u��\�u�q�[�T�|
���7��d�K�9���L���(�kϫP�`d�A�x?��+��AiMFN]�m4�p���p�y��i�L;��\�r9~>H�
���y������O�K�g;,'��6�fqRs�8�hh����e8}3�5.\�[��A�������ig�ZTKm?@'f�������`>�7;R_�8^�o��݋Z\ƾ���/Y]��?���fR�3�:� '���D#I��sO�T���U�����[Uj�|w,D�Q�Q�3��݇�p��*������s��[�v�]�.L�ϸXB�;�j���m���,ww��?�&`�����ǭ��t];��c�)�1P)j)�QY��O���(�?G~�*��-tt�0C�smuPY��w��0'���|$�xo@�M���?�Z���]m��o��<j��*i�Q������m)�XtKrQ�pj/в]
>�8�֜� L�o�Q���5/�ѐT<��42�F�'(E T�r��9�O�0�z@pV-�c��B��/��x�U�tQS��κ��}
oo�2ҔJ�QL6�8̎�!*I��~�r��Q���33�C���?��J�5�w:D�`�f�,��Lϸ푶9�|��!nR^��3/��j�Nls�3m5Rk��Pq�r���LW�HW�g��Y>����¡"�F'nS�2+�h��l������L`��)9?����T0������!�+��e�6 ��$sQoRH)������퇢Y�~��`���<���N�o�'7����*�B��G�I1̪"�