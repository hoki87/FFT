��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ���������dI `!��d���|��Qs��+��~�ڴj�/8�ꉔ/�pb�j&ǃ��^;�iÞA��kh�(��q�cD���[L��n��!�(�����w~?�<�j��-�x�s[՝�X�_��gZ�
6�����ɻ%�V���Km˸f(3岻J`5a2Țp�(ʣ�VI�)�kQ���]�!Y<�@�7�U���iۀԩ\_^��,�s=�L��B�~���Y>�g�甆e�� �T� �]>N䌎��x�KZ��)���Y��;9�����M$�N�N램s������%�����싰w��.�`���jG+��rդ-	���"e�S��;�����⼥|9�Q�?�)��3oO�OgXF5O�*סs�at��e���F��@�|-��Go��MP��YaJ��U��Xl��y�"rE�-FF�W�gf��]�t����k��Ц��QW��-Y���z�|B����pJ�7y>��'*���5�4� k6��=i8^s�C|�Yf.��1<y%ſu8fmQBG���[����������<�E;ӽ\txJ�,�X�o�+�F^� �ӝ��D��%_�X�4D}�kBF��J�Ͻf&IMɤ(t5�w?���;�U��l�e/�X��<�3��/���ip�Ii����l���_)M�P��v*P}�a,yeh��1�dA�a4��$bv�?0�H�@ԡ	T�:Q����;��Σ���)�Ƣ�k��t��kd���vl�x��k�6E�*y|I=�4���԰v��Ji���
b�*T"�H�+��W�/�+�K�^ZH�y����x����n0�Ai
��{�7�-ɮ|�3H_�	gɱˀ��D	|���c�NK�|�����]�����	��{�Ĳ �BhȢ��9�N���>k�p�J�������x��9?v9N��F��F�+͔G���Y����Q:�w�{?Q`���RM�����I�Y�jϒ^��]�B������ɖY���.A�	fp_عb���'��������y0�SA��Uʔ g�ޮ�O>y���q֊R����@oB`��.��h1���^�V��=!ݷ�z~A5��p,��1s�;"y��#�����P �D�/�"�]����"�Q���lf��F;�����E.�d��7�B���$�+d[Ĵ��!]^j�!�?'$L������g����G?������0�s�1T�P��n�:��_��T��Xt�$�B����[{�!'�ð�P�w3tY&�Fi�f�{�0��9��mYxw;.lX7��U
�ѫ��.�U9q�^Օ'0����� ��#S�j:S�Ku��)�ɹ6�S�~or:�L����'�{ȅ��y�L0����?}X�����D�t�]b��`�X�e?�B�2�{�W���/>f-�i�t�K��(�Fߛ��tnf��w?y�����/�UĲR������7nr�*D�r7�mL?�ؤ�<�	���u^�����׾��kj#ǭ����#�#����ܔL�A��v2�`#��a��������>�	�������=i�(�T�#�&��(f=l"�Ζ���J�	g�8�fZ��;W���u�hw�p#�0��������!m�:쮺�iB��djmX��J������cxWQ`8��J��]����sm�w5�U��\���$��*����mQ&.������A�jۂw�G�'�K��`+�H���n��a� ���;�#$���2	>"���' dq��WnK8L�G>�6��;y#2$f7�o�
X��˷�/��N�T[���·��]$`B^fŵXI�*�E�tZ�nWK�^d�g�h�&Py���H^�@a�����f�hK�4Bxh�X�8B�#��ĈYo��0Ti��9�z���<vZ&�8������$��F4|�T�y2f��}�P`�+��Mҭ�r�Z�%CZp!Q�j�H6��u�!e�)�غ<��]������9��c
�y������7��g�?5�`�r�E�m_Z�K��}"yD� K��8zxVc��K��?�w���<�]`.�u_��o`�^�;+��o�V�w|c�,[�s^�Vn���9�ǝư���B������K�=y^7�Y��ȼ�F'�ml�U��]���﬐�h�����	�0�&�eF��%a'����4���!�w�-�c�:�R�W�h�	K�[L �p�-B��Ĥ���O��_󃉬%j�^ѢH/4~"ȏF�Pq�X�|�S�7���6��ẹ�������H�R����ƜC�� %��cB��Ӈ`z��U>��F�cD�f{t z�J�Ukn�m�3�(�R0/9n;"f����XD;��{Ź�b��	V9-�jR��߿��ݨяl�S��5��c#�V�<��^�H}!==��\�g'PR���H�:��9�Ā���i�N�����g71HTl��tA�Z&��I%�(:V��˂���qÄ\[/"D�6��L݀���Z���Bi_l��_�v���,�����ʦ�d�a<�b���[I��+㜱���A�9�S� ��`,��7K'��0c6�"k�W2r�7x-4,��B9VPr3����*�)k-2�Q��)|��Z�Y�8��gyH��q&���)�E����=��.r���9�kq�/h9Ba<���FY��N��c��OFګ_#�$UG�*`5]�x<��+� |�oq�r^}C@����7֑:v�{�U��Bj��XQԑ�(i��\��7�j�-��+)�s���!Q�k?7a�	(��x���#����^7���?]��O��M�B�>��u �R�렍�>Zxx�����o	3� ��]��2P]4%	UI�:*G��f�Ϗ�~��%�%��?�F���`����_)�b�pԢ�s8�e���N=����1|o�q���/���&V�q��z���b����K�[���������9�0V4#�{rל4;��7��}�%�y1��nWW�\#���&�b�����[q*|6��3�z��L��G۔������A	h2��|_����C}�H62�ɎǛ~����_k˃�|���iA.�K�T0�/T��n)���2�ƕ���]��HMtTVG��d�i��p�UF��'bOtN�ef`E�15"�!��p����� �d�|���3f,�( _j^��|� KѪ�aJ��X��c�L�=��#D��s��`S]��Y+.r�G�'HvO�Z���O<U5j�FLa
L�.��ى܇M�_>�*���D-�!Y����t��~�\˟D�u(㮒4�z#���:�ҏ��m��M4��*�4	���_�E��
�L�߁�"6?�&���G��pͽc�K�(�q�H �Ƿ���|n���b�.1h�;	�?�������_�ӡ���7�v���r��Q�B�74�q���(��5�˃�b�`Ƥ]����ʺ4�JM}}�=���K��9%=>���S��T���ͭsz�'-����F���Z �Kx8��|HJc3�����N�@��i\|�[�%9�Ū�^��77Z���� �3�U��nI�JS㲹�|�U��-���uϛ5�SU<�xCl�����-���3�_��C)_P�D8������,������� �n�b0W��g�w_����A ��䵉%��aH����̓z��\�����o֦9�;�Q�@�YH´%�j���R@݅`A�����i����q��]?�i�&�]@ ��5�Q8��t1����V��G#�U����D�*6���a�Ӎ>��'�<�ј*W*3�OP�̰p�Uvx�>���ٽ���2e��R��`^�[?Ӯ$�G'�C�3�ǡ�(�$q#��zۦ����y_��T+B�[�l%T���`��^����|�%"L�Y6�*�҂]�<t�m�����x���Q���C�e��&MZ�T'�f�+��=i,g�`S��k�w;�ZM��~.˄�a�̲��5n8s �K�9�0+��'8�J����O ]��u��%�/@6�dlp&I%�W�����[�gT�[��e0*~κhp����X���EM h�?�Ts0S��3�e��HG�J5�j=x�]s,�#'Y>"�(��P�c���%-�To�v{�����+d6�Ϡ|&`��[~���x�'S	�^�.ՑZ�Q��}V�[�
�x]�e��y�?�a��ѳXK��i����U��kZǼ�7�s�Ƚa��8Y��͗���?��I<������t!H�I�2CO1|,� R����D�G��T֢�j���uM�����^	�O�����y�-��ڟ
�\R~ڢb�i���+<��K�KْE�Ɵ�Z|AD'�8�h��knX��-4폤߼�&�����ǂum׆JHri�Zlmx_�����Z���K-:V���
m�D �T�oĄӱo��Rxd�\�w�Ss����ݡG1��##�0�+�u�b�7����x��������r&d�x��Y�������1Fd��W ��=���"�/r��k�tc�|�"���? a��x�S�`*}�)6c��MI��~�WCPu��׌��Rͪ ߽��߲3s�m;�Z5:$��%(�f
����-�2��64�!�!f�|���޸�p��˵ʨ����E]H�g�s]�Lf�?5.�l�U#ٙ��s���w*�N3�+�5�P�ݔ����x�*�D|h������!�7my�%�U.ح�n���b�՗�r���W�fؽ_�����.l��l�5�Ε�d7o�~����T���^��$��xMm���d���F�4�8�)���o>��� �6d�t�h�'���D���H�+�����aiu=���B�4���+=���51t'0�Q"���[��c�ո�SҺ�>��Xr�|�B����fR��S��]S��>�̉]zq��^t�q<z��v�hR���H��&ǚf����������E/��;�.�?��k5�HE�Ē3�#�|���Fx	���k�n!C���ɻ�0����rn J� ^���I�$�U��;��(_����0�@-�|d|/�,�Ԏ���äRq<;�#���B�˟��\j'����ܢ)5T����'F%$v]�
�c&�,U�,Z�� �m��l�j��F�c���LJ=G,��g8Ry�$^ْ>��
%������Ԁz��²,-��������a��ߎ�Ư�|Rlļ��p/��F���hw}��C��o_NԬ�,QvF8HC���v���g�������sgp���*�8NCI���h��)�+�wp���7w�Y7k�,]2��
3�!�݌Z�)"E��`���;v���֥���/��)m�����Om^�[D�}��g��(�%�b�QX3NY�1�ު!9�ye '����H�m�=�;�ӻeP�TXqӯA���.����s�g��L�|�&	�V��u�\B ��@�O�YU��c)�GRT�fD7�{��N'�o�R��/pT�w��:������d��a�yE@�hA#�����=B��䎺3u�� �F�2#�� ������r4aMe)cc��Sn��VI��Au0=�a��N��Ze_�<3 JI�&�Kq��^��2�Z�+�u��K%<���%�th	ˬK�q�Q|rχ֒B���Ӛo=Ea��M3��q��||\|�Fl�!�y��C<�3uO�Ho��Vc<����rk�������7�1L/<蹺N>�x�Q��S(+�ʨEI-|o Ж���/�Qڞ���U�'���q˔������:;�O߂�;Uw�b�=Ca�h�y���=�g����H@E[WJ�ٖ�,Ɉ�P8�VǠ9eZ��Μ�d?{�S��c3�pp�y���uHj@�KnЋW�ﻥ�Em4ⴱbr:�QdUZ �PiJ���iO�и�����%"��۱���d�Ai�ڇ�����J5�kX����g{dl��1bT�5���֟��5yM�sǐ0�	2���
��~h��� ~�Ua�8��긢�����9-9��[WE����Bl5��v�����j�R}���A�!���:6�d%!q\&D�:�-�~b��C�mT�l�V[0S����ڼ�Qk���5+e�B�c�vD*A��A�ۯon�͵�k�*X���Iyv(~Ҧ ��;��u��Kݣ!Q�&Nَ�ZIP�{�B6��k�=���كvE�-�Q��%q_�eh�&/1C|�w�H�Q��,��i0�x-\�2��
����ݝ����&�~hZ������H�e7�G���>[��y��
Ɠ��ͩP����8ĩ��?�D�[��V���>0:v6�
H���oĲWfcQ߭_;��h�������޼�������D�9�Z:���*!&Ao�8�p;��z�3�#q� ��f�+����ӷ�|� ���F�"x|G��E
���R��O��]x8
~����D����n�6��y<�r��XV'j\{�*TX�J9l�>Lه� Rr�'�јN�
:˱[E�Fn��|�q�:��C�Ǳ#P�����S�W`��CZx�l�B	�%�D��	3������h�u%L's(_���c$�tBZ�Ћ�<�����r(sh�(,h��m�,�* ��0'�f&��ln�e�q���������hp�*��CÓ�7V�3pG�=U���Y�+����|ªSz�ӵr���i���$�وS�FAu��ŏ#�P�ah�ug K�#��Ю�x^����ZM��F���$�����2?�"mh�B]Y;}�r�SB��E��<����[l�0��C�}�Z��r�8Ouw'nU&������'PF��� k���&T����$�-3Ǟ�2=��k?.���A��(����E�k������=i�p(i|c�� �',by�4�D��y�n�Bw�#�oߵ�v�w������)8j�{"!D�L���?�� ���ִ�Bs$����=�)�d^�Q�}-Z)[OM\�������N�׎�/QS��_�q1+1�{�wZ�X�]�-��M�M����8�]�u-�V�v�����Q%au,$�c����2�Ŝ�E�0Y��8��=��5����LE�B��R;h�M�]� �%���~�نO�r��չH�����n��'H�lPI�ޱ�����J5�x�xO@�eћ<�J�C%�p?-=�� �o������2� ?�ke�۶�<�!���Z-�c����A¯G<$ ?��#&e��_5��oE����OA�n��@�ܣ���GA��L��a�n�!Mj�wGѹ��d�N.�NS�R2,��A�-�:�Ʈ�Ӛ�����e%��Ƕ�[I��Cv���g}�D�­�kF>z��?�6c�`g����0@��w:��0�L���n�y���co�x��^�Y��1T0���BJ,#n�X���d�d�%yn���܉`��ɺ���yx(���"'�َ��ww�N��?rfPޙ�{�[��������C�E��|���)�����Y��9���O�wX�S�5l�{-�)Xh���V����_@�QD���JҹW�g8j� �-J�����c9ơ�S�L��l�����:M.(���A�c=�NKMVa�G�C�5��3�U9Q���VS�����-��2���	ޝ��� /ߒ��o��"7��vA*HFܕ(M�)�{,���dſ�u�,V�X-��|֫c�T���z�(`�Q��4�9��b��+KJg����!W��H�A]*�@�i��.�s���f��Y�T��P�e��5�^��Ů������	cGΘF��� HT��ǔ���wi�������2��!Q��ץ ���!;�^�^l���Qm�(�����e�$��;��Dk�\,�V�S�x���x����� {�t%>m�X���aeB#������u�p
:+�9L��_�P�1�N�$u�n�Ӂ�<#x4�HG�+\ ˢ��ј���_\��2QƵT-���z�x��}lM]�}����=TI	!�V���`����!"��QVऔ�-4��0�]X��'g�;��i�5La`��	�=��G�?�7y��Xu�(�StbR�8�>p�	L��3}Y=B-n��w����A��s++:ݬ�w:r�S���=uy>�ؤӊ��6�Y�D�^�0'$OО)������?@�F�Kf��=X�8���[a���S"�v�ǚq���A�R�P*�{F�ߟ졫������ƌ$5}��]F!����v>��y����c� 6/�P�U��h]�Ɲ(RZ��Fz$�
d�B{;�p�)�:���u�[�N
c��2���-Ҥq�Q�R�n�ßG�����ڿ��� _�zq��6�u�K�n7*Yכ�.�G:6�X_8�r�cxC�S�Jǵ����l�,�<ɡK�N���qm���O͠��L|p��?>E�/ٽ�򅳛E���;8ƥ ��U��AT�lt�7���:?��{�g���������	���&�i,�\�º�2�1 5�_�^`�����!>��7��R�پ�b3Cp���Q�m�#��S�G�1�b}b#�����'��H�wq���wl4@V�i���#�|O�=�I���c�+�C�heߤ\ڍ�YD�t�Y��d�ئ˪�4(�m���Y>x�s�h����Mv�:�z�o�	��M��}���/�at�����>�)��H��N��ׄ&wuÑ��:&�3�p"_C��'�/��4D��K�v|8�5B��y�ڶ���OKs��>*fG��xwE�x��b�W�U������Dz)��&�w��~��]��2�M#�"�u��8�Lq���`K- {ǣ;>zY zP���@���*��d�-�v���!�9�ʿ�ÄAKD��[�{j|��(�)�Y�[H�F?���ԍ0�����e��r��	5�ݠn�w�l\Vk��R�ńj��D?AO#* ٦�{����Q�%��ն6��-���QKU9�{:�R��"H!!�.��9��_��2[�D�ų�bwJ�C����x����� f�Q��0�hzأ�S��19`�bޓ�:�ye���I��fS�tv��d.���k���[8��U�.�ߕ_c�3��)r ^-λ#~�
_7i�_�ـ��B
�u�E�l"���#XWpb5#&�b��XvV��b���:��W(����L&�3ǝ�X����5����~�6g^�Q1���G���m��Z��XLX��� �Bl��>���m!�|؃�Z(�u�B%��a�4�����'�e�hC�z��Ai=��YE��^�>>T��^��3K6"������8J;l�q�}wB:�r�ȃ���]=\�64��R��^�k:�aM
.����k\5�u�wG1ds�W��x@�R_款݆�/�߈4Z���|�`&��i��IO���wQǤ7!��
L�!�⚍�n�.u7m\�`�)�c"c�U��:c<f�t��k8铏�b�Lcв��5�;��'�n�*����:�(�#��j6���OWpV�)�*ٹ���q!��<�Oϐlm�}hݸ�y�t5�����ŉ7w��۰Y�#(���j�S�$O��m�4�-�MiV�q	H�Wd��%Z�����[�� �%���Vx��	5x���T!���^�
�����W1�hf(6a��\��w.<@5��F<q�I����{<�iDK��)���w]�!��!)rE����Z[T��M'����M9���k��jΥl�{��G���==7T��,��m����߬��ݍ�S�q��-pU}�C}�?���럣�@��<��䅕~J�׷Z�b�Re�> K��zl_�������׵(A��!^�C�G����j�Fsf?�j;J���Vrʹ��.?5M�N��쇺pfB����Y���֢�8h���̌;|H�G#�]i/�K�Df����B��O�Ye�e5G�zFQ����Ƌ��FU�p����-d����G�
�.�^nA�Ł������o�}|7l'@!�B\��*�E�zz7�,eI���5Ø�����T1�H��3^$j�/t3N���&O�~�U�"LO@"���hLٽ�׋�F%w�TJ��S�ٽɄ~u����,����)M=���b����'	#0�IH�I?�o���ЇH>�~�����r�hy<��,>�
]�������-�|x��>�:8�w��=��.����������J��?�.Y��s^���4%�?;�o5�:�tq�s}<=	����E�n�9�f���ƾDf䑛5A�bH5&�����%ڞ�!��12�J'�����j [2��b���SG�VC=�I_ڹ�cD�:\.���D�QB�B���Y��ge\�mo�9�钰?���xW��>���j�/k+Qz���u{�Wݴ?U�;ԍI7��=Y:��OF]��g��
��e�e�P5Wt'�|�]uJ�����lt.zo�9��K ��F��������$Ѹ�Lp����_�����7�̛�{A�삻t#��ἼL\s�0k�;gԟ�z��т�L`�����x���Z�F��?�p��}4�?y,��S�0+s����,��n�o�F[n�@����D�H��������p����f@�]�u�Ƹ��2r\�p�ҋ�qZL `�����"^�v.R@`�܃�u�E= �a��%e#W@�Z����KFE �%�/���J�>ck?n0���1�E��k��
��E�=�yw�)l�O�gX�e��ś�5�	`vu���w��pg��t~*���	n�:��@`�R���I�Psڶ��<) 1�R^R��Q�V��T	�&�gȫ�N|Z�;�>��)�Ż`_��=/	��y7�A\��ۮW�9��'���ѭU<�I{�'�=[H6׏��U�C�PJ�r��hc/}��	����eN�Y�s����4�]�Xj�A��>G�|{eV���	]e�ze�Y�K�uk���0�c��Ft�����u6�M7l�sʿ�T�� ܎�r���97^�|� �=�i��s�Wԕʒ�f�sF��X�VK�ӀN.�����1"LG��X��	�+n�7@����Y�Ǉ���ה�,�R��Y�y1��\�bjm�?Gdo����rQ�dd*����uA���n�w=�aqd��#���� v�l٣;S�w���q��V�⍞��n�H���e�iJ���� ^�%5����M����^_�s(�O&p�7�}N���DX�K4�y�p��L@���T��?�͐��	6ZAr<�Ve\iI��,'�����hm�p�QG���dl���e37���b3�ep�8�L]�l�.���d��T+�#ƫ%Z%�C�N��X�23��Ũ2e�p�3Ɓ!�p��CZt��CG;���"�<�,�9���OkG�}(}k_�L���5��&�?�y^���Az~��L�W�NgJR��Itڕ@"�@X���݆�� �% K���k?��N���iW����omx]y�5���]#��}i�"���"	����~k�S��l��@k�� �Pe��%J��C���_�-RO�@%�t������U��s��"�X�UG�R1'����T|��~�����y�|�(��)G� �Z�g0A�
�vQ�H��ɴN2c�R���4�����`$�Ii7�7}�EbE���5� ���ﳎm�cF�/� Esk}X��[GSz�v��k����0��N�4]��ţ��{�p
i(��eO寘��D����P���&���v����iJxj)Ӽ�%99�9
��k�l��Md��1�>��mĴ�V[J��+�i]�c��ዝ��������c�ho�Ow�����|8��vw���D�L�=Fk�C�Y�w��-����pu[-c��nQ����C���II�<���]�*�AE�}h��HI�y�Y���mH�����S�4�&��E��w��q69���R����Ȯ�~���>%,@�Ļغ��ׁ"x�@0A���F�,�JRRzo�@nFt�e���B��z��_�¦n����{w�5Ӥ��#G��Nl�ɠS���shc#�$���������Ѫ�ʖyd,du�n.��,��	��qj��j���0�/���K�*wy	���J��R��#���p��F�ӎ�>�u��Tĥ\t�RgS��u�oq>��o��W��D�e�g�9�VT�qh�OI)aL,`�j@�)���p\���+YrP� �H���G�Nݪ��Ci�c��l�6�8G����|������΃�9���Ö�
�dQ�`�=9�ӴX�
�._�_�g	%�H"ԑ�6�0WW��v�a���֓��q9Ϫ<�Nv��|B�����~���p��{�{��
��a� �^��	�Ѱ�B�|bY��u���k5#œQ���K}�.`N������k�S�׾�����+=���:����ZNV�, �Y�k@�Z�9�a�[� �<l�9�m)q�,\@^?�OQ��4�:� l��ǁׄ�y[!:
v(�޳���F�E��}�O]0�T��y���?���#vPq����LC���B��8�~��\��\G���=�3�^�Wa�� '����1�c�P�����G�F�K��y i�߁����?��JZ�}�[9�"V�&o�"1�j�7�:� ��� {�2 �[��{X�%Ht0ıq��f˺�:y��q~�2� ����{����
ߚ@\` �4Z��XEJM��#ؖi)�M�y�,<^o;��}��X�`�^9�Q�i���҆|���=IXpS�8Trњz/PYXZMc1�����l����9�6;a�ve����ǹ�0�j`Gj�ƴ��}���I�Q4@�^��(����٪Ht� �A��j �C�n�֚r ����Q�a�Z��)�Π���N�!�qkx#��~��0KZ��>ܫ*Zp��&�VO�'�-� �"Z2x)_�,�+E8)	���>)g� �;_��w����~��G�p�7
ՠ�����D�X��$NV�z��0%�Qo�F�����׸�����N(lMjE!3��a�pݺ�e���9
x�NҚ�@����>0j�
f"ƍ�j�}�q�������'*k�i�Ч���KE>1=�`r��g�&���ܫ��H�H��0���E3�9D=�Ѿg��ǁ'�3�a��ڮ��~L���i|����p��QIT`͒��he���B�#X����]d�%yl�F`�Yf��,"=b�"�ll�Q0��G܅׶,�QN���_J*�&Yt))l����	t���F"�l�m&��Kè��&����OF\Ћ��BSL���7�	�����+�%2g�"E����M�`h=��P@`�_ə���f<.̻���c3���Kǳ��ր�O1�~"Ӎ����F��:s-*������.9ZӫN��a��k�b@:z)�� ]dv��M�}ˊ��ݭ�մ�$��A"��S�6?��e��n4�
Ƙ ���3��M{��ܨ%����q�lyK�^��<�:=xii��0��������$��Śӊ2�(*�yR��8rk*�Q�`�8��)qEFT+X����o��m�YќB@����#3;e����@��{	�����~�sc6�F<k� OP[-�Y���Z�x%mq�m�g�^�s��-&�j�O����*<7W�%3i���Xh��T'�.���-P��1�y;�Jƙq^vs���*��x;��+)ˈ8���j�#F�"א����W�e��/�:���2U6��g�v��m���f�>r�Dx}6������$�ɷn�7�m5ϩ��S��e���
�������ս0��O΀6}�E�
^#����1�K9��D�Uo$�p�qd�d�w�=�T����L�P��k�|�٥�q/#j��\�|3��c��#)�	d����?8���&����S����V|�'-k��i�J��󎠼Vׅ:bW�\��=�V�̓Zʳd�<�����.=TԨ�#rmC�%�������P�/�����{��W�o˥�w��(��'�O~d��{�-��k�g��A #��~a��]4��Ծ������$�X�̷`�wZ�e�9x��rr˔��J�r�t��b�R�S�U��<ջ>wJ��sҀ �k�=]�_�5�J�j*�����PU��4���6�k��� ���X��	�H�:��.�mb)� ���e@f�w-���b|:�	/��$O�������?�`��Z���{r�!���Do*s��!�
i!z��Ͳ���%��E��Ui�YGܓ��9�܉(w�m&����TlZί��? i|�G8�#��85��l����'���w�?Z������+24�v6�\��](,O"�I'���i��}���iBn=�0�k��ŘՄ�;�j��������S-P�4E�5h���4��T!�*lZ�,�K�^ӕ��xK���	ǻ�� �j�j�R쒛�̭�!BP
�vŞ61/	Ň�עuB�Oq@v�91{�`�T	�6�v%����;�v�0ҨU�_��~*��̻6C�6~^��I+�D_U։_dř W�|�3���Vr�`Y9b�_�[�:�,��h��B|{O�� �y�,66}ݤ��n��t~�U���B�v�L�M����#0G\�ƊG�
.��Xp�{�ˍǊ��/O0օ��7���ia���<�U+����ٙ�=�b����4���>�Ւ�UL�� �"x%��VU]�_��q�9N`��ZA�e��C�ͭP�6(�3�����V�,/�^^�Z)��p����+ ^I�bF(��/�u�̨z�#䞩�K��op����L���l�q�46��k.����Z���a�ퟩ�SI?����%��f1w�\f #)bC��6��!�!&��*�"�m��c�>i���D���M��%��������esd�x\^�t?1̨M�c��Q��w��X��%P󇦧�7bO��^DRx��o�d���j�`g�Z��蓩�n�Rf���U��$==)a�B.���V�M���	���ƹ�P�8s�B^���K�!���)C�f��h�6�� Rݻ��"���}\δD���6�2��^ A�y:-^b|?�	�b�_оs��j@���CϮx����j	�#�HGA��R�z2�O��Z�����2KAx"E^x�霈�H&���7BMrwQ�B���~�8��C��`Q� o�	�i�^�y����g��p%JwWo�v���n$�*�;�)�	�E�V�em�N̈ IZ�S�_\N j�x��E�BZ0H40���k�W�r��n���}j�ͿR����+$X���Pg�DV���1���2F����.+D���\qo�;z��!+ ��Z/��+
�I�;�%Z?�w~���v��X�G=�Qr��^�߯Y�/����O���[�������/�W��QqG3�wZ��?Y�!�2���݈��y�m��aX�A,x�M+�(�F���y��/��v����#@�p?ɱu��-g�Zؤr��=�c-�b{=�l=V��iǵ�?0�E�3����Υ6ֶv�IJ!Z�s=���Y���nHZ��Z�,J��&�J��4�}�|r�g�+����3o�
LJ�%�h��T�{N�BM˵�O)��f�⥙�m+[	q�Mϗ�x��:���"���]\A~F	�!�
j�Mf�	�~<����0T��tG׹ls�[��=7_��
'��h�����F�B����\+�c��Nb�\��^uϽ4�f`��1!��M�5Շ�B�l�x��3������7آ�#�%vSzc2P�Eo��u�.Am���s6X��c���C
1p��&��~���	���8�G{��rc7Π<}eê8������p��@�G�D�sP�H7Ay?��;Ef*w��"=/K���	4����d�yf1p�5�)^���V�Vm�8�'rP����K�'8�_w�u���Mm��˲n�y4�ɿ�E?;u;�
����D�7��~��)=�\5�l�V�-ۢ,��<v�H�7,��e��:��Ԅ�я�d4�\RxZ	o�d�jm� �������\I�4����?ܷI �D m�bJ��{PB����D�w]>}&�a��(X���_�ԕ�	�V҉ɇ~u+�[��7���۾���7,������u�tž���3�Ő�D��N:�2��=��
/�D����TE������ț�n�rT�����I�'D������ܝ�~e��|�h���L"�f��B�w�O�\d�8��?])��6m�ǹ�� B��Gҥ5�#v:���,���@3�Ϣ�B�nf��ȅ��j�Ԫ��L��b�ÿ�ʥQW7���	ֿZАз�Aң������uP��#����=Q���r�b����kJ���V�߰���L��M�$e��j�.%N '��?}Y�NՋ���@y{ �����/��(uX��7�ƅ-T4{K��0��t����£y�(VJ����VLJ��Yi��v)�š�p�;�����C�@�v�ܞ��`��uC"F1Z�c-=���N?�.s6�F-�p����.�e�����`42w���!��4�N���iЂ5�8O[�PA�[ď�/��5P����<s����!�?p�ބ���n��ﴁ��&"hZ9lN����-WO���=����MƉ�ۓ��(J��-��{���5�d6P��\/iJ������A.:n��^F;mL�ӯ�%��y�����z�`�^Z��Xż"�z%��'��"Ed!Hd-�`GD(��a�*F.��Ya	�Y�沦�W���~�����[����U@ʦx�{"�ȕ-�����-��t�O]�˩@��8�8�W�0��Bʬ�x�ҥ���^dGU5L��?�Cz��*i��1��O���XCamW��(ذf�@2�DV2,{mYt�����8-��{_;��mFAK����ǹ;5q�I���NX�)��We�ҕT?;��߽r$�;Jd�c�R�x�L�� �$mU�s�nݱ�'@���]ĭ��q�5�_���O�J�"R�\��{e�O#J�/�c�4�r�Q8��_^��2x�P�c�PU�wF_nb���>�l�'Ƌ�"#�w3o,.�r������.S���-�E@K&U/��Q�0X�{d>�y�?��"�C�!d���\3Q���(��L�N*�\ϷKd9f�3	�4�5��nn?u�ԏv�2��Ul�����l�Ä>�}�V�͉S�/G�}�c3�q�!~7<w%�i�h����%�x�¤hv�9j��	[�>U� ��(�P���~���K��.9��r��Y���tJ��t!����R�NԺ��%�\��w�,�Ş�w|����F̈�"��}m��.��;��X
O�+d�ó��ѳ����!UN����34���P���	fD*�@��[�tNNk�3�z49
-�.6]��tj��&�Z�e#���
2y�(�Y"��
y(M9�1��)9�(�fP�A����6���81��*n� �HJ7kqu�R_�m�=߿SL'��9���8�)L;�g�b責A-.m�x�q�8
�2x��S�"�l�L̫9�tf���2~�*�X���u_��Dx$��1n�G+��F���_�h�[�|�ᯕ�r.�.u��?8"?G�yR�&��L/��LX�*�`��K�6Lϖf9�"�ʾ8�\p˟#d�B`���x=�8&��ݟ��J�g5 �A���=[j<����Uz�g�Qՠ���tq�L`gt�I��te���n2lc�����_rwmTF���8������Y��HrۭXw���ϔJ��f�;�W����6F��B2��<�ټ[�O��+~~�x��l�6��
�xF�L?.��UL�o0/����v�YJ������S&v|�E�r�NY�^�cx�M���p/	���	�����s}��Q��MQk�~n�B���&� �RU�W y��o_�:��f�:G���ou?���R�u|y #�\�!NE���� �M�\ꋙ�B~0���z"0����ւZ�����gk��R@2{�B����4�T���.�]��t�O���H*�ɘ��y/\[	�������w/��^���3B^����K�	�R�����1;H��
-�۩�7�F��Ðc�>�E�[ř��� OO����7v�Z ��o����"ṝ��4�u��j�f��Q�����Bf�p���8��z6�낺1�g1_��d�}����k2:�u���2B4��yѐ8�.[��ʧ���W"le��(4��M�;%D(�W=`�%vV��۰��K���"悽��Ѿ�#Wǿ�GS�A�@�d��g��S-�4F�Q?v�Ng�u�l�X�([}[��}�۲]	�u9�~Y0z��� �d��S$O��q1��}�G%Q�K���,N+�Ϳ�?c��S�`�6�Mm�I�'��/>Ʉ����)�y	!��KHH�'.��w��5���j
�-q�vU9Z��#��i��R�7;�\�k�9\a��k(�t�\�(��N�q\�+���uz��O"��G�5�T�l����Ug��j��� $����uQo�  �J��hVP���'�-��)�����S7-�0�I������N�-���i���%R�p��{x��m�9��d��U��?���"'��T+� �lƩ��=8�j�ޯ1ٙ�Ge��Ts�&��G���9,��sZ��2Y�;Q=EE���2�q��r��-�Ǎ*�d2�S���-��{"�do����;����BƷ 
�H��#	��hp�H�6�e��];c��ϯl�e)�p����.��m?��ed�bESr�JB/�͢?�D'lp�cH���7����3Χ�e�L�m�A�dMw4塛rjj�]��pRɂ�5��bcF���]������U-#E�z�؀	��ܿ<7�|�R��0����%.�&�EXk�G�Onf�A�����$�7
g�[�S����,L���t�䚻*�E
V�,Y��(ϟ�jmJ��F�!$��I�o�-�x�ѭ�g�A�%$9�_��ф�|��`,.��Xȹ����n�Ȟ�A�]ɐo�;GlO'/L'�IX�;��v!x��o~����AK9�H�1
i�]=� ��`�Mc�$EKo+�Ҧ�KMf�Bx;���u��is��tY�PNJ��Eb?��Bі��V d�=Kq}_�h.zդ��!���P����)x�����"��]��8��o�Mݲ/D�W5�0�Y��B*W`!W�ҍH����>����{��)�R��)����j�ҡ�x���Q��ou�S���<:h�y��u���?	����Rv����!Q�a�%P�鬅\��[�㙴��4�y����ΰ?ښT��0�;4��(�ުѮ�)���@�Ō8��:��]�/�+��-�̤|]�SoLDP�o�w�UL�4��
�xg�h������?��n}��W(����Y��jk$\�%���.��J�G��Z��@،6Qґ���2l�x%�JI_B	�ťR�`� D���M��s!��H���G�����4�L���d���)
e��W�4`1���B����[�%ј��:z��	����
��2�!fP�mg�~�U���z+>�mƃ��t��4��wt�๮�sEZ�nKQ'T�g=� �O(��v	F��ӓ"cT���������!�Dꝡ}?�����3���S��D"�7�=�v�p{���;N����#��z�o;�.�*Ԑ�"!wv�4-c���Z���e��C)?'�t��W>�)��x��l
����� �e%��g���������\:h�NO�@��kP�ij�~�t\8�8�,:-E<���9 �ބHE��]���
������JNY�yETu�F�;�A��LA�Ej?���19�C[A �Ӻ�ۗwW�n8�F�
��~�Xΐb{\���y���7���O��o9?���p��MW�H�+?����ۣeSWaCPh��Uks
qk�-1q��Y���	z��||n��.�3��U󧇲��q[�ε3U>�f�Ŀ�S?����09��B�@�&=����1K�y�H�]�c�+Mt����S�!����pW��sz9�|*5��\U�1�m�ݑ��V
iAav%Ob����9��ò��{�{[
=��L�ض���H�zM6 ob�����.l{��_̔����ŌS:��ÿK�&A�
�V#M��^���]ҎM0�1���b%��%�z���&.r(���m���$�uP}k
�A�(Kj���M��դ�(����}#=�]��L�+�KYa\1�d����g�g�h�+v��0$G��o�_%4�����O12����^��TS��z�_����H��|�L�f����0�������y}H�W�֨�}�%<����U	9���b�`���[�@gx-�+��'%�;�#�|��q�li��uꉻ>������m��%���B8�������U�p�.�ޠ��L�a����|�A,?��_�����uR�=�B���[��q�}�]��KV7'4N���@2��zڈ�dn���rj��H�B^���i���0���i��I���7nv�j�zK3��K7�@C�uU\-�zho�#�^������
`E?��D$9b�Z.�ܽJ��|��l�b�5]v����AS�*�dJ2+��0d{��s�dg�xs;�?3[�zZr�-�j�G�>z�A�����o��j����Ϸ��Y&�Vڨ�nH9V��[�D�Q"�)��fp)�r���(���N��7;}q'.E��:w��72��n�V/�9۪��C�p�a"��8�&)ٜ!�4�V��,*]=o���c7-�k�z,Ѥ����--��Pa�OR�m�J�Ф7^W
��1,�L>��`�7�2e��u�t�3�o��<:k���.<��ɗ���;�9-qbwG%c��.�)�($�� �:U�Q3�eom#�p�bCVQ�&���1p��ߑ2�#��	w��b��7(�z�?�	=�@5���<_�pb�Y�Cd�����N��6�9���EE����1;�׮�ڑ�~��9�Z$���R�`n����xT�^a�Q��[=@�����ޟvx�H����-ͧ
;�s�����⽉�@��@L-��F�b{�޹=���ѿ�c`>hZ5�K+�����Pm�����M]ٽ��E�\$���n0%�9�z�Ӥ#�-ҹD����-&p��|��Q�n;��I���,j�󒩮j��GZVm��Ob�@��d�����Y�K�����S֛�?+��i��C��Ǽ���L���)z%�@^I`�~�2xb�Iޜ=���V蘂DePrAu�Y{�U���H�*jT�o����1ܵ�@���^M��T�Cl�j'�N��ZY
�Y�F�\�)J<����H�n����6Y)�1~&���H�h�0�Z&����?����ɕ>��.l	���z�#]�#�;9Sś(�����B�Ds�"��E@O ���b��D�^q�/A���e�z��	����� �A��Q�}����.V6�bυ������x����V���<Fh����SJ�+a����~�����P��8�n�m���@����jۯһ^zF����b9nrB�����K�c��ۘ(uvH��n��A�q�q����4s�X���E�ś��q�E�������)��o5�O&�����m��+`B��vo�: �����>K�TC5+�h����L�Q���f0�n
��+�Α��L&��+��W��Bj/mX���
�0�=�oX�;�ݦ�1�-ɲ9��q�6���*pX��z�����~a�!��)�o7nIV�%+�p��}�rf�&����a�3��ﰋ��4����Tm)9	�\�h�G*5�@�
��j���d��rķb1�u����N.�4Q=�)�F�'�k�x��}H:��KVhO�%
�:��m��98Q�/Z�(w�˧[B�4+�׋�f%�|@~Ƀ���g8"(o����Z5?�}�}��>�pc�}E��V<���̹���`H��S��٫�N �x�j�6Rv�
ܵ3K���!�dT�q��=����(c�A�����2m���������CQ],�9�&FP��ڒ�a��[��(�`	�i�*�T5�\>��_��v���������@`��g���f�5]s�jSqO}m,`���:i�Z�Z�h��g��?�wW�.R�5� �@Z;+�<��(˵��?ڌ�a7M���Aa��~3߮�:��A��e�,/�����M@��ް�~��I����\酮�ָ���b�:�J��oJ��#N�o��9��U�s��r��Bg��mk�N�ex���D�����E�ļ�70Ja�L��?��~�D�k˟��>3�wI�s!m�W`u�}�׼y!�N�N�,b�����*Y���,+'���F[3=��5��SQ�W�ܠ��Ӹ�y(:a8��"4<z�(69t.&�]r�b�����GB������y����%�R��Lwy�@�ic�Q�7�)�5�����,jI5O<ޜ���	yWV����J1T�QHX��4r��>X4L���%D�\����9�:��F��~��a)�ΰ�e���U����@t�D(��gϳ=$���.�U^- `j���������h]�V�=}�&���{|�EL0~zzB��F���7eZ�l��L�l{k�����\7�϶�����s�����z)��X���D]�P�g.���Fjh�J|#G~S�G� U��o)�(�ֻ�E��=`��n�硭�bT��?Y}6��A��̓^�R=�@ĉ�
������W��8���L`��>&a���*��T; hzF5e� |`R컈,O�G.�� u+^m�m|�BJ�roԫ(&�e,�_RfC����C��0�y[5ZtY���v������{.��Һ	s��x;��1!������u���}�qS��\�`��+�6X%B��a�&���#��(����RK��J'�v#�j3~��T���Z�;*�[�LLV�Pu�M�ۅ ��~J<v�<�i���˺�o>��<���^h�P�������59��,?�F`):O��G~L�L�!�Ǆ����� ���$g��t����u��n&��N��ƢIKy��@�\ꔱ����Ϙ�p�������se�`�slx�4�K��4�}����m�F��_�L4���>�L��D��8����s�s���~�Ag;���ek�K�y�d3�c��1��S����a]��*"���L�wW�EĢ�@��Y�Z�a��'��B{����ФΖ�����Sձ6Ȅ���@�(�Tc��}��IN��ݪ{�:�N��^ta�P𖉮v�,��<@~�#T����XjUD#B����B��ze�
m���<�l�_R=YgxY�v��k�~Ҿ(�R�T���{��������~(Q��K�!���8���%7T�2�fd~��$Os�E˰Y����y(��;5k�v�	\�q쫩P�&b�[Z=
I���4-�sb�n�kco�,�)�&O>V�*�����ս*A����ȏ&��֕[��݌{��!$�G�7�"TU���S�l��S�Re�N�O�"��O��	ݍ�Z	���݅G,C�d��h~x����޹
;�C-p�<q�q-8WR�Tx��{�,��yF�Iq��j�e����b㌝�=A����3��?;�)�_���[�����$��'��H�����r��j��Md�;X����t�iG�Qׯ:��H��"��oL��딅�ゐpPw��љ�r����?�W0t܁-�p�F���J%5V��fA�0�8e��;%BM�CN� �V<:���5�xT�@z���
���$&�$��/PU�bDN}w�?V1�'�߄o��S �56 ʺg��s���e���׳>�F?�� +Ug��`1i���<,A����rb��uD�����.�q�����_�I\}����+�ı��C�k�˖�#\ܝ�j����9.cˢ��B[�[�3e�u@l=��`�� ;>����:<^�	�dL�&��o�G�ߵ~��𮟬�4_y�0�{ W��l��$�Ǳ�P��@��L�b�������׺`�G�~��2<w���bU� 2ޱ���f�?���9DgHhjj\��|�@��m�x�ʘ`���We4����6^�_:��_��Ŕ�NA�	/�w��7�*�p��M�o����c�1WC�jp�X�9 �'�F�b����9].m�iߎh�����G�i�$�LX�sҙ�u�[ƾ�|��^�:47�=�@���`|"2���ňl.l�8�p�Vۉ�x��b�	�@���I�b9��k����i��LV��P���@o��3��O���	]�PY'��a�G
�״��ԢE�����U�T�d8u�^t@a�ٺ�PV�ɨ����|Ĭf��j��<m�Qu���Lv��:7)���8����n�q�Y&U��T=�*����'!���)��6@����|�ʿ��l��6�߬t5�e���}�)�i�2��"�s�s��!��@�׊��m���TF'NK�x*�J[_���#(������NMx*��M������UW�.�S����1�˩%�,Pw+��~�B���H�Q���]4츤�sr��k�;��,�E�ֳ��1f@}Ѳ�r�/���y�5&d'7v�x�3]����T�M��ؓC�[��M c0�y$�P���� 2����~C+8���7�T��E8�H�L� ����n&q���X9?:n���u�����[��x����6�þng�?-�>6�YF��xG�����z�ٷN媥�g�j���N��dl��H�_�]mb3]q�ۜ>��;c ��=�h��ܛ��z����~YU�w�?��%;K��S���3l R��>3�HS/�$���	�zi�g#���gb	�����s�:��kZ��{l�
q,�F� Ա��B-g��������w���v���*�H�Bn8�0@t@u��{�ٛ��0�������d��2ڊ ~��?i^�u`iYL��3PT�)�u����fo�H����*�B���s��|+Al�G1Զ��_���~���=o��Ř�0|�t�0�sT5�r~&],X��>�,$j:~clC���&�(l! ŵ(y4���	C|٣ir����uЁ,m�˜��)�g&�ǥ�}��9� Uy�_2�A*)]�~��R�ں�H�q�0VQ��c'����:6!O�1�K[����.9�aWש�K�E]��|�����x�G��M�d,CF')��0�����K|鮞��UGR5�]c��k��݊�����Q`�"�<��G%.�_�s����+s&���	�T{���K��p����B�Z"�fz�X-��5��C:�*�WB� N�#�2a�7?�Mfׯ�T��Qh��<`D֍�)]�ji��=IƁݚ ��[��QqW�s��!E��! o@���ٔM[����ß�P��h�TѐX ��oʼ'?�t��$�� 
��7�H/�Wr_��0�,p�-��יEn�T��rг���8/��H��b�NM%��#�7�����Ӭ
(B�*~����)s�N$;��Gj(ո�fky_f�ri���u�<])��_އM���3W<ueW��F!h@������䘲k[kF�T~�O;�E!jj�uZ;EI	@��ȃ���̹P/��y�kB�d�b����22\X,;`��a���ԧ;�[UGU�;!��rXV���-=�dRK�&�~�Z^;��>o�X�4��4�J�FRv6�����P���(�6�V�Z���ut��?��a��.F�õڤi���+ɖ��_���G�9�u���W�n����iƗ)��/��G<�W_1j�<m��(QQ��1�o[G�!nMwr����^O7��9�^�)�y���nO�_��Q��������a{ye�Ʀ�a�?�|؜��f�7�~�ښ�@!�(5��S��7������m�6M�P"��Vhz��>u6G/�	�n����r�qT�꽶�ڿ�������zm@ҏW��������6	j���G���GQ�N�8��5Rvz�)=EPҺ!����k���e���L�v��d<V���d�G�|x6�k0�c��!�*=���&�5vQ���Z+���9��Ο����]��@`EWh��Qz�K�}�����y���d;I��7`ha��+�"�?��ڞ��뒅P�8&
���[���߅Cj��0������B>�XV��
S5%~o_fP���*��������إ�O�t��>����1_'��i�z����V�F+�w��٘\�qX7~�G1��ڳ�_#g�O��nVW�����J\Ph�'�%����k��/g��I�B֋?l�^ o��V�ǿ���e���u�����"�}DJ9.�5L �y�8i^fg�>ڝ�Ρ}9w.?4�AG���"ۆ�(�>|�f�2�`�`11}I����,Ȅ�q���������~�v�,�,L�w���'j�h�*�	}4���x�g���n�,c�mՆ�����ӆ�%[�s֤����|�� 7�kzsD��=�i�x��Cy����~5~���D@�T��[�~0��`֥��޾8b a��o�G=X�g���P�i�J��f�Ĝ�B�8���S�G�S-K���c:5=��ZL�J��T�.wh�`+]!�1��f y��Q�z`i��:j��*xT7e=��ӿ�����s3�g�z>o˷���
ω'�2�� ��a�^t�ʗ�ӳ�姒aZ'|m���D>FQ���Pe��fer�0� u�b"^p/B=���Q�|d*��|Ŕ�k|�nZX8���N�i�C����7n���S��Inb�݁s���&"�r�FΓ��$��C*�[rVs��A+i�6��x!
�I��?��[b7���'��ku<06n��uok�ϟ,x_�1\��1ϟ�&؆f���#<߽:�H�Tf��^j��Aܻ;���I�n�&��,��2�|G��E�2J^�/"�z1$�/$_eu���/l׫���\�����#�-#�H�v���]<q`e�~����$6M���(@}���X�<�4(��W�b�2��qcUl�q�L#�@jQ�X��f��A+q��&�'�Y���}��a"W������X��3����և>�B/��|�m�Z�7�d;�O���D��a&ІR����������%�&0[!�1Y�w7�oެ���0�Ic�u���D^�G�F��i�!�-讑,�P���,RA
o܍����{?�`���V�����;�m�Whk�>�.�r��XeX�*SyBU��{},r���<[�5ά~G�$f�d���t���V �^��	��!����=��4��s�?��f�F*�`:���#�e�f�[��Ɔ�6�n��kT� ���G36����w0;���/��i��RL����B1HD�͝5�͂h����I�Nu�
�`%B���bi�ł��C�䦵��͈�|4����B�WZ���?6�X�Cz�X�l���o܈���n�L��s��J�D�I>���_���h����E�z����Z���x�b���أ��K���9 �yGC�e���EpN�B�����h�xp��ũM��[|/�/��)y�Nڔ�σY����S��@�g��<��\�e��t�����%��kD�4�NBM�<�� ��:$�Z����R�J������~�B��.3gt{G1����1���(w��r�#�!�=�Jϰ���*�nҐ0M�\o��B�MSK����w)��W IĢ��@��M&������	1.T���0���Ż��(��)pC�G�����A�� Ҟvc��̎ �|��/��R9������ʴ��!|��5Y�ʧ2�+>%)�Gs�=>J�	�daO:��L�A�d�,=�ᗟ!gɻ5�X�|R,��p�>J�+~(j64���~��6e	U�
#{<#�f�ܟAA���ǄQ�����R5���LV��0c	���?到�	.;i_1QC�W�H���b���j�(����Lٗg4z��@�|��W���6����3hn�X����J%�g��u���R�쵚�8�W��-����r�)�<�"%>�z�������^�. {09w�.*7��~�����Po�v��)�} w" 	���S؛�(�9��|���ؠC�=��XtG�}.�']��Lӛ̺gժ6�y�]=�PC��5"ݪ3|�x��}Π���֢�^�U<p�����Ћ���p��|�r�,�b ��,�"dK!�I�Ũr��8�4 ��?7D.j�D2��/�^��7=��Ď�N��۳q�����vaI��i']�X� i-�;�������<4���/%	^��Y� 	s��b�y<�i���@���۩����%x4��N��P��m�]��V]�'�*�u�^�4����a�\f��'���~���r'�����إ2��h��,�Zq3-v�B���֜�#��D�eˑ���W�t}�)( �xF�?�$��$6?b��#ԇo���Xhm��ߤ�f:�D��Q��N�@*������gѢ�R�x�9�)C���@��Y�"��������H�W���Z��D��_d��+s����]� s
yFq}0^�Ƅo�N��	�m�;Q���(Xw
Q��{o�Əisz�HS�޿�"/�R>/�u�<��&@Nm��f.p��h(�
�M���p9D����c���2�2@�.v0LT}!�P��E{I�]�ۯ~���8�s��XQ�K�w��J�&�*Ə�}h!�p�}��-�>B��S>hU*S�;��WVaj����Sf��?6ِٝ�z���P�e�B�a�#����ׯR�}Ul��F�M��길����o6�ۍi�S�R�ʲf��KT.=�Mp����6�r��j؉2�FiN�����/7`��X��%���(U��BQ���`%ߧ����6�^%�Te��N�zdL���L�Od�}M� ��>zٱ�R� ��V�f{������&Zn�A�1AO��i�w��EH�ƺl�_�6$�3Z�:g�+7ʿ�?w�'��1��tV
GIo�����J̃y���ލ�I���K���FyCgF	�%�+s�K�l\��l��7q"�tp8���Ha\g���t�55�����*k�B�h@���c'v
���X�f���l�"M�
����>/5d�WU��+P�k]�D�L�8�('�p��}%6JO�.�P�@�E1<BNh\hI�Ң��|Ԓ��C��;��+
~��뉟Ly�3��Z*��d������_�[0��,$�>I�3V�T�q������I��cL|�qmȿ'Խ<�8֪��Q�0����y��!���?�ZYk�)�
u�����+���033�ʗe�'��%`X�5D���7�?
�.d?�Qtġ	}S=F���8���ޞ�r�&��&窆vm�=blqKyp�Kh�@��r��Υ��uG����"�qO�,[ע=��zE�GK�ds
�Θ�zl(���e�#���"$/�ƺ�_]h����>э�����\������#��1��z1?���	�q(�w�8��̴�6�^��n}6%�5�b�0�D�.نp�� g!+X�u�;�����KB�B��l�w�z��dw[��"G����	w<Ǔ�.UK-�r������z|u0�)S�=��
uR��L�R�T�tH.ю��
9{Ht����Aq����*T����d�T*|��Z��/TmK�;��ɫ\v�+%/Y�]��nf��)ۃ\摒s�����F�	´r�����:O��; ��C�I���UEN�^��T�2�E�/ Z�����c�.羡��

f����.��*���Z�Q�y�HZ�$�
4E�8�Qd��pUu��u��C��۾PU�����H����t\,r��+�L��['��H�P�k%�0,��^��g$��q\NG��:\�J��1,t�q�	(�$'� 馦���'�7>����]뮮rޢ��	�W VN��� `h�=}.�?me)ѥo��Æ%U�7b�yS#�L�+�cJ��ڋ�5$�c��vl��'������P�5�)2\躕；c����]|����$j)Q	��=���U����]��!F�Y,	d�&���Oc`8�!u	��>��d\{�R^�z7��}MB���n��JF[����Qzށ<I�O���U�<��]�z1�Q*Z��̒#�g�����C� y��+�[ʻ����ˊ���l����\���qO3����hW�tm��V�W�z�e{�Q�tb���4�ߖ==Y��t)
Z�8:Ѭ*��
A�bp}Q���/�	�^	[h�Ara��$>����LvJ=x>[R1C�S°�(�� �`��N��I���7��g�*�X���tE�9�>��[������Q��7��O9�;O'���F����}�8�i/G*S�뵍Qp��J!KN��;є��TI1��&tB�M�	26��ݫצ�L���k�˼�j�������Z�!t��w��g.�����Y(r���+�j�V2�
�|M���N]���:ь98�[fu� ���]�����<^�=��R�]{���e��y�E�c/=P�e4aU߇:�U�`�fv����_	��G0�T"�lޚ1Z/m��荐�8a�_���.�yq����g��r��A�m`��ڐQ��SlAph�o���>��]u����Z�""!L����8���o:SfR���#�����C����f�����j�Ӏtc���Y�:�/�Q�-o���ID<a������k\���C�=�/p��Z���B,A
2
k����X9�)OQ�&
�����3 *|`�X�Web���/T\3��ˆV��+�#a��Uz�XWH��݈[e��2��hB�h�7���0�q�/�����B��/��I��d�y����b��L��*;�q6���2��[W�i���-�q���B����zh�j�:�`��u��M|�ez6����E�\h��Bꕝኑ���8�ΉaɁc��Z���Y<�,̬g7�:FxX[A.�(ȵ��4�e�?_�����c&�DH��2~j��)���w��Ҁa_�.����"�[<=F<�"�Ju�З�;���F��D��Q��e����r`��x�ʿ�U��-��x��$���
���]��iR��iD�-�~[���=���٩�l���M��C����J��p�o��?�M�}S�n=�~������v���K���/`�{��T(ݸ�''��`�����&��FD��M�E*�&�`r��B5�7��w߯�v��w��o��O[>`�2I�����F��<4#�Qp��L�U���&a?����x��ݒ��[w��&!4�+�,����*�Y(Ε�H;�D��3nEmN�g!m�~t���i�нJ�
f^����=B���C��h�����n��ǡH�B0g����|@���`�ԘC��ů�L���Z����? Z�����ƌ���!A�%���Z��s_w��񿅻��d�Ui:��`��YI�?�$�"j�~�{Q.=�7��."�wÉV���������������8*��?�p��`�M|���u��-ǀ �՗/{]iM/�r�S��a �bw��by$�$���f��r�E�l����W&q�<ZW�A�������"G���T0WQAv:��A�bS�4�}^��ۥX���U'���2$��W������˱��O/�%փ��<q��p��p�����>�뽯l�k����������8��M��|�jƝ.e�/E�s7'�x���j@�Xxh`����(�Y�+ƛl��$�O�+\{��S]������=m�4O��uP|�����
aص���m�%���(0�*TA�my��[�=l��O�ɯ�G�g(.Y`}�-n�1��j�,��^y�sJ�,�K����56�b�S}̭H�gxN�i��ߵH}4Wkz�� �d8D�+���nr�qxvu��N��[���y���H|���g����AfwQr �;O0X������ް�@eGҧ�^/������?4���%��I��֝D�;{�zl�a<mȯz"� �#��GKH���|�Q	�y@�|�xry�v����GW��[�D�5��#����j�O��ETOrz��b�X��'��C�%o;�Ig����`�96{}��	���MlTBvodF>����)rK�=��:�Y�Y�MB�bL3-0뒫�E���݌�D$�u�ի�?��7����ӻ2鶓�r�8�Dв�F�	R~M�Q^���q���f:��	\+x2��(<BJŔ{�M;�s�D���S���X`
Q3�ٚ<1�-��=C9�t!�yt���:U�f�o$�Ծ|�Lѱ;�v��Z�
���3��o�K.o�؇1u��g�=	���ZL6r��_g��|Z?z�nډ�CB�/'��L�N�q�a�UG���{x��R��I���Õ�HEe��}#�K��:���u���>�R�΀������[�Yyĉ.��̀���si��|�?R������w!���H��:d���@�o_>��嗪���k͝J�H��)�!�\i�1���_��sPu������3ɭ�<1���6���ƅ�/tR#�s?=b����JAH���rE�8��`[�>ܜ3I��ɚ7��#o��W2�p.7 p��[��6z֣(�<��X�ݖS�k��H*��fx0��pC��Ky�9bCQwy�q�>d�Y����G����A��b�i2-G��u��bm,U��[r��NP�ҏ�L8��c��Zt1�j3�0F�CٯpO(�ֽ����&�ծ@klG�X����Ԉ�ӏ�p��=/����*������и������*^/U��rU�L��k�՘�X�_)ٴޱ��aG��z�I"��U$��=�4����啚���
�Rn�$YE��2�V�^i ����@<@wO�i ����$��c�Q��~��F;�J�����eP��a�4~W��aχE*댘�1� �UQCn`A8F���2kw��X���T;+CP��7����f��������eD8�(�ᙚ�$hKK'�d��&A�_����ȃER�/�*UG3����L-�.&���D�H��l�Sӑȝ���(�`����9Ue�%�nL&>9b#�c�:;����L5��0~���� o�"����<���A��tژ� ��V��J�#O����D�h��	�{6���@-�b��]y�Z�{��.h~ORT'�,GqV����О�N��(�i7�I� 7�x��2#1���.�@�N�s��P��$�5-��1o�]�4���t�0�����q`ŋ�|	W��t����@7�A�n�w�j�!��0�=Dn�_x-�S��N������2ߔC�cJ7���V>:g2
��U��Zxcߐ�s
�!@G�Jvx��wY3�����le����Gd�(��X'M(\<�����`���+���d��pX��U�%3lc���:s�c��E�&��g�5�H��/�c�˼�wY�4Uҥ%T�KIUR��W�($���B_�h\ad?xOa!��=[��?`̖t�1w�nM�)d���c��/����bg�G��H|�bxҸ8���;J|��}��	���M�LZJ/��>��kZ1����
�\ ވ7��g����1�%�*���e~G%��G\�Y���o��ט��v��Bp����H�}0����B-�`�|����鷾���=0kU X�+�lMd�y
��Tň��Gc�˝����(Z������\�EL��M�K��r]�+�Bi8�}��6}�,�7���CZ�9�s�|2JY�-�L}"�`�wDH,�ҡ��(��ꦕ�~3�T�Rj�3x�&8:,`�M)���~�Cp*���֮�z��+���b�H��j<��g��m�I��_�o�0���W�G�]���jL�"��7��Ϩ�{��7]�c���AГIn|$�lD]tB��j:}e�G?{XI�����o����h�J��"�1q ��m�E,�䕃Uks�8���$3�$�M��9×�=����}[r����,�A_ }�do��냺*:�d��(�M7'��.Si<`^�D��;��'�V+�{&��{��-�5�.Z0��H�������%c`�δ������gan,rdv���/������d&+W%]%�'��#��$����M<e�uE�����H�SH�:zQ珡|���5{��E��~�[Sr��6ʹҙR�HJ���(߸:�HU�L�",x�I��V�II	a	�Y0
�V�{0��KV�.4� ������ZC[>Բ(�wj��^I^�Q5a��1�:�:�ºs��fq��_���e#�Ց�R��)����N��,bƂӈ�6��86>��ر�]�O��g&���1�1Ҳu��EM1��0��%��<�|BT�QF��?@c�6�����~�S�͋v%���I� |?>+}���51��%[&>Sҗ�v��0#4����+�*}��mC�pL�U�4�^]>����Dq���-^�6�f�q��}*LZ6O��2��Vu��J�O�����%�Px�oW�{+b2X�BE��
��j���@�|p�;l5�ʶ�.�,2S�������h|�<��Յ���t�`$�aWx��Y34	���Y�ٛT���*������,9x�oū�'���Y05e�����s�������B�P�YJ��m����נ�B�٤�U{��~"�qw�-�����p��j	Gz�9�	�l��A \iaݐݩ����1;�&���X5�t�>�j����C��/��	B��T�K�	��L&�۶oন%�$RJ;���F~�PXTN���*�}�:���|���	��}�ӏ튞�|��\�����(��b��@��$0&��8� �#C��"�.Lq�{���澮�z3�z�����jH�^�8�^Z^�a{�K�v���/��@�s�B||��� P�ɈK�0��
����O|�򏃭*`&�v����N���h��EДp�ʫ�?W��H}���\K�Ҿ$�$� �v��T$%5���s� A�O�������ɋ��V�޹:ǩ�K��T!� �8V2-�U&�(�D�[z������ZK2�wc�B�)���6�E����#s��@�ƶBj.���ԠX&5�%͡��`U�*|8b�.���i,C�I�ϼ��W&]�͇��Z�è����Vݷ	+aGP��AB�d��	�<�~�rt�� pIu{<-���) �����ؙ�K���K�A�Ư�~�!t�M��M�G!}\*,WF@��S�74.�(Q���>|(CS���0�R>h��(>�=Mq�6��A�},{a�}*L��_�)��sv)!��a����6��^Tm�Ԋ��d�>Pgp*��X���4��-ܜ��^�c-n�Ҟ
8m��=�_�Re����h���mj��<ڗ.���w��@�l��O��+������4�d�{
��p7���|W�cƨ/?C�S5(�:�}d��K��0=�bP�H���Z��6@�x�ϑ)�a�_m�����(��6��c��xn=��*T���^m�ڨ`�Źt�>�= �p�"�ӂԕz��c�D�mT�N44_C	]h�{ ��7Sd�CJQ�GhH�y$���4%��鱭�.ψ�k� 3��{�f�8r`#��4�^��MDh��P�Q(��;���V]Nx�q���N�L�����tk|�m�����y�2n�n�)��r��^�稍���N�MI�\Ե�s��b��B�A8@��!Bй�ȦK+����=�SA|�%�'����v{�sUA#�F�b|3=�C< B�gTt��3m���=��BP�2w�:�c\=�����E��uڎ,�/%���4\wfIN�Bi���b����~(q�[B��{wY\q3�w�qq$�Z���%ǹ6�y��VB�:>�6>��
�C�o#I�P�Kӗ��y�^!dY�5�i��S�O��G1����&m�$�/`?�e+�[�@�[m���L�e�Ƙ�BvT�+%�H�g݋�H ~`ԃ����D��k�3���U޽2U#�B�Uj%��7[�g��SzE�E�hy�'���W6,�� ��h�*9�1<:k	��� �0M��SL�I�1���)�%���``���wU *<���ȊV��r�M龨s���9,߇���KJ����u�K�a�Ȼlr5�䤀s%���a�x
�Z�aR�Rȝw�\��O�z'-ucG���[a�+�L���v�Ο�.��E��4��|���-�o'y�:�cW�|�F6~�J�����-���(vK2(׉��>�=�K���X�,�>)���1׎��-OY��cJ�ǩQԬ����o(9\Ou�T �N_���
�������)����(��>͠kA��)*�O�dbʛ�������c�c��~8���4a6]����m�H�A�I��� xYD�gW��Z�ɭ9ڰ�ĳy�q��%���{�P��N���U1�����֓��98�/���%5�_��/0��%'w�R���t:�D�����N-�K�A.҈R�ʝv�{6�)oG�A��9�}b\zmB�Ght��X5�Am�U������4�O�b�o�
B��>�ݢCџ����P��!J��,ӟ���Ab�ұ@�f86�T��BP�K&�3r*���<��8U��p�Y!��*>ن
�8��yZ9�?'5�g��>^��"�!����<�k��l��C6h$��E�?�"3.V#f�f�� �X��F��S�::0���_�$����`Ȟ��`�R���O�
Ui�v�+�`=���X��z�jMv�c�?���kyϜ;H�����-U�İ������@�٥�'��eh|�����(���U��؀�)z\:���s�t��rhYz&�T�ul&����f"a)�#��7�X��5\�'L���(S\OE΋Z����S�n�Hi���O�Q҂}�!N���F��ye ��,����4	�V`�|dwc���Ϳ�w����_�T����2<��ӮsZ���ٔqZۆYai 
�ΐ��uv*��@�Kj�@����kJA���O��0I>N�Ҙ�֝2gEc�9����ϱ��C/?��]����k���;����	�}�z5�Jad�)6����jو��ԉ"{'6�@�<A'&������E�v7{?,���t�H�B�[��X�,#i��yƬQ�]��\3So��|�_�.s�E��+�d4>-�]��vDB���S��Z�N��}�'J�JЭ�H�� ^܉)�o���U�kc�ao���2+,F�FfF��l	aD$JT����1S��Y�C_��,I-�ξ�1��>�8=%��/���)U�����>������G�jUޣD�8:��\g���h'�����w^��U���A�w�۬�x.��%j��U��m����͕��r��zd���kR�
�.��kS{KD���a���,e]?���B���x����w/��R�1Ȫ/7tUzJni��N�ր	B5�v��c�"���5wX�yd�HM�ih�@�(����~D��1Ԥ-����80�9s3`�00d@y2�<��|�<f�Gyd6��K�Ά� �"��@�3��so�� Q�E6R��֩�1�!J��m��ƅg�<��}�x���D3��$�]�HP�N�i�ʡ����}��&�Q��xF�]ؑ���k�[q��3&:��*	Ϯu���:����F��y�m�f�u
�E������Q���*�����F��o��oء��-���h.],�=?��>̖قG0���x�
��eOȔ�[1L�3«�v�jM�n�|�l�s\h�pw�ń�HŨ'd.zs"��z�W�5=i'Z9[OJ^)Y��j�_H�>���Ñ.ɟ�jEk*ٲ��	�?f�r�-��W�	�tH[z	JiTr��T�EL���9_ي��)]/#��)2���܌z��M�Ud����c	�f.��U@�GɊ�+e���i���9���D�H��c���\�K��O�,�hȃ��ݲ��o_5�pޱlg�~�����D8Y�@�3��?W�1:܀gV�y�׍	�:l��I��Y(I`b��(ECu�_��獥�M9!��=�
V��A��dp N�p������/�c��V�;|<��;������6���o&:��_s �?jb����9Zi�Uc?�%Ypg�]rZ�<�:H�G��caJؘ3�*�B,+�MşVnG�O��5��[�ɀ�d�&��iZ�?�-�1�H�ҳ� >|�mP�������)_��H͗��	��ti�9�j6v���ż��xf~C��^3'�},�J�2�
:�Ć�{��H�vT�����7S;�z7�4eC:���Fv����kqM4��oI�Q��eu(�G�\�K#��Æ�����_z�ӹ?�f�q��~�G�D	o4҇5ۚd�L�����&(lS�G���}���&����۶�q�ڎ^D��γ�j|���d�Y'͎���BS��ݳ ���-^������t�5�H��֨4IE�잎٘�5��S�V|o����[#E�<��~�B=�X�n; �v�w��*��V[�p����(�<g�מ�ig���3���KR�$]�S�է��R�e5��5�TR���tZ����)$���z��������	\�.-
�I<{��G�K��i`:��8|z!�}�^�e�A�Vr��1&��]��a���5v+(�[����� pB�`Q��pob�J��Dׯ��41�"�OPPa�tX��>l1F �	�v @c=6����Gm|�/�iKb褜S3e���5���B[ �zrP60:�h�.W�;}��Ӯ�Q81���U�bװVM�|CY���>G���Յ�)�)��hm�MY���n@wь�t%v+������@����[�_�I�?��5�k~����N���?Lr���a!�Z Z�p;u�i0�6 o���ú.��wr^�� �@���=��),v��T��v��Rꢊ4��W<�%ӽX��f��%!s�m��a�E$�5^	x����^���/��M�$Ae�m}�������ڜ��rO���<��>&���6�b�oh��(%p�q����B�����m�W��O`0@��L��EG�v�S���:G��>a�O�;��E>��`�ohaԏ��S��V�-�}�Y�)%W\�s�ܺ�u\v����$�������J�q>����k�3���Ǻ$l�>��l�������|�'�g��
)4�v�*�4W�+SPN�pXz2��t%n�h��c�2y�FX��;3QU6����w򗌡z�!�ټNؑezT�eH�,�3���q	�������X�
��U2��6M>�9Hڦt2�G�rAa<Bƣg17�I����*��OBM#v:�V�l��#uJmSc���6�����
<4��6E^�\�w6<S
7	�k�; [-h��<��D弹-e&<~ U4U���e�#�?gzo������5���}r�hP���VL�F4�O��s�]�SO���l��Akj��dl7���\O�3�lR?P���Ɯ����h��!��4��+����|lIiA�r֫
z��Z5r���l(PG�j2��
���F'ٺ�q���{��#W�j2Xp}��w[JMU����Ev#� ��F��&C.N�Ǧߦ��`W���mb�G#���FR��9O�_/�3@���y�x���
��h��v����>T[M�a0;�`��"AG�W�r��
;�;��e&u���MP��֢���L���ޒǣ�ŀ�tB�Nte�[rV��E�Z�M��+� ��
���G�MhpE�?�{�mQg���D���M ���a��b0	��
"���<N�گ,���Dgt�&���GD��D��]6x~BF��
 �F���[�~|�Ruq͑�a�+��9�R��w?�cW8q!6���^P`�lS��|l��g�4uB��_���>2�g?���?��X� lԘ�85	iֆ��+��DL%M������br�K�@6�Ab�:��uZ{l O��7M�X|�7̃��}��Xx���S�K��Tj���|Q����-�9ifB��iD)�'�T��@mA[w��H�Al[��)w6Fsav"g���=�wQ�.t��.5HJW��\'-�D�}wcL}�Fz����6.�>�k�4��c"ZFc�4�����r�VP��?�C���,��u����kL��/
��*��ʠ��+��?�W4���W�P��%��V�>���i��'i�J����1c%O���!��{�٭��oLq�Ѵ�Qa��
 A��X���Khy�f�ؤt�u�C֒v�5�:"�,K����'!Q �	�G�)B`*�ͅ%Z�
o��d'M�i�)?߅&Wad:V��᛬��ꮽэ�� �NM
���̂lٔł�u5յ�<�Y�O��*��
d�o�t�����<&bh�d$�ҺOe��:aRߐ�BY�1P�.k_�l�}�O�'yY�,��� �k��2�hOfd�xs��j�K냎�}�&��3^z�޼]$&Eܭ@�%�c�SV���U����Ҥ;��\5Y}Y��Q���覨�P���V%����%�������C���*���6���L�.?��Q]U&�ơC�5�msM�F���P��t�o���"��vt������k����3^������zh�N���9
Ur!���^|CZ�}7�6�+�3��fq��H��?����K �b��?~L��l(tZIM�6a��ҧ�͞�2��a�d��	_��:���w�`����֤��p%����`����3��Ǟ����ć,�m���ly�	��^���h�B!]|]
�����?l�\h��({����z� Ά��?��	Z�mRHPOi�ҫ�*��Q����7��9����_�͈=-��4 V)��X��kQ�^�3ݑ��td����!�#��"�����17'ڏ %/(��N�8���i|�,�F;�,�%C��c�`PK���(��
[��������=�kS?�j�ޤ�C�HŏO3pLpɔ`�G�]H�*G�ϔ�VmѺ]�M�����:��@?y����rB�%M�,u囗���a�Be��/��~)�2re��ȱ��d|զGDK�@7'؎R����R��-�u
y0�]�ٜEj����۰��%y���܊��D]���0J�n�/�R�0��3� @�T���t����o/�p�I͢�{n*^m2�Nye�禩3�k�3�'d����2(�ǂ�������0�d�[SP�i�S����Y�s�߅W��Y��\�^K�Z�	�%β��K�8�	��atm.-�*��f*�4�ã����vm&�x{����F���ӨiFIڰKS���Gt��-�����X��S�1Z5�n�/u��q���� ��D�"��"�O2>h���Z�/�p���H�.GYa�� �C�Pd���T:���r�� z���eTqMJ8��A��Eu���?$�5�������s�=���.Wm*W-	�ڡ�����&��2�b5�鰭�^衞�d&��P�@����#�@ebl��#����ΜI��o��n����M2,u�w��\-��;��c�������≙��Kr̔nj��(�2���c�ـS��Z���i���?s}�_�g�=�_��S��u�}�w�#�II�]um_��t��փ4ղ��	-N�_j��d��"{��?(���m|���e#� �[�G��`�:�m���R��8V=0�أ��T��OP/��+tmʴQ(g&���5�)�>�.���`�U�=�c7�Ï����r%�{��SR���D��w*���l�gQ��6�P���=�	�>d	�����_����P�ǧ��JП�����W��ʹJ9%X�v�1'�W�\��� K�j�!J˷+]s~�2y��KQZ�L6d��>��:��A~˕ګb�c%��'Vj��V�L�V��p�?�ӽ�s7?�*����7_���`u���`%}��\9hx�ԛ�������|?E�e�������R`ZP1?����ѿW�������J�.����hu�A�`� ��b�F7��-H�!q{>a ֬6��k���*V�ܳ"o0i�\Z��F	V�ig��쪿;�N���L|h�P<m%D��J� ���=θ.��q��-K��&��9�A��:s=Hih<A�@Hh8�1�=6;"	s��1�fbb��,b�@޼��L��A�alg�˝����*~W�2^hQ �\E�hG�j��~-k����<Q��̇���)�]3�~�^#�|�\������䇤x�E���F����2��F� �;�6�����˝�Y�j�,�ꊓ_��7D���"^�A
z��� �T�wF̍���/�d��iE�ɩ��⻙1��kM�	�2��ú4�z4�å[�b�Lc�oӣ����S�n׻�9'qi��]k�먜mt����(y&�E����9KW�B���3=y�EӃ����)	���������%�ì���g�9�CFU)B�F��j�1�3�tG�M��OVt���iS 1)Z�T;ciܾ��W#�ӧ����͈�8!H,��^�qk��k���\,B��4���i1��� ������@������Y�4��,ط�&!D���p���]�����$D9�}��	lFή���dz�p�j���p&j��(~6�vI1�dQ��������ٮ(�������~���&{
8G�t���G���`����	V)���4@R�ɿ�s��j�,��`X��>$�|[��Gƍ
Q8�	��M-���%�WlP�b<�Z
>�$�:���rn)��ƒ�;v5�z�PR�3���8�$��=�4F�*H[�l�D4v�p�y��kt�2�K[]�-�En��ŴR1*�B�R$��X�x�7�^ǱX����fU��۱�@�Ypq�u���6�L�tg����'�0&ab�!�(��Lc�����k^0,a:�k_j�C��c���@�H�/�)��@�5��qYo�0<��*.��I��ye�
��xV������-��u�����TH2H�.����7��`��/u�kk1���^UP-� &ł���/ܼ⼨�z���d�5�V�ً�?��*������n!���L��}�數j�r�-;2E���ܽ#��߫��6�v7����ňi����	��xZ����_��jn�c� ksm?�C��&ߩ�3q.� I�=�(�D��X:�e6ݗ6���>�J� ���O�i/�,�:m�6_�E �ʫ|�jJ�Żܩ�(4��m/Dԯ���t��g�!��Gf�ܑ8�!gE����w��:��Y�!S��u���������GNZ�6�S�<�L����JHsrK�e�A���Xs{�����q}��TH"ʥ+���f�(����F��du1xP�Hj�q3t^Ź��������HX���Җ0���vݻ�{Z�qi-���C����&�fU��K�:_�7(�ߒ�Q�+�Ov�{}`R%'��cS�I�K�����ǨМ˛�"!�O@� ���Y�JÍ�<W���KN��h�U�!�s��_���8mb;����sgb�m�i��ȳ���l�40����q��ܾ,�b���	����d��B�������5�ѽay��r�F�d�"�#;iK�u��ȶRl��b��O�+93�0���Nߘ�~����f߃Z�8) �h�Q�!�#��w�i>��¹�Y�DN�h&Һkt�ԧ����O���g_(�c�6���{^^zD�ޮ��2��I�4���s�&��@_&W�4�B�1t}% M՚V�3����q�ʝ�owP=�|A��8 ž��X9�/�҈�����29��#G8/�v���%�E�"M&���$[RU+11�\�d��$�?7�0����J�?��q|���z4���\�y�����\J��0%R��Z����^e@D�B�� X����e��E�||������O��x/�1~KmY�#0d�c&�FX���T�k,#z��͚�˘ѻ���T�2���4+�W�f��$30-��U�����k<cȶ�k�ʫ֧�v�"{Ym�%�}%I��M�&��$�i�jQ�H�gC�b����C��cș�k�˿�jʔ���j�؉P�q:���,�,֣�$��hg���`s�ɹrN�AvB%5�ߒ����`	� �.��p������ݢ���ş��_���F�~�Q����0Ǩ� u�E� !�`�)t� ؅�}�gߪ\�GIUK���������p;�]�����ۚ�?Z/V��*�T��U�ə>˴�g�������Y:��@�p��d�+Iw6Px���w�ŝ`ܽ��+�zMT-YyS?P�V��ܶ+x�ᆪ�*��a��=��0�_t���D�0�7䈋�[��=M��S	���p\̀\D"��;������r�����UH^���r������mG��8�g�C�����r�VxǌYTM���e�
+�9�s�4o:�5|y��������o��M�W�KFWo�8s���g�����F�&�2R�\�$���,��o�Kz��᠄�3��d6����#�0?㆙¡C�1��)в��8��=-����r�c	 E�kpq�&II�,�6���Z�����x��?~�+g<�!X�Kv�=ӛ��r�;[��R����/�L`�s��?Ezwt�f�}�g=t�����(E�<*�����Q��>U[��M2�^�0B��J��L[��tB���D��������i0��)3�f�ξ�W��+���u��{��ӣR�vw�I+z�lo��J���H��v7�Wy�!���h7�(�]3,�"LK�C��@�;jC�xq�3b�C]���%�[8	������9c�/�`�S"�o��T��ӣ��ۜ�/�rV�b�.4���+��M/P��8�k��O���i	�uЧe�?����~+F�fz�Px>�WM�$�{c��A.-����Ag~�x�M���-1X���+�O߄��c}�fzg�:�w�� D(�X���ؒ"�����G��v�^��Ŭk�RO�֊��M��%����|^���jcz-7��K�L�*(���T���<��6�of��(l�cr�#�M(~b�Mđ1�p��_~���5nN�=^�0FY�!^�Z��U�1S��~��� ����̦8��B�b|�H�.�b���3��B8+�qL��<���<��5U��C�O� k��y����C7F��v���$�r�=�����Ct��s5da_���s�Z���{�eM��:>�f����}3���k0/��pN+�͸ ������K겲h�U�s�<h��1�zτu3�����-"B3�t�\��!�eAv%}��:'	�ܞb�ل*?�lU���W��eꩻ��(�"δ��3�\j>�9�ruU�K����eA��������3].a1XWf �R�>��\C)�����7s���s���Fؖ͂���AgO�9���uF0�Ld'j�'Yg�!����%��9[��÷|xjA�I%���k��+aj	���߮0֧F�J6l�+���y����a��{쭽Mj���u�>�rr�i�`�aa㿼��*����vw��8�<����軴����^��ΝT8l1UKVY{���שi`��©F�(W�(V/�cl�G��cE*$I+d�y�''>W� ������Ut��s�	 �1H���K��=>�	׬#��/Ա��w-H��` ��%��*1U�X&ݬIH94�"�ݤ��������🲁��%$O1���t0������!=�v� �E������wc����٬C_���l��Ͱ��X#|����D�eL���%�,��:�"���1-!<JI����2g�j��9� ��J"�"�%������Ϫ��n���9�;hR0A���lV�.'Ӛ�`�ui[�d�4�m�ڻy�ұ����1��ԓ��miC��YƝ�?V����Fs<�����D��by��p����K�W�J��a��,�s�z<�P�J�`⅘�yp����5�AT��	��u��y�~�T:��+-�� ��N7���#�Gls�:��-���ԥQPz�E�յoe�5l�A�<ƽ�C��x=aJQ�?Y�h��T,�ꊬ��9� �I'�1lݗ�46��ߌ�Ǒ#HV��������K�˿Sa{�"n^;	~�t(���p�+ؒ��s��m��Oz�2P=�zg��2�[˭A��_�k�"D��nL�i����8d�[�fS�Qؓ�����D����]s�Wۊsp��׌6k�rC�9׻%�=k���t��^3�+�Hn&Kw�^d)�������z�ݣ�� "R籍���m��f��ş�A�����c�P�
�d�����\+	�GY�ݰ-�eʵ��A�\�{
D����T҉1�����Å@���FK8Ɠ��I��ִ�����>����N9��-k@AJ�)����O�3���mu�P� �juX�y��!����ͩ.._�����J�"k � )͊���3+;�~}V����W*�a�0b�S�|�F�I�-u8�ʪ�FH4*szZR�<r���պ� U�u\�L~��	��| ��O��,n$���'ҞM�e���+��8:5
�i��&oɫVTe�f��7a��Z�]ߚ�9���#��a)�~���T�O}�$uʐSּ>ó�*ʚ�
���T;�ԝ����̍�d�Z�q>�)�bmW�B�����ȹ�
�՚�@��ܭ�".���ts�nO犡.�Rr�v��T5�y�r/�`Fd����3�pS"����|7c4��%�=Å�g�M�/`�"�
2�b���`�G��X��F��_��<DL	Bױ��p���giW�����	�s2��G]сoN��4��YΦ5�0.vG�<ȝV�"�"�*��'�^�4�����dL'���2i)O�e&ޢ]���^�.��z@8���/r1p��#�{�iJyG�N*Q��FP�������� 1v�KX- �u���){C
����{��:�`Qȅkٮ8D���6��+u���WAӊ=In�ݱv�k-
� �O*BH/n�j��, ���ph�j��/H��98�W����4=-�	�0������
4`az|�K���11���D�v۵"u�`��MjfN��w�"m~������ �UXQM�cA;?�=	Z�bIB�� ��9�)6q��;�#�"Қ鱷��u�P>����~��Z�B|�]�/)����o�~� 󞐘Uɋ��-�1���v�#'�%n��f��K%W���&c�r���:�*q���������\ޚ��y�y�P�N��� ��������]d���.�dF�����)\P!��qf��1=cwS�39ƾ,������1�=�x�Ǵ�3��8f�R�@�!��߭� 	��8�Pd3ch>��D\���*~ �X������}��4�N���h�ByCԥ��)�Qw�\��t1�cjR�K@�]��E��yq*\�c��f�h��]i�3�4k�C�t���T]�M��t�^V�!諈B%�?�����5FO�G���������׫z�%���t��6N�ș�k:�cN�,��L7��u�E�*�O�{C+n��[;Ej& ��'e����V��� �V(�Z�����6k�2�^�Pq��ն���ä�:x\5�M,�� �]r�I8�~'ȥh ��o�_�r���������K}�a"-I�kz�O���X%�#0�Z���S_<1N^����`��3k���H�q0s�@�|ۈ�CRE)3�{&F��gO�c�z)ң�M���#���@`.lQ= �Z��c�"m<�j3k��/et�vM��ܝ�,�ZU�Rz�&>�	񵲣���\�]�1�� PJh��IZ�}��k!����$���_8R(Jv��;�����&U�|�x�lt$/j}����|���kL�p\2"_$i�aD�1��/���ϻR-Z/�_u�����|ɔ��&ABY��~��d҉��k�!sĭ��βׇ�n��g�v�&@5O���v5�Y^�X$���F�OƂ.���K<I�{M�����q���v_��EF+��|B'͠���x�7�e�E�{9A��Oc�A�Y�	YDw�4�Kx:Do��/UP�s;���RG����W	l���c�?9���tZZK�#�r����ne�4�*�xF��1
�/����-�`��<�����]�I8Q�����j�#�% @�?$#�+Z���D�,M��ڔ���F�1�/)OZ��^L�A�C||H�S�n<[A^��з���Ad��!�=����Z�N�� �>Z/F6��~�7\����VO�_�Q4Z�\j�|uD��#<˫��������%hi���W�[$��C���Lr�BL��0���W�`N��0�u3�W �U�߼M�;�~�M�?�õ`�%w������yx�=��+';�]������éǾ^�j;7��I�h�q�Ac�P=-6G�i��W�xU}�>�t�]!�@�{u �mŽ��<h�6ul~�? �}+�����t��s,D@&#w/�o:L�%(YL�n��0����auD��8��S�����l��$���^.�7�&f�1JǗ��-�m�)4�Y
>(���w}DA�Qޮf>��>aqXQ����-y
zo�'��4�dD1V�#���x���#����FR�ljc��v�8��j���}vN8�YI�;J����tP`�k`X���i�c<i�v�u1ݙ?˘�O{VG�+�C�E��LT�B�&:���(��*�3�1�k׾< ��o�(y���.R�+�'�R�$�\�3P���l��g@�[w��PĒ5u�b�K������i�
�g3w>���<��tO���F�^��n/����A�2�����&�AM��r�"0L���ƣ��N&�'C���;���x�Y����X�����Q�埚���C��]�Qx4j��Ԋ�^���[�M�	>?�G3{���o�yL�3���+V�k���Hr��o5�j��T͎�`=����n��o����A���5t�:�y�p�{ ���#�꼼�0��˭Q�����Si����i������ѩ1aug/nc+4�MI�ű� �-etEj�TU��b�H���zZ#ƿmj\��k�tu1�˛w���̙��m��jq)��;�)���*�鸑I�
L�>�)��돁`�_T���Fa6�Jy*zW�sJK��u�ܭ����\�''�S?[�t���Ӡ�X����0�zQp������r_W�0=}�-^��%�}�d���h��8#�x�;2W���%-Q��	Dg� ��L�0�`_q�?軺6�؅��0���rW�v������|%��гmW�#ٿ�/�� �+��jY�pܺ��G�}i���;��Z�v�r]��K,���'��Wtyf��'F�9�~���f]��޿��A�F��I
��%v��e��i����/ĮX��������p[��} ��Q)3����	bh�;(i	O��&Ngw����`����1���v�q4rzeˬ��`��Lpu����g�j/8�\&4%�E6,��1�ԅo$B�~�a*u�w�9��o���\k�~'���L� ��s"��I������\�w���2�N�6���-��г�����BV��p����2(lɬ�V<��߸�[�Y/3�]���%_˕e�˛��C$��F�ƙ���mĶ��5�:e��"��FӴ��,��WY<&kY��i?l�^3�����e P����C$p��ݶ�1��u�-��^<~�q!���V�V4õ#/R�3٣������ʏ����$���05'X��̈ �3��%�?�!t}��0!>�ŷ��8Z���7f�"b8ǪK(^*6ጦ�<��Z1GEǷ�V"h7FWlL[��,��ƀjr�x�]�>!DUH��B�
T-��}x�H��_X�C�76~uC�u�5�Ӕ�ْ�J��`�|XQ��]ǋ�Y�܈aV���)��3AK]xؘQ�%�В�ܢ�R��wK3�Vo`!�-^~O$�by./n����Ė�U��[��r�ו�ԣ���a�4���q����d�<�[pP�ow�+X+5>�Ü"�F����K�r�II���E������?i+�v�Rٹ&z;��ʜS���+p�%o�o��Sc{U�1v�9�(4V*/���$|��ɰ���<ho�
��BB�"o�iя� ����x��t��b4��Գz+�2	d'��b~�\�:6��|.�_h����)������$��Tٖ����~�w����n��y�X�u��>i�Q�C�qS�>�~(���Z��Fbi���<'��h�`��i�'�L���d;_5u���	! xH��%}����ly�&㏠p!���@�z��ĉb�+���N�P9 ��
A3�ӈ-j�5��$���`��\G��sUC;��~�tB��CNg�:�z��a�,3���X�&#_��3��؂#����le��PzIj8o�)¥�U��]X�d��pȺ��ˣ7{�*��b[C��h7�u��2�J�/u:{���af� h�wD5��C c'T����@�KO��SB�'��$�!�f`�ֹ��u�����}[�=�8υ\�}
��^mJX��=��l�2!;o�+��RK���lO���%�&�H`^zܨ�x8�p*#�@��b���g�8�G�u�1.1��ɞ#��36z4��\��=��Z4q����R�s@4�B]JZ�g����]vi�6��=�|���=�7� �X��J��.䄢��B�fMb�����7W٫���J͓���}5�5�Pe��`��uH�̝X��!{��H���f�=��"h9�j ��8��d!�P������A���*�X�P�����$Dy���=q�B���֜�+'����W�	?�?���)��R�k��1C�Kn��\�b0M��k��]r��_q?��I~<O�o��&3����*b+�/� ���C�T����� >[�qPU߳ltn���Nj�)�?ה����Ⱥ�Yfy�x���'囎�n�ij(�_>&q�S�qG>g�Z,Ѿ:W߫��UK�������d0�r� -^�CN|��:��O2J�W3�����h�7ȟC6&�xP?J���M+�3��{�ʤ�U����%j�0����#�98���%&8��B��Y�s
r��q���ܔ�3��p鹉6���;�j 9� ?��*��K�^S����L�~�푆p.ғ���@F��Z�������b��,���U�p�+��FV���_�cF�j-|��q�ĲD�ui��v���95�V�̌Z�J	Ӓ�V�x����wv4�tF��c*|���x�P�6q��G�����
�#����*�mZ��M��/��e�GG�C��}��h�mX*7�l�;��+���D���D~��$xK���ٝ������'v��\2@[obi��-�M����
�ӭT~��>#�3Iz��h�9s��Z!QCDU靶�]o���I��uj�Y�~O��(<��ʎ#V�cqVO���֜���P�uuvъ�z��CI�-; 0v�*��W�_ۚ���_�Z3L�l���Ir�2�ġ�"�;V����P�	��&�qH�.�o+�߅��(i*v���~5���e�#qhz`���|��*�=�5��Z�����]<ʹ��]�l�����z��[��mlUϹ���ѽ[:sS|_g��]f�_��]ˉ i{�uP�������4v)e��jQpǀ7�f�D�l��֧����"��@���J���do����Y_���p�S����3ݷsb	�P�E��7��ف��˒��%嚀���G�~6z+TB79�����#֋�t��eo�.�)��2�A�<W�Wl��p<w���҃����T���s}�����t��W�18�N��eE증
s�,��Qj3U����
�3Ϭ��.�4/u�D�7߻�Q�C5��� s�8ob_���\�)t@գ�p�!����n��'-2Ǻ1ߩ�s(��Á�J#�Es����Y}�y7l�_����b�u�Ѹ��-2u�����!�HD
"�)/�7�U͉,$�Z�y�>t>,o���Ly��;�!y�EE���>�wJs%�Y����g����]�������s�FE�*wS8a�	ij?��l�����}��d�lLΠ71�/�������9}y0������.GW*jH��ol�k�?�t�It��֨��v�P+'�L
�ޘ��婯
���F����r]�^͢ﭳ,3���I��
9p2�����sE��w�nI�j`�i��-v��bDI���May�td���a�m�������t`�����-;)`�8�K��pq B�Yg"d���T8l:��+o�6���������S��w�����������N�-iMrJ1��̮1�dϠ*�����p�f�����Y�T$��:p���*]���^��=����O�w���{V�R0�r��	�Q��������/���$���R�f�W�	?<��1x��֟dQ�@S�E"<Ry�1�@3�����)�z.�a4ݪ�2�a9v��<[�J8���(�O..[�dN�s���z�]Gꑖ�֛���ώ���^0�P��U��*?P��;1I!d�J� ��>����"�%c��k�r����ЩcV!2A])���y㞟tB6��v�VTre�a��b��%r.��Z[&��Iv�T����'1w^]��a$�kv���#�U7��!%B�뷠
�ǀ�O�ݸ� Ȭ
��Ns/��LqMӋM�\�v�h�H��o�9���ҕ�
0E�pW��tm�i>��Y�_���ga.��^A��8���j}t�̫�uR�cXy�s�$D�z�J�/�y_[7����~��Ĵ���5.�x����xȊ.1f谡B���Ў7+U�*��mr$��%��W�L��(��dB�`ka���a��un�Md���ؚ��Ć�8J�N�{�X��{�3�(,#�E��z�'�"K{���&ͦ�%��&s�!����-2��L���Y��٠���Gg�
Y�i�ҥCef��2�/y=�lx\��N.��x��h��z�7�ZkJX�i��Z�Y+���W#��s�wH�����i������@������!������܉MeFڑ���9���a��G�Z1� �:l}%�~��fH /������Z��ܷ�F@@�(f��<_�+�u���7R�w`6�����#c��MD��29.W��:L��إ��
xU�k
������J��L-[е�i�������B�%��
��H��I���@����t���b����A\c=z���sRp���C/Ƿ�j�]n�W���LH�T�CA�D��"&�����~@�U0�5��3k�o�t��͒뼀 O��	���Ԗ���.�����t����Q1Vg�>:��ih� ֗�kUҿ�}_��Q�����#��L��u4pLjΤ�g����$��%Sy���ݔ�|10�����n�lQ"G��+bZ�����9(�D��5�&r�a6���$%%O�KT����oŻ�O�||bx�vf�O	��F�1��0�����:"_R�j:z+ $.o��+y�_��nk$m��ݟ�����W��(�2idh@J�����1"u3zT�nI��d��ȓ�o��eݞCqL I��!m���#�=D��Kp��J=$���XT�(H.�c0�ڴvh^a�b��^�tb����ǘ�0��}ͼ�bP���e�r�Ws��;��Q'R��\7��cf����9�}�}���Օ���K�4�D�jǯ��+N�^x�|]�tqA������5��\��s��gp>6�!��k��D�R�>ؽ�3s�h��,	���� �;����[�+(V*%-�M���U3[`83|�9M���z��gj:����Z�K���-;qI�K]7ﰟ����-���:w~�@&�BL�cl�aB���SD��=���3�Ƈ�B���MJ���B-��?�9zuᏅ��7��f���CA�3Aܾ��+���Z\�'&&��"B�Y�0�A��p��Sˏ'x�����\[�����ã-���w�Oi���J�Q�o��2���C��,�w������*'F��&���M���J�3^8ŏ���+�@j���������Vږ�p�H���	C�1N�܋p,!��}J׺#��GF �dvae{�F_T�l�l\��mESU5z�
�/c2������mt�{_-	mƮ1�|p����#�)�H��w_�<+5Y�I��!� z����]P2ײ��z�`��f��ׅ�A�������
"��t'���s��������Z�iU(1���t��Z`��?G��jG���$rbd�hv0��B���M��R�{�R.��~×��ǳ�$���0!�6ܤ!���Ur���{!�ѓݴ�Ⅼ�Y�Jr=�WR�D"���! 7�I A��7\I�-�\$��3�&���ek�a����s��n`V����Q�}d�S$'*syQ	7b|�r��1����[W�^���Ȟ�/��sZ�����ڱ?��t��!���1h�s���]D�嚎Es�n��{���#�ҝ?���k��)_Ū�����ˣ�o ��X�W���� �T��ʨ;z�gۯdY����p|���#� ��v�*�,M���Q��g�OZW0���9m6KJn��ҧ2_� n:X�C~��o?!h<Hz���ƭ�
fD��L��g ��pp$9������@iTV����Rq�@�
��>�o�ay ��(c	��:�;v"k�w�|�پIp_Y�څ���C�-7�u}|9�oL�FL�����X6 B�:�I��BB�m
B(�Y��f�[����gv��u{��p��#��J`l�δWfg�bCl����=P�̋�����݂�0L%/X;! @��x�W����e��=n��[����v1�V���N�X�~{'CQޗs�h8	[��M�@��/�m@�u����xd�v��k��ZZ2���V;�9���i�)�X�"�yf�c�̚�cuj-u[(O�5��v�d���W@�it�����AyU
�-�N����	���ܾ�z26;y#y�g��D;�g�*�u�+Zūx���+)����Z����{)�Sz���_	cA��Y���O����x��F�=��-*9�MP10�c����x	�S�'�g���p%;� �ܫ�<�g�U�f:�1�o�"别=���É������.F4X�z�p��p��j"4�>T����!�9VFƔ�+ViЭ���HSH�DZF��&ޖ����wyE-�d	I������t=K��n�N?帴9g�OU�OĒ�wh?^h+ �Co:�]�F��t���
ʐtJƗ+%��4�*����&�M~j�0�ȷ}�D��N�fpb�$Ϛ��z4Ȫ�Ymv�(z�E��w$�h�[;.�J�$b�_O��*8���Os-��\!`2v��k9K`(�H���4��vvwF��!�����μ	() df�F��iT�4S��5�c)�W�h�"{L�x�y��ў��o( i�q���C�y�Ѓ�M�O���AD$oz�$t�W32��br����U]�jh|kq��rp��z�u�0��k�>V*#9��)�Q	�%3�G�ΰ�n�FidKճv@���iI�v7�I��IC�}���j���?<���Ǟ����Yk K��ge��J-	8�XXo�#������E>�����A��3����!��-K�R�/Y�x$h�Un ��RXH��d�.�v�v�E�$�i�je%�*�3{q�c;� j�R�%&l�}y�8V�ڠ�������ń��Y'f>f��|��+�S��~1�B:��^�(��������<��Hb��:��5�	�y��b�8C�q}�p㎷Tlƽg�G]��$n*}o���Ԫ�%��
�ɖ���y����#oGΚHM֩G����$T��W��x�DP"�~��Sh�c�eu�?�sx�f����  8�rNr�4���7o�\���z�%	�*z���G��)�L��4���Pcͮ�n��O�)���x��]�ELAa�_�\�������w�  |Tȭ�C���Hw�#��Uy2I#���Μ������Tw0���@��f'i��*��I��"��\�񳼚H@�f���F2��.�o{�	_2���ŵo�Sz�\8
.�2���\j(��U^�1_���������,�MR�y�O��s�r��V�c���ϟ�bX�s9�Ϳ����D��c��oX�L���b'?��8fl��!!l�X�a���s���<��O���=L�e��Ʃd����s��w���MR���>��3��/����ǉ��(���gF�Rֱ{�_)o*�����D���V'( r�q��~�,�� �`�m�w�̉ ��zٰK;�Ws�;������d�� �Uw]7���	 TyWU�ۏ# ���� ^}!�����4BK���T��
E;��9�&M�psE�>yLIq��R�uz�2��;@��l.;��✰4�s<bڋ�
���|��)�Nі�4�#R�PӚ����܁�9����f�u��$�d {W��_�Ϲj�jI���2�������\�C��Y���C_դo�Q���q�[�n��gYz�4�*x�0�ڐ��~H��:�΃���"E<$,�e�([�<���)(L��P���ɬ� zA�L�;U6�J-��z7'�Y��k�	�-%/k�K��q������[n�Z�G��s�F��Y,�g	�Q�~�YbL�A񷮂s���[�:{r��-��ir�gh��@����/�Dh*��L�~'R6f$?`1c�)�I��.or�8�y�^(�Xy[��)zبT����eT�:�3�\�A�y�/����b6@��-a2���s��N���R�g���ۮ�'� �J�H�*�U�X��m ��jX�c�l?~b3�}9i=A�8>�cd"Բ}̦����Zt��D������=%���AQHQ�Ԙo��;��U���Q��5y��z�-	�UҀ3�M���2�*r[M��9�y��N�bF��zc6;����Mn�oT�a�h]�<�Z�S��b%�Ӽq0����ƨ��ƅX�/	M粫;�z��H�4�����O".~�Zy�SE�^|y\�?!4��e�ɳ����p�EJ��ϻ�>_�����;K�!$�-��2�n��2�{S�i���S�Hy�i��2��V�j-3 ��K&��}�X�!¯�dVҒ=�:�>�M;`ҵk�MÎ�\�2oķ��<��Y%��]�/�S�/ď��lR���Ȥ|��WN�s��Ԁ���BD�k�ٳ���X�!��� !̏O�v-�N�7n�ٟ�RZV�H�aS���3�J&]=-�S�1�NlMS��!���饈���	'a��FaӃO�-����;���0 ��a��?װTǍ« .�uQՏߝ�_OQ	�Ԥ�+�D��*8��s,q��)�����ew�[�H�<Oy�%N3�I���4�hUH���7���7S���"!��dt��w|_12�����~�:?i&�x��d�5.R��b�D̆��kS�H�&��*��B�@��I�|s%��ĕ��|�Q���7�ֵ!���YA�~���)��l3���eg�E�N�ŉB�G���m|���{�s~�F���x��ɨT��m�<�iZ"�ct�>쳰�8����f��h<Ď55P���������׳e�L4�W�{�IJ�Q7�K�q��/D8���Ia�q��'c}�&���	/��͋��!0�C|s'�v�\����^ޕ�T����pz��/H7 ~�ɽFf�ZJ�:���vMK��m�,Q7S$�N%x��T0�W{��R�՝Zj����q�
3Z��cեL�O��Պ��I��y�)J����z�1JB���Ʌ�Hjv#A'D��wLn��2�1���o�Ui]'�ҊϿ4��M؄r�!����b=���n���I���%B���O-=kG�R ��t�Ѻ�������.(��Ou�bT�X���cGMz�m�����.�s�ޫ@^�\+ayrz�X�WI~׊�'Q._X����I$��b�yݗ0g�u=���T���b @�sJ7)����L��B!|��s*L�0վ)y�9����e{�u8q��[��l���ig]�;�ofwn��;���he�8ˍ�w�u�LZau�tjC�ce*F��v*?~I�k$�M?�����ֺ����Ka�B��r��N�rdc x�՛��~��le�~���!��&RK��mmO�F������w2I�0[�����7�Gn�y��W��d���f�ۗ�ע���S��8E�c�V���)��9T��ƴ���&�y@ZJ�d�ͥ�l��Sq����D6�#��� �e�<���HE[��)���,��Rw���ױ�Ͽ����|�����38����jSL7aX�bg�a���C+������-����t�4��~>l+~+�T8�5�[M|c�u~����{,'�JX��-��ӧv��હY��^��R�kߜ�Z��IW�s�.Q0~۱�6Se4�j��H�a�m��8���hں�RIg��5�O(+���(���\8"
�b����@�����2mb��_���%#�/&~R��1�E�}�:��}P���N����Z�T:nQwH;�����Hӹ�e>�P�~`YF�4p��thT��nm���!t�����j<���r��Q���{��g;����'�%��Y��&��e�1
����0q�ش�@p���	#G�C�1N��Z���{F.�E��L��}���i�Uv!wt�X̢�c7@=�u�9+�|ĭ����]�S��4S�J��s��<���ꣀ	�0�,Ŷ��7M�I���}�8�$�{K"�/�;��E ~c�3*����5N�QZ�J�d��2C����?�lm�}���!֙y�Ȗ�K�.Ёr̞VĈ���Q�
x[G!�� BQ�9�^���W:���X�d��̡��/��_ONÅ�S�u��DuW��>�nQ����v���ɾa�o����� ���!�m.d]�C��q��ek��t��NE	x��*@��AĶ�c�+Tә�$Ր����n���Mͣ���C�o�h�#����� �@�;�'�h�aY�����b�Z�j�5�WJX!�3�`��B��.Ar���m �:(�-�� �B*�IƄKH�赏y Tr�Wc(7!�4��o�r�}��^Y|T?�[�'Mh�!�[,�1^���F�G<EIc�A��J���� �{C,~���	$�DR��?UZku�/��'`N��ʓM,�Cq������V=�d��J J�����(�Rhw���5���_��)��
2�/�����]��\=����Bӏ�i���ۚW-��?V|wbf_Ơ���J4� ��>q]���$��������pA��O۟���O{���/���O�u��IX���Q1cY>���8��G��^�Lނ��⎪�P]D��m�2d6+�h���6v^�E�rV��:� �j<Q�"?*6�m	�祬����ԅeb=�� �ڲ'9ä�Ȼ�fx
])cXR��֦|�-j��/���z��:���rrL0G	�F���
�Ӫ��$w.����ȂJ�UAPV�w�:����}~�7�SҜZԞ1sD�tQ�4;'���[��a�9A�l@,���?	���;�lJ+�YX�%���C�\(7{�G���и�޽�L�ȌS�	� [<)�lS�|�c�����l�%}��y�߷,t��9P�O��̶@�tO�ɨ'5A���+wo��\[���*��+���4<�s�9:��)=�1���XZ�O��'Tc{��GD<�j�h��E�(>䛵V!��+�T��[:Rw�]'�W0�^��L�k:,e!Ņo�>+4Z��΃���F5��mg,�h����Ye���?� ~��+��`�zL
��K��.����Ⓡ�$vv>x!��O6��Tg���YR��M�O$4}�D��=�d�$ �_��*	�'3�H�􅽇 u���]ԄK��5�f��A��O�ſּ��U�P�	�zUF�,/�vCbid��9�W#lF�:��d���C3�<�/�lT�mE��>�XӃЯ1��^�{fT���fIJ� �?��4�x
%,�:��"���u����ܗ}���Vh6-��A�oz���� ��C�ay�p�<��G��� 0k�w\����]ph�_BX$Uu�����#��+�t6�jp�GT���V�,�ؒ���Q���A'W ~O�۲;��� q�4�2�n�[�9�ı6�"39%5!�_*E`�n�; *&�&9�A+5R&�c�I}�@[��*��%�������zw�_���>���aN�A��"�����6��?���5��h���w\��gBU����H���	�L&�h��o�.=6�NA4'=�~.�g�N�bډ
�C,�*����,l��`��WsP����*nu/���i�#�˔ P��D�1ĸ�ӕqn�W����*��@��׋R�����p��ۦ�n㮪���&�.�8�cu�)�_����A�ҋ�W�$�=�5.�QD�T��,�v�K��#��q ּ��[�+`*"���N�����kB���/w$m� ��B�qɣr��}^�F���]H�#�=ov/�Z�`[��I��1���bO��Y{���+����3�&���Y?�_��.pzK�Rіd��C;Q�}��g��o��»�&�x�����mBan�t��2�tSKWDQo�
j���'���W�#��Bޝ ��O��9�R��U�'��\������yn��oźJ�c_�@�Y�5�^q�.����4�S/mF���4}����}*�S�=�A�!�8�OM�*�C���n(��k @��=��I �߱]<��$Z%F�J�D���?�]I+���(���&1��I�?�����x��P�}=���"�jX�`�A=��Ή�@��Mg���ڳ�YV�8�r0��ß@�c
�A��m�:�'�5�@?-� Xցzm�LS4N<���Ox�`E�q�����("�qpC�#��<�2���ʢ��<��	��?M�ˉx`(�j��|u�,��\�:�20lL�R��P�C::p�i�@�� }���T��F@����!��/v:M���u茤��譏�E��`�dN|��nTN;�����}��俄�MbJ#�����S����W��hu^���`W-:��G��ˉ'M�;C�
�)�a���]�!�w(�V��bRr��B
��C{��ؿ5��t���s�>�g ߋF=�5���dƅ�zqr���u�n��
�f����_�D��'-�	������Y&3?�?魻R�� �]�v������&8���
�@Ƨ�|��c2k���uM�E��2�M�G��'�3�wq�B��ም�UG�� �ᓜ���-Cރ0Y��;�����a��r|Q�ʒ ǯ��@��� ̞sK��T5��=6~�4�&a��Av���}0�.���Tө=oᕥ�pe�t@L)��{�������ck:�!f^��D�rN
�Zdg�TϥThI�����\�S�m�N�/�&'��n�O�0�u�V��j����nmO�sV����?��]��Ir���V*�x�֋�w��x{��͜|�t4s<����p��~+y{>��xDG	��T(rI��H]�?����<^�t~Ay����::�!��4�Mn����3z�6O�=��f�*J�B;��T�PI��4�d�����.*����~�S�>M���b��+�`~�e�7p!S�˯�bTx��t8��`c�B,b쭍�
�U�F���u?O#<�ZH^��X���:F��o��	���|�kto�ي�@�D5^+D}_\�i�wj�ӀC\]�l�קm1��}c^�Pi^TN�[z�q��ؿ(�B%4l`v����ڼe�YN1�ƱeľO{&ȩ4Y�K""����l��y<�<P �U��e���	Z_��LH�L?����TG�)B�#su�{u���+x�����$ثap�߲���Z��"P;{.���̟[�(�s�֯��P]��E�>�\ġ�T�FԚ ��i��D	����G��dc&��N�����oWU��4:�~\�ȑ���'+��_�C�p]T�Ʈ�KX��"#\�Z����3Ω���3m��(�G?RAyU��ٽ���'��\V��;�O� �o��m�}1d{.
�+u{y��ƥ���9o�6�� oq۞�8p�o��pY�Œ���J�ˀt��3�ٿ���uR@�����_02�ʋ2���(�+^z~'-��`"R�\ӧ="��ibl�'�V3�G�E����ݠ+�������IŜ���@S���c�J�@�-9[��"�1܉g�;�J��/E �؇U�����X܊$�p�^i�:��Y�s�^��8�Z?
~:���ii�	ƭ0�n�_;P��_]������q�t(D�����_��� ��J�%���'�A��9��g�be�1��e�R�%�r�Џ���=<J>M�2�Y��?<�bjY�":������K��(8Ҝp��լ-�yw��I���סvCo����jn@Wq��x�\�[�H���dj�c���&�<���V�`I"�w*\_#J��3;�yqN��`a�a΄	�*��3K�Q^���,M����-F��O�ST+���GQΚ*�e�q�����k�R�,t���Z�n�Ϛ[�d$E�Q��Gr&�ʥt\@��uM������Y����^�T�a;t+�vh�,%oC��ap#����d�����[�_�=삟�e���ç!kdJ?[���� 	/È��U������=���*�|�
� =�F���� a�~��/2�DX�.��B��`��$Np[S@\�g�)�Z�N)���V�(Kԓ�	BQX���e�&: dQ:Ș�7�Ix�����>I�9�T	\=��x��t��̆��P���Yt��8� ���b�
�!��?}HH�ʠcGG�?�wlF�ۨ�uxg��bU��,���}���T�����p&:�z��r���E, �.)r�N���h����}ň��Ep���������پ�i�*�b�s.:X��"�	T�u�x3�
��4����f�U��,p��g!��Ӆ���{�rg�; ɩvuJ��FiZQsYu>"Q�u(�ќ(�?��4)b�E
�����].�U/����18m�C�"�j��]
ri%&�ٯ?Ț�^����*�V�:��H�R��+��i0=��j����x�d��|�ݲ���_LɓD%N�����*"��
G2ˬ#q����߾��Hd6�	{<�s��\Q��
U�k�b�ߎU���c��M�χ�Bl����~�B*�<�ZK-��0�E%ڛ�N���X/.�� ��J�ڂ6�*~�@���.��!ͯ�=p�~Dn���t�@A
���1_-�G�%�x69{^�E����4�-�n�y)�rzAj�E:�m�.��||t9!�>�ܦ�Y�멚�f�b6�ާk6�/��������h��"Ӥ!?N��p�sPC�L6켾C��e/�=SM!<8�i��x�3
�f3K �,`S?�D)�����t�G=:��ˈ,��M��@�¨��#��U����\s=j���-q�e�Pq��]���q�o8��hPS@��!�>.h�MԤC�$E!k��J%��+v#�0|�W��	�j���%��u" �#��A	�ɠ,�{�8�,w+�<P�Q�y?�>�Ct;J�A��ޏ���C�R���3A(>Z�+:5��B嗯�����3b�t�No�ۿ\R,!�f+�2�S�C�} �qZ�������̃��WSc��������n�}d�6�3\��J�GP���w��YH�^TC�[��jW�Q�9�l�<��F�����svp���<SzK�xs}m�����$w�o�����~�n�>��MZ/qdӏX�Ɩا�������uۏE�w�V��r�ҌmZ�:Z���6�Y���C`^a���~I�,��IGF� z��\�]&(�vRtT.@x#B�%'&����7a�8�8��-JFÍ x,�	^|��^��#S�om��wd��	���2FEo�C؅Cw+��p)]
C�Ä��a%w1<��^�d�e���p�vBn��4o��� �8N�	�($�{��ٰ��
Q��Ȉ�=�H������ޗ+�닪"`2P.l�
�+��+T���D�-�)�D�E�
��ئ�_jο�gN�
�
r��R��Rn1#D��4I��g�h�����	�.�`9Jq�]�! ]�$-<9����͟N��b¾�BB#U=:w��|�F8���ʏ_�a�`�e��m��S	gu�]$tV䶧�J����|d4�q=e+� -����|�3��\���&��Bt��tXNم!�Ýe������
�)�M?��34g+�4�ȌP��E:��-6�$i���OOG��X�����ڼ��=gCi!D��c{g��I+�30�ag�8p����d˝{���^��P�����ِ<X�X�fУ�@}Q߿���h`�r	��Y����QX��l��}��HB6*{e"�U��>���ˆ�Ӎ0��) zZ'F�T�ĥ }<{�kg^v��ֵJ�k����� �����`���v�Ax��\�FJ�%���RJ{V	�i��g��� c���k����W0
^F��a7��μ������]�>�����ә���&i�,����l2���	�Csډ�:��v2��8�s*�L8�РVp�`��g��yTKv"�`��	�]�u�.�ܙ�(�t]><½�_8$�:z.0�)C�� X����K�܂� 1��]�A'=��nvGqp^��ZP6�7�B$➩�_E؞�����ӌ�GPٮ!��Q��Ds|^q�'�iKZLF���3g�yٞs��䙅��?['#��-=�N�����޾"[�O����䎽׍0����B���@��o�DR�j��>��F�{}�=[��Q�����fC^�(�c��Y<u�=��OU�%*|D^�XVd4s� ���ؠbqd�^����U��]���I{d9��{�s�烪�����UB$����ɔ�EƷ;��}�������sR���P��&�-�2��!���~l@��Ec���=cI�0`������J�e��\�31��Յ]�ى���� 5��B#��+�K~���U�S��`�9�#��kk�%���>PPHI0�<7o|5t�[���8m��G_��K0.˨�[�U�G�=8
1������a^%����4W ~�R���&��i����/:)�\� =�A���l�<�0��l� �_83����g=��/A�m�(�F�#���)Am9Ú# �g�R	�-#,����>(�Gpv��Hŧ^�=h�A>�H�5�K~�EAX�Y~E�1'�%���ښ
�S)���A��
~$�������r�-y4:�^ 7)]�U��a�4g��b��?BD�|�!�#.�G��UŬ�ZS��[ޫ��ʠ���3<݂7q-q\��u�1�?����-l5�o�wq�		�W�.f\8~�wl&� k0	 �(?缛 T�E�{�����F�E_R��uA��2�D&�ޣh���'��=v;[�BH+c���� ��QƖ�y�����7�<N��*�~Y P������S���
7�'�������s�D�Z��;{���������y� h�)PF�Ѭ��z�b�xtH��2���I��D)�wکf��'��o�������<�]���&�W�hr܌l4�ohdM�VίV\K�ΐn���LwY�j�����VL�B*m:���C��R� 1�V��7�٧�����=*�t,�9��t����g��$�a��q�LH�#5�Y#��a�)�Y�>j�\�J{�~��4<����cە��!FM�&�zD��2;)�ܛ���ū+�ٚر���m�Fkﮋ����j��'�&�Piiߍ��U��V�]`gD!�oAh�)i^j�7�Ne���͑tȺEQ��X@ �vM
���%���G�Aބq\�z�\��d������2�a-jry�wb����}��}v.aZe]�%(��J*yv��06Bj�~[��{Z�PX��T�}�VsS���/����G32E�����VrGCᖨI�SV&ýi��YQs�������	!va�n��q; �[�I�]Tkg)Y��%��+Il���[L�"W+�>�,�g&^5o`��9@�O�~��>nY����m`a{	xgُ�CE����ZŽ8�I�	���A�Y΃�ś�̚�}��i��H����f�V���\�b�ӎ�;=�*ʗ>R��{����p�����A4�B���!T�WF�p�ws�gzC<V=�a�:�B��ߑ�'2�f����*��B�Oq����,U�8��	j6��좷}�?i�&5Gy��P4g�k�i:�]��t�#cN�Yi���{�� .*�4�C��vK� �C[��w��-6�P�}�1�P��=���#	�����
*f�Cȋ���O��N�J���Ȭ���ᖡ{�XX�d��ͬ�z�Ke><�}D��r�Z:0�ĥ��8��7�0�޹�+�𴛮]��3ɺ���E�s��f0��ONk;r��"�;��9�d^�����?��Z��A,��������V@��(�&0mϕC����w��Sww3�����2�� ?�ʁT�|Y��!�7�U*����j�@�NL���t�)��k����{�<��5h� dt�`<�����T�pQ�z�Q%B�-��ش�������n�"Ɠq%�R1�MLB���w�aa��1��;��@z�����eg\��XH2��rh)g�yu���N	���g�d'��T8yJ��a�5�6`���0��m��ڋ����>��U	A�����ڏ�j#�#Qџ�+/�lz�V&���$Hd���??�ݪ�1\�SV{3��׷{(�����zs���}��>]+i�����3����)I�?&�h�J˒���	K��x	۸�O���C��K�L�� ���.���[t�����b�c�h$]�����j�3ȫ�e�g w�=����zgx�[�"�l[~�f��'ɼ�`��=�s�,8��ahra���=fH,�#I���ĔJj��«u|<�W����#��k�4i\J��$E�?�yA�LkkyO�ׂbdԨ^Xr��QrY���M�Y���e�'Sdbu�f�q(&�T)�(���P;�������&��TX��W<!��W���@��C�H�#[�w�^�+Ha��}�(�н��~����w����sӹ��%v�'�bF	y |M�3+*)P���P�̏���87k��w����,��&��MN�qĸ���:]��+g.`�/WĴ�&����k�-��f�"����o�x������H�R��|➄a�k|�+bډ�M3�ʰ�ҟ�j*ޝtن��09MV�W��Jd��FIJ&;�p���x���G;F�T6�}D>f8UN2*k�����}Pƀ}Q��>zt���D�u����D��P��lw��;�
�L�kgê�LJ3E�]�G=��S���,��:p$ɶ�'�@'#�}-��--RbŊx�'~@0Q�� =�U����`엷�{����} �4L�%�s�len��.+�E�����JTo��o�R��l�CV�Ӥ�[���rq��๪Kڙ�}���u� ��2�+�<�E�<:W��/0<y�%��))va���9</�pP�t����,)4#�D򍐗4��Cr�K��
51���?Ix�EV�x=�t�04gbo (^�J����>�Oa��N<O'����������R'xXܑ��Hs:?��/��i�֩����:MѰ�O߫��D�pl�]f!Itq�Ȍ3!Z����{q"⌟�K�����l��6)��"}R<nWR#���z�5,�\X�T�8p�ɘ�+ϴ�2sz�eB��gn���{c$$	B��[w���ޕ�wH��9��S��H/c�f��#�[��Q 35Q�!Z�G���2A����e��|?�%�	�S+s\]B|�����S�K\.�Xp�(����e��y�
�d�)���M��:KV���!��ƶ)��CI=�G��{�='cF�.����$�k��Hw��F�A}����+����|����%���/����>S0x�����=�Ї�
Tr��L����h	����s���,Y�j1@��d����������1M!�>������ 
�Ҭr�����K��@�_�$��}���4���}'�,�i�%���]:�aƝ�-�� �.��3�Ju��Ss�=�he�N�\�k޲�KX��B;��,�d�`��:�P���1c��=���:�FU�����{�>�E�?2V���]�~�	Q3St�T�P��$��^ń!fx).�v5-E�\RǍ
�`�eq��)DC����R��g	�Ƞ/+��.�Q	�g0��H{�R$�Գ��C�4��$ ��_����~�3#����_�1��q'P�	�� �������Yb�->��{=� �z��xe�례k�Ԅ׈V�6E�k:H*�ejv�I��3:��qL[�A�	@(`�l��т����j�)Rc_�J��W�{�^ۓB>I�q�`/�[��
�f���D��$��vu? �9��c�SOF�:���#ԅk������M<ZW��� ��{]�4���b��&���c'*I��D�Cʙ��<��re����}�GԴRn�;*�� � j�Â�U��ЁH���W�M����9C�9�""BW]��ds
I�NH2Jw	�)bשR�K��	9�!f�@R��Tj��H�hj �����EО9��~����-׷8Q����=��ʻ��ŝ.w��/�=�;�~����*�W�*Y�ϳ}��dX��"DQ�e6���f��L�%Й����=|��e�YW�.�S[����r�����dտw�}�r�J�%�Nc�i!�����Cu::�1�涧�)W?�����1��;��]�d�g��~Wqu������v�0E����ݡ�i�z؂ `Nn�eپ�}8�5�����F+��ȵ:~ʛR�Vq&�)�F�=�K5��eq�t04Q�⤎AK����9�]4H��J��2�}@SX���&t�=�*�[ ^�.�=3�,2#M�.Ѯ"�%���emsn��� �	?�|���2���y_���)Ƽ������R�4�r��E�$�b�of�3*Q�&�g�������2R�<��'�����:�w�@&`�c�4��̱
��!S%hPz��'�;�K�o�+6�}>T�=!HQ{�d��N�`�L�,�$���N�9���n��hr#�l��]�Bud�0��R��_��� �II׻V�%�	V�(�~4����0e�0����W�k�f�_�	Pŀ���̳9�Κ,����7��UIS��ӱl��qW�[�wxe���փ�%#�B*XAkV�9J($� �������g�u��n?�͚��UD<�{�<��_`>t�X��e�kt��"��#j3@�.���@de���%�hRo��D�6�t5�h�{y�vר�0@Yq7��RE����X�W(ϖ	��X{�k���9kF�w��޴��_�z���ix2����d?^�JmO�P��2�"d�S���v�Ľ	j�D\�&c��i�0[y]�v��mk�U����t���o�ퟪ�����8�����;~�賀4շ��!�K��PS{����+����G-C@�����9�%�x�ZO�DG� ��<�5�/�|����D��ęVϽ�u�,b��������l���B=��HA5ל��7\��'�-�W&z���;Z5Y:r�D��1��<�t�+d(-�ꈧ�[�����X(E�����<�F�����p{�D�LQB�kg�Z��7Z^0p����'��I��jk^��@�J������v�4Qe�2~Y�HX�ר�F�e�#B���U��c���K�X�M���2���e�,'�!+r�8Y*���!!dVL�g�o�aw\���(R�΅EU�wVH1(�Hz����یD�>]�|aix/�P�D�<-�X�m���|�a�}��-��ԗrh�\�:���_��r��͸�g�1n
J����l ��M}�-����X� ��֩bC����a�K��q��JȦkk�*�_���@KeNV��]��AJ-�϶��W�kS[�I*�H,��М�i����|�����`p�x�6$�0U,�
��
�m��G�Y���y�n �8wR+r.,e9GO��q&��#U1-�W����D��mͶ!-q%3�2�fQ�j���[k(.���2����� @��bf��y�=�T׍I�-6�2ԩ���9�#I����<�Th-6j�W�����IB+~K�yV��U��%� �x � z�
|��-ἀ&E�SY���S�W�$��Kr�j��g�~�3L��g{��Z$=�3W��������4,�FsC��nP�S��P�-]epg��g���ү�~	C�s�]�5֎�ku3�5����|l)*S2="Na}T��#��ɣ9���.M�"�^A�:�>�T:�йy��8��)�#�}{�vt/Px�5'�=���p�� ᴯӈ��0�DC<?��0mjv�1�9V"+�#�à�����9s��+����UUr��ʢ�q�|��QuP�\�@7ZH%P0C�>�U�:?����������1��
�L�}��]t��ܖ��o�A�6	�S`7��.%��#C\�E:��Y��n�B'I�/5h������M!ʅ8���e 3��]�s��ɨ��ٗ��?_�h`)�"~n�q���Q�է�'��w	��z��a�6��5��5;N?mv�O��.!���u�?��'ȩ�f����T�*L��0*��[���hAdu0{>{�������c+�����i{����ľ��ּ�^M�x�� 1*�J"���߅�X��}]� _M��ܿ	��N�O؇�˸��cU�\P����iR-��J��<cNé"�>�4I�G�����S��RM���C���}zTߧe){aY3h�Q�t1M��
U毰�h�/���ڊF��,��-W�pa|��(�d_���+O�,'�_�l�?����$����y�h����խ���ihB����;�'G��`�@I�<ؓ��j��%~}?[��$bŞ9�����!��95V8���+O�+�&��V�%����w���!�с�@����C��Ѓ>O1�b�"0�F餤�$��O|,�iW1���^3����C�i�Ͳ��x[�9�����5�~<�~&N��F[�j�3�q����^���D V]�_x��~��֗:w��_�^�'�Z�`u��H��a8���XvQ���01D�B�\ԗ����<'��'A�}GlD��¢TY�N�'��r�vVغ_���(�X�=��>i�S�0���}�u�
�uȿ��|I6�q|�)��M��L�Fܡ����yԞ���ؚ{���vmm�W�H-�5x�=��J/���fb�
�*�����{&T������X�Jt�Ma�`rzϗUbxмY�U�rhҰM�<d*�Ջ�a��#��e\�ʀ�(�`��[�ĥ�Ѿ<��rc�V��
��q��۽=�N%���=4k�(_�{i\�gRd��m.�"��͝m�W�e`ᖖxs�qh�ץv�S8�TQ�q(���"' J��>����4��z0�H��'���>A��������᠔����� �+v�fvC�yZ�w?bMp9��>���@[̧r��\�v̨"l��po�Z��B�9x�K��2;:DMM�WV�t��.�w�	��P��=�6c\ܡf�v�*6�����I��.sÇ��?���4�5�C���4�!��e�R�ꯞU�avp�)�����n��c�JT�A4�%����9 XV���Y��.�Ft�+qPY|�:D����)ڢ����6E�k��.�TV���ԧҤ#s�TN	滘�$휼u!�J���w#�R?�m=ig�_Gc��t��ũcH4�����m�3q"�:6�-�ē�ڲ1�:�*phs	�G[�Β���F��X��侒LG�@���g��YK���dC� G��H�#�P��[J4�b<XW�j�g�M�pC�*��rG��eU,�WV���쪵�}Bn�qȓ9*�H����sCc���(G�^/��9g�֢�?C�p@!�n�`��\�U����*mdG��Eo�������h2�2G�W��yu3�0u ��=����`b.��o�Qdj7�i}���!/��f=̞i�g%����~�q�1��]��6��"������!���4�|`��Zq�6�����.��pV��-U���r���P��D��.��l'Q있2�<��g"���HW0>�K��?Cʪ��[�N3�^#��7Y�&Q;p��w�����Y����X���OKD)7��g^����=g����"*��m�OGE���y��-�@nP�9=�ڗQ*�W�����Ջ�@����-[�;���mb��&��m���-����:�'
g0���5p��;AI۶嬷�����%G0�c
7Q
�7C2�R����)u��7+�B�gi_:���m.�G	(�Z�L�O'q���j`^%Xȩ[���1�`I	wW�u�G��,w`�Qa�8�gۣH�B�{�/�w�.�(�U#�r�^/�b�����QQ���>Nl����Ѯ���F����b�Cx�"{�c��ڷw՗C%N�x�����P����2i�q]��*�ŷ0%sy�ѿRf��m?�t�
�� ̙�s�F&��@��TH��1�%��{�Y�[m���R�����$�
6N�^.�n�r�.�[�r	'R�i镔di��^4ǡ�T���G����I"�~�Ҟz��8���R�ǜ�g@%�(�[�����K��<���Gwe䭎�HR�63��L�9+����\>R	$ۭq��C&������t��FƩM�ic���k��L���o@�wu�tM\���ci��,�^�)�L�#9���[��뫒�?�LC�[΂-�SJ�)��ʆz.PФ5���������r��i��1�Hy?)˾ϰ�$��?*�/�)x;�a׋$��l-��[�}���q$-=�*iex3�c�zŬ��'��*�W���v�d���Eq�,.xOH��Z���zl�+ަ��[�p�c����}?8YCV$�J���=�s=3��*O�49�0�"3d��Ts?��<��[�5���Aj��NH�2]��UŮ��ؽ��^g�N��/�\��p�S]���:J_Ƒ�X��Q�7���"�Ƽ�{QR�QF�m��u�j��PP����k��숵q��[[��W��D!p-������^p׊�8a��Ѥ�D�K�-V�u��{�{Q���Ú6�߼5TU���b4$�Qރc�k�9���"�})D����G�&r����B�I�Ejm6J�2͟ȇ�}-v<sO)D�f(�O�5e������z^&f�2��tFQ6���n��*?H�Y��ԳHAE��s֠>XЛ[߃0���`��[��&�sYK�&�8�"��A�
��r�Ɩ�>�N1���dL�a�R.'�,�e�Ƌ��E��>�*o��������HaM͂ozFz��-e�����7ɷ�5v���i�M!2s���'��Gw�nWgH�
_������,_�_S���6���M��LF����ȹ�F����*�|���I��n���IǀͰ�������+�Tb�R��y1Dc	���A�B����"& ��&�ͭʚ�d-����;%�M/��W��}H�<+� 󁹅BcEkf�^���6�*H��l���g�e1O�����DҚ(��OQ b���~�Ճ�0���1w��~c�8�k�Xf�Zo��+)!�<EȋzTV��M���	�U΅�BbՁ�v�ه��kx��g[�H�J�����?�2}M����F,�޺x�v2���T7������R��?|3�w�E�0˜��aG;Y �J�Y
��-�
�2Ym +aZ�]���0bq�rn�Z_�]���h���gxS�S�p�#np��^h9.R6�}�C����M�":Ӫ�/P5N��Y/a�ߑb� ��#g�k$�|��v�ؽ���8U��魃���
�] ��/�0@&��b�,�\�?[Y�����J�
����h5P�]��G	� !�u��M$x���VIΩ�-��Eޜ�*@[����E<�;U������nc�LL: }�A�x��v� Z>�a��"��WC��[��o<9²�5�.Z� ��	WeO�� �_Z�{dv)#�䇄xC��v�GX�@�&�_~�O��`���P?0>�+6�}���0P�m�x������:��s�� �8���co��A�MR�zd��n�Q:Z��|g�����FG���89i�����È�H��<]�%��'�6p��*���iǳL�y*��2�R���z�1�Q�Wҡ�nU��mk�ۓ��<R�&�����ò��qN�2s�^C�b-��uC�X���l_5�)��QW�*��mЎ[���$�	ES��DM��~w��ƟE�&���[��jԯ�fN/P���ecD�>-��ո�v�w�R���Zd�X�K�'�*�$~'/�U65�a�mO����K��]}(��5{�tn^@��|xb�O��i����z���l���z��F�[&�w=�_&���0�f��6mM�u���2`��Mz��\�\Ջm@eJ��P��ˢųY���DODL�(h	>��պ���*wAF���4���˼��: �ng�}�/����O�0��Y�՝�Pt�W�b�����ʃ�T�ޕ�	Y�y72��{�B8i��[�g�^~H�%��z�mrw���AΕ���𜜩���/6�@e���I�$���������� j�;	�&�â2X&>Ĵ��V]�p
ʺ����
G���Æ�#%	|Y׼Uo ��{*��!R�%����� �	��%|�����hd	��#o����(�"_���3Xov<�𳺖�O�n襷s/�[`{���1�=	�#a��s�ֳ~��d���1�*gY�>�+r[��e� '�@��)T���g��<����WϢ�.>xڪ,�Oz���;�{��m&��(���'
��F��74������l�<��c��ە��'�B���7�;qB�왞Id�g7�F=~�C�n�6ِ��A�#C�n��;I�`$~��!m[����¹�N���Ȼ�{�� c���b��5�����Nk�&�Q�O�et��O����Z@�f��1��I��\��;j��Ap`^<���S\��H�*UṴo����2�aA]��g�Cǳ���"P�^�K,��H��x{Y��7}:�&����hP\R�Ζpj[,>'t�a+n�h���1�Y�酖���[?@�s]��u!Sf�#u�AA��&)�^�y�\�մ}㭚�V@p�c���".�n򆥋��:&��._���R/&P��=7�K�e��SxI]5N0P�d��NѺ��AH��Vؖ�m���&�L�6S�4�%���μ�*�zH3����*ODp� K(���Tf���X���.P)�壥��BA��)��������%�sk�e�7�sRBwa {Q�v�c7���fq�Cu�X��DR���8q�:�Ro��u��	%��F��o�&�#_0%ߢ�B�QG�X��Q[��9������I&_E	�ƫ�w5`r�@�s\C�����l��ְ���1�ŜN�����e ��>]�v
k����ų��W��J��&e�N�KN�5[����*H8�^6�ô:ݭm�V���J9��k�_2��pú�E�����>1�!.O%�!�֡/:B &�8u���?�	����Z֋7 &�>.m����r��Y��� ��KI%�j��V7M��M�zd�MCm*��1e��'+m���Q:�@�zq��<����3}Y�ڌ+`!!��y�A�p-f� �ǝ �����ks�4P���<,�g�Fy�˗��%~��|hwJ��5�ݐ�}#�
b��[\��+�
�BE���\%�"\ݱ���I�}��G��/W���_p�>t��l>A}hI�ĸ}8t(�w�x�Q�Z�+�}�봧`V���t> !`��|͝ u�;�� �aƘ�.�Y��$�