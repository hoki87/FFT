��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�#&��#�<�������N�4@S�y���zM�|=�ٜ�K㪼"���p�A7W�JIvw߅� �of��Tg}W�t��8�ɺ4َ*��iYJ��$-��m%w'k
auˮ��:��/��ڛ�1�)m;���05�5��>c{
�B&����uM��n',��M�QC?�\,s�&�����PW��ۖ:��744�S��<�,�@=m;g��tJ����
=+b�n�vS�O�R�/�A�D�O�o�G�Ħ1�$0r{_���ғ1�V�d�o������*���v� ��I�����5��*�q8�E�穈G0�G�E|;�Ϙ�V��4K�����t��Vi���!�j�Cʙ�}�cߖW�u��3�񣚢2��zA;vX�Rn
�qt��U���w�tۯ����P�Y��֨/B�LR�]H��H�P������M-�Q+��Ƴ�V�׬�lL.��²�*�Nv�����ξ�YfV���ﵾ�a�0����q
/�c?���My�.z�,P��x$�]�bGqZג��o����$��~ꊡ������(rU�Kn�G5R[z�f�i|�|\+=&����r�9m��G,9���4Tk������)RM�c��Zū׉)�_��t��ۢ�yF�v���	ʯ��To�%�#H��T������q>|�*��6��5\�4��% F�� ����|�� D�+�5f]Fa Y�k�;������o��?)+0�q���_�PE�aE���ē#��ʄ����e�����o3�H��$�jG�����(��>���h�dO�Ys�$�q��/���������\	�Q٣�����%�(8�b���4o��I�Z���ۯ
���a�Վ�(��]��4N��{2�O�Dvi��S�ʧ|�5 R�Iy�NW���𶧋�k�凾l�]�C3�����n�౫�����-��v'y�L+"Q%��_��L5�ԐҺn]5~ W�A���&�}R�Kz���np�J6
����π#����f�Q�CW�� Jh)����v9q�.��y��q(WZa��s7r�G�P2b�Ex`�N7�7��lP�N�N��G����
�Ju�fM��T�m��)�r^}C�y�rX򲺜�GEE�~��w��/"s�[�K�~}��vdڍ5�U�o���uw��
I���$��՝K�C4��)|7k��~�d��_�ԍ}�\��|aN�OF�w��ɻsQM��]o��L��G��\f�&��A(�?�p� �\�|��b�@q�����׶t�`�����q^�p8oM�"�4v�Vo\xO@d���+oM6�p�����!�wGq�-b��\���o�r����cb�|ps�M��H���!A�tW�#q�I�|����U������>�|���j}<��I�S5����ؿ7$&q��� h�YFy�Kt]��+\���W��k�����U�e����y�]�|�?f����I�kl-����ձ��{�0�t�&Q���3 4���a��Q��i�x>�Ŗ�t�~���o���f(D#꧊��ˌ/X�ݐ?�	��ױig>���&�,v-��~>fT��u�1n��
l�TP@�]*q��Ђ����/4��s�q�^Y�Gʸu�q�^B���~�->�X�M�>/��a���SmY����ǭ�f����.?��IeI��%'�O�Ԟa/�zc�~z'���[a�T����Q��Jb��	��Ώ|�G�?s�R�ʮ���IR�f<ƻ	_��8�C�͖HC�����$���h�@W8��&Bւ�w���+���gQ�x3?���.7���9�֮�έf����&��ܠh���km�j�2�T�j��4�T��� r�<K���4`��,ű��bK��E ��O�x�å�4uVq�t�eΑR��#4a��0�Mt�7jEO;{$��jr��.Pg)&u�G�ؔ	PlK0k���]η�EB������=苶��(�h�9����3�8B�9������`�w$u�uzu����i��
�v'i�����W����1��O�!ie���B�����=�9t$�c�M�w#`�~g�Wt	�Jf�Ҭ9�oj�� W�����%t1Le��X`�&ZON��qS�$rͫvkP��2�P<��Q%����- �a����J����|�>O���_0�J�}�����ąm9�'����I�B���	D�[�T�r�5>��o X��p�Tt��UH]�n�ށ�r$�0ztƾs�mYE̔cФif�V�O�ћH#����J�1�z�&�=:D�}ʡ�	d�0}8B0"����Ä���;L�N���� ���_R�w͉�w3��Ŷ��%(M�fi��@�~XX��e��t��2R�z�y8��"�Cf2�����, "����~pv8����򪥋���wP��:����qY}G:��Uw{Y��a������ⵤ$W�x���fSS���"ov ����%��>�0��D�7��� �}�NW"|Hu[1�xm������9	)�1���I���@z3�K��|�B����umZRvy���/M�j3��k�Rܨ҅PR��J*1p	�W���~���sa?`�w�����K�r�F]����h��Z'af�5Pݘ92�]&|�T�������p��mV����k�Nw�0_c%*=W(��tE�K��f�X*���[����	������ו�K�	J���(�R�B������V��>�{@þ��]��U��J?�.��^��!��WBw���%��PG������ʞ���>�K�|V%�j�@���/�U��^�p�Kr���YUʻ�����}tf���,��Q���jwܛ���o��(w+|t���CZS!��i���^6>��6�N�$]Z��Ĕ�U�������F`��CL�J�K-ȟ]�,y���`��w�E���_�v
re�m��zjw�C��ϔ����po{�6J�QTߺp��J��;���Bh�̊?}G%F�W��SV�%�ՙh�Dk_P"�ǧ��t3��
_���h��".���V/�hIX{���rk�Nq�Cc������X�'p��S'��jä��SX�?>�H�)\�Z�)ַۛ��;6BF%v�����i[Wc`J�\���#6��AK�(��%�P"�X-���k`��;&�ڑ�4��ɯ.)���L�<K��c�u�ò?n]�%�^n��k ��a�iJ�&�������9hd=T���q��q=�f:+��!��J��{��f�WܮӆN$��_���k�:f��k��Θ7��v����^U��s*\T�	Z%W9�����'�+�v��8+L�=�z�o���8/;�gn�fҰ\l���̘��QH����=Ql���L�t��� ��߻An�D$GZ�(<P�]���(j!�z��Nߗ&����i"�C�I'�7<m�!��2Jٵ8��w��"V�g"C�P+av(��o'�~�~�2��w��(QbO{[�~o����&��I3�J�_�$L���k�Q��і��k��_4�M�zd��t��Y�
qh�G�a�~وab\�BTy1��|�"کV���ʓ+��ԭ�V-��n����;B��{V���`ǳ6�E�c�%�c=FfZ>M�F A�֍�s�T�P�0z��2/I@'�@8�F��R�f�/��k�_p�j��˯�ܴWg�� Eؼ���FI/�	W�0W�E%h,�8�%�dM��|�{�w�G.4�~��_n�d�!��5Eڛ	q;��-���T�Փ5��5uSAT����c�Pfz��>��L	/�OĻI��K���x������&5���V��t��v MɃ��:�p&�6���U�w~�I"��=�C�Q���6���5*KV�V�L��ϮW��5s�Шh��4�f��aK�j�S�9�@5�������]�Տġ�[��VF�\���,U�щ�I�&��x����R���4}:k��� u��[�@�~F������:[%�ea��	!�j����\�q�&�޽o�D���AzF����=�ÛI 9o먇���\�Xģ�"Px|�U��k!�A��lwp�4�vO��C��7T���"�3�5�a��� 8�J�q�f��Jc�YȆmC;�9S�����s��\ٞ��~ي�Qz�҄_�q:t�?3����) O-% �N�\X^k�d�
j97�M��a%:�ʀ�e}�9�nx�m��O���n���_d����(tғ�]���s����Ϸ�Fd����j�����^�1[iP*N��Ϥ��P���tu��|��Qp ��:����;�ް3u�ȓF�]߰�"r,��^K��`Hl���6�O5M�$䛴o�}�:��Ԅ��U�^>INT�L�"�+K�&�na7f�z�:(/�u�k��Fg����(�B�5�����KY�ٜ��HH`�<G���v�Մ3Td��깙�"U�{^��,��l]ZS�4�USwZ� ��x�b�Z�y�4��*Y��ʊ�oL�ݘ��'�O���R�*�/j��۵�De�3k =��΀~��9����aVt軪y �%�Ə/v8�QM#��~U}2M��A�bh�W-b&@�lE���'��#2��1a�g��@����_ќ���O����px�xƚ�~|{�*�)�G�3�uz��P|�QG$O���re�uK.�B3�s������d���9.@������"ى)�<��5p�_b��*��Tz��WO�H��v�d� ����63<�B��pז �Q�s��F6�*�4%��ۺ��sW����@~�z]_%�����87R��*k�����G��ޭ�i��z���6��]��x��b�tStR�DG�y>�s��鶵mf' x��̟O1�B^�p�~2�S	-}aip;�HW�
 ��z�>":̖�@sAR�z-1�"�̔S�s��E���ϝ�@�fK��$	��!�<q�dr�IW�6���x�E�����c��ŋ���'iU���(!���A����|��Օ�*'�r�Ґ�J&�ydD��xbZй�� ������-���t+��M��Ī�ZW���܆�HY�8v��X�Eԙl����4�p���MW�y�e$N�;��(�=�(��S�	�������9�5i�n4iY��9���stbDV��}��d�y�%3.~H�%�T�)�3W��#3���-5 ~�.�1Y"��Y�|�b�%�yB�E�t�*$:�!�(��]�FzĮa-U ���]��Yդ悄ڶ�+�z�s�COI�	��Q��#0ϋ�}pH�bb9xԤJN4y�����I=���PM�,-�x{����n�%��O�@���H�4�
�4��M�,���r/�.�����[p������W-�W���U�xj|m�!��}����pE�D���!�E�w�!��ٙ?���FΟ+���UW�T�:x�&�9ͣ���^z?�;>��
g���n��n\��`��@@�
Q����"@7���h�zB�ޘ9�@=R|MW��|3eஶ@6��$�S�BU��xb��(=�qﴨL�)p;�"T�����;x��HϠ�>ͧR��cb!�{�a�u`�<����yW�*.W�lL�a\�a0[����;�ᥪ6�a�ӗ� ��q\-m�_^^�a1w!5 ��]��p��?�݂"�ƅ���1��+���V���-�`;ӑ2��.�г�C������N�6���Ղ4�,|�R��xV�R�>L���un�G�\���x�7qWX��'ie�o`nu�I�&�l�sP'*���`K�>z���x8�7i����^�ըD�(��q����W>���b3!�%R�d��C�]8�v%��ܔt���=�a:'�����_MM	SɬGqDO1~����b��$!� ��Gh ��]
�s�-H��BF�^@d���;᭣H��E#�dN��f�5�֫E��(��2�S��
�b4�C-�p����[O�O��F2}&��	�E{FnDX67�ͩ|֙3�g��͒v�����_CR@} �`�^=d�bn�0k]��#��;�0gr�|`�����H����ʔ��F̱���ۉ��o\��fH�=��`�X��p�lD'4�p��*�[`�ݜ>@�Þ�u#͐�� ��G��\Z��>�nM$��:�μ�ߓ��vFI��ef��-Q�q�yJ���pA��<v�{���5����qٕ��Ȟ�+z�4hAp`�u`���u:��4���4>~���]l0���)�5�O�E����k��e
"[�y�X�BJ>V[u��Xp0 ��P~��R�wZ�j�ѳP<�t-�̾���}T����H�X#�R$��:;�����-����}�Z����T�f������� �]��|�Ǎq��|�"�gi�gVQg��=�J����X`��L7�G��V�6�g����'�^T{g�Y>�Q�a���vW��J��Т�H��4�R��*���c�Y�� �ӥ��J�p�h���~�>m6��WC�eYJ�T�!-+���QqU�~��@�v��:b�h#�f?����-���ѫW��㱻P6�Q���r�FgS^���>Q�r=uB�$�:���� )&�=Y�~ک�J��ڞ��j|�ŵo	%�!@l�[[������#�+X��1��(R����N�D}%��w���K�A��e��e4g�oN��gCj�(����9��%ѻw�hP�
�u6n�&�'Gw�27F�,2�2Q�#�(m{�O�]1����{xw衈��W���u2��(g�(��-�����";K)"=�ۉO���l�D�9o��׾б;^���Z$�A��X�b/=����f��d[�͟�Ø9"r�H�?��?�H�Rv)9�϶�R?~������1�ؘ�I|
�:s�w�~h�jF��[ld����8�M�.��W放j��r��5Y�W@�ho����u��'(D��Yxe�p�su�'D�kTv �_�w{�C���[�>����`�z�.J\��{�}�Y�\<��k�q�G;%�ư�m0-��~�q ��k2�d�֮��>��b��T�Je����<)��R��r>�LH���V��TO�؟�+��cnI,S'S��a3 ��/�)�xq�N0�����w���u�1q*���	���&|����+�0�V]����!Bb�lf�������R�,�%	/�BcMf��TDt#��;�ڹ�6��I�H~�f+T&hM� �Y�5DC�6�kVB���m��}�]F�Rua<��s� +I}B�fz�"����b��\���&وG�V�O�POрFsϨ�������Ռ�8��VN��cO��a���Ǩ)�K&��֌�r�&1��֚���7{�3�%y<��`��s���y����C��M5n�Ml5��)0X���!�buCѡ��\�� �,��h6>�,���;Z�@��0'��\u5L3V����Ƹ%�_��!���<�Z@����'�o\2���~2�:v�j�0��@;H>����;�Y����6n�Px���ͥ ��Z����� B�(�[+���«���qYW2ev�Q4�x��[�1~o!�&���##�_J�{��?�٠�Ҥ��@ۍ�Cm^!-SpŰ�0�桞OQ�x�d��3K���5�����a�A��?�G�����gc�Jz�x�y��@Z+����c��cEDe䤭�`Ȣ�؄��i/�ܨ`;~��1�4L���:2V�L?*��9i���ϳl���?S�&O�Kɱ]�/ T�md~�O����W���A��6�A܃-T%�[��itb�*uS(ՕA�/��㝚��l	�b�:x�4YH[�#\�ư�)���nO`	K.zn�v4��H'\���%:)��b9��4V��	m��bK<v�7k���o�Z�C̉��f�]���~0�gԟ0���*~�����M�f�ˬ��hNF�P2�D�O��\m1� �c|��4�["t�F�<� m����"�������0%U�p,3�٦�M֯[�X��U�Ch�g�#'Կ�duN�	gr�8[�pDp����ȗU=�}��9o @)��>����z�Kl�ءhu+
�/��H�{2����^ ��2�2��鷭6jzZI]B��t�u`�����Za)����R��L�u�0
E�}���&����&W�q��"�@2�����*���
bBaZ���q���x �ftο�;���}���k��.�^4���dr%����_�T]�붬aI�"F"���@<{(Q��1��*�h�/7Λ�O�3�aaAп�i�; u����0��_+��0;��6��x��y-����QJ�8Ǵ��:obx:؂�!�����_�`u[^s�"�)�Y]9�m@��6iVJE|n�ENK�K���tҔ�13��F�O��"(<��I6�S;*F���B�LgN�������ɔ �	x�Fe���W�"�
�t�����t�9^��Փ�F�v�BG��N��ׁ�Me@'t��_g<)�?@��yV�a�Ċ�fGf�޻�R���>�>��c�;�Qg���`�)�6��t5X:�6�j�CH���fJ��{O�7Y�]!!'Q綼� �q%���[��uH�r�`:5�}u�
�3��r�WR<RX��Gj��j^,4�7�K0aTR���,KZ�I�S8��L�W�<ub�Wn+����\�H�P�i�rI$�"{�e�Q��<U�eo��$ؙ�`�WC]eo����7���z=�j%�D
E&AX��y���s�1x��qR}�ȻNWK��Yq�%Kk:H-�.\���'Z$��&d͓: ]�f���t�Cj�� �)��� $����hg��{�����z��јR�l���h#Z��-:2��rk�n���p�3=Я\�7n�_�u)h5C70A�x�s,T<'�(�o���� ��`E��>��wX�_��R�V����I��O�n���O�I9��&���󩉽��D��Y��/����eȼ���Dj��;��
��nX{� ��N�H���	��4��$Y�L��ŨD. #o���4`q_�!�Ů���.xhT��o� �W��J����W���B$k�@Fz�ӹu��`��L�㫜&����S$��RVOE`μ�8l���X�xA�^^҄hn�>ё2;�G+�B�Ћ���l.}#�A����9�7�Pʡ��j	V$���CNQ����N���ܶ��ː��޶q�霗 �%���~�R!-8%!WaI,T.�W#�>}����s���� 1���$�`-�&�җ_ce���Pb��E�^���BA͊)��XvA�ɗ���i��1md�#���c�|�]��#��=�O�)���5M�>�#��L���6���]Āh���V&3��ԓ=��rt�ּ�����,�'d�@ѵ=�x�ՠ�>����t��o_q/nw�d��F��e ꆎ�S� �o	�>i��@���L!��e��l:khY�A����b���u7%U�܍@��H	\EshH,t��)�,�W&M]$W��LZ�W�b�r�$�j�-�9]����s\h��RHCp��oЅhQ��b�wf�R��P�f�+mnF=�����~ɉ���K�[��ywT����!E	u�9!G�C�L
md5�O��M��b�'ta� i T��ǲY5^��� �̱�ř���h��<Bo�������0G�6AV	�%�#`��U_A�7�"�T�P�w
*�ϋ��d`T�a�-��f��ñ�]�`U��m��U�}��"5W�W�G�t�:��U�(��˫6E����fJ�)�M��ݚ6Y���j��AƦ
��BHɩ��>)���u٫���͒�3��:�yS�b� �d���+��	%�V�ԟA�{K����M��|��X��Q��q��r1�D$�*6G��c.��S�[���\iӍwf)ڜ��Ku�3��~0���r�^ ��k'� �˳�
���,Mbl�uL�˱�:0����+���G[��p�;�"��C����Aky�������3~ �rAlx���,��jdH�k˞m;�ؒ����w	��o��lC�0#57f~�D�I�})���}�Q��;���4lS�s7�K����J��Lr�`�E��^��i_Q_�NŹ�p4��򀯓Y[a��tpPm2G���k<��-�J#Pi�ӹ4�`Y�h�@L�E�=�?��E0O�=(H�KRҵ��!��Z�*�k�9��LѰ �J*[���ԇi�P�#O�R�%�X������Pd�nj��o��d��(�����V�z)��{��=�V]Y#Z�"��n �b��xy0L���Q��ڊM�sK���8w��`�p���C�=�aQR��Ӛ2%��N�Λ^ST'��0������p:�o}�hz�.�k��r^���	�Al�R�]T#�K��2�}���R��vUB��7��]��]L*N��6�e�6���6�/�~� �nM�@Z5�#-ĸ�<�A�D�N�j\��Qo���C�g�ު�~�U����$f�4��.�R�8�KU�E�y��#7�DŁoq�P�����J�|�Nk���+u1�\P����5�n�7�F�>������h���P:zQ%ڷ�(v]�HIֺ;;G�M�.[E�^#���<;{˕���9icFR��W6��[&c���O6��Mįb�ҁ��/��	EG�&��;���xXy鐟��اd햤�0�e���W���,%~5;�4-q ���Ƥj
p����� �Ƴ���Y��/��9�}�Xip���U�6��v�Cl�D��37?��[>kc{�Eh���T���ښߟ�!!��8l�%Ag A��ף�·�+a.�[z��k��ӟ��+�	 э��^kq��ֽE�i�)�� z���9��!WTV}fF�V���)���֏�y��j]g�Y�e��;���ﲠ�gwjY�&��d=#<嗼[�����CpW:1?��7G�s��0�D�t�ww����Io}톕-e��f� �~.Ə�nԐ-��j�r
�Y�Ki0QJÎ�!tU�����<�۰ uwM͎��x�Yz��l$�n�P��$�4�ϲ���]�A��L���2��Wt��{���l�%)x���FĜ��MvO�4��N���(�.��7�H�~�ɄD�NV�a ���ӛDVp�dY1��w�H}�#=n�&�y�˂��)nI4�\廙˧xuB�~���Ƅ��$���W��>:v� '��^��;�4OA��-�p�:v�v���^�4�[L�W��{�n���a\}����P���E���h<y�2��Eu��Pz�maET���7&�e�raN	������Q6{�T�\@�aN��JO��z��K*�[W���w��*�������y{Pa}�z�CheOp���^�����Sk�P_�Ғ�j�-ڐ�K�$�RM����i��Ue��g��+^�_�!g�̕��l\�g3��QWE��\<���cH@��U�8lR���i�����=��jjGc�.C��|�c{���5Ir�ʄ��K�x��7m�!�D�$sƅ��PO��|ʭt�\"���Ys�ߵ��TgH��ݖ��!PX��5��=VuE�q�� �7��k�׶�Mυ�:	�:j�U8��$�p�
N`��˝�:�!̙:��@w䪿���gnᑠs����u.Pq0C(hg׭I�_8��v(�h�΢��Pfv ߼�$��x�<KQ�t�
��}D�ת�����4�`�\��3��K��z���r�1�v��$Hv�}߬nI�Qㆤ�H�78߳��k�� ��������ʀ�u�^���F�a5�f�`D ��D���TQ*���ޣ$�'��Y�E�r�c�Y��D�Oɿ��a}���lB
����׈-�
�7��Lݳ�JtA�Y��}Z42�}&A[��lt��G *u�b�ԋ��)4�e#��bgي5�R�M���n�;����q�G������Fz����d�.�H8:"^Vta��О7%�@��6��zѮ>��>+ѯD��N����QAhSO˳����-Y8�ԪgHIj���,���e�{�H9y�[��ɭ<Nڑ�Jt�݈����J�	^Rņ��Z�D觵3�6B5�h[`W�Y�L�7�5T����ά22��"U��4	�dS������%ď>#Y��^�t�z!����ϥk����Lo4<�;��,k��Pō��y]�F��7f�y�x��6)��C j�P������n�W�S*�2�OuD4�8���*�<�����*9�{�����?�������6�K��������Cx9����~�.b�����V/;[W0>�Ѓ���U�*�C��Yh�O��_�Y�c1l����92�tB���DkUkp�,ԼnbO����*]�l�p)�"�A({����D�b��t���n@�����T+����To��6�ԛ�`�f�Ə���*�H|�`b<&�G���iEN	������I�UJݠ���T���հ�z1�B@�|
��CW��g}�/�a ��>�S���ʀ\���Aa1�oꛊ<LyӪg���P�����G��>jy�H��[kƴ�_]�7ĵuQ����,�zY��:8�;�{�C���-3u�cU�̞FbH�����U�E^���π?���+�o7�t'��888(S���y$�W�������������.}�^���|�� �oSY���:VƔ�N+�P�Ʊ��SL��?��
��N�ǩ?��9N�cu}��f�J���j�eg��&��
�B����������"�����9��C�i6W�o ��r�߹�f���sJ":Ҝ�Ƥ�Ʃ�+�l�����~�U�V�L;1���]�)���.55�� �/B�����`z<���Frg$W�%9X��ͱ�k� �t �����fCL�_-
�����ty��!4D�L��tZ���Ј���}�`LPf{hB�_�;-�aFEFC�,q�*!�~"�ъ���\�Z��o^u��&��:�\��.0�Z�e�SQ��}B�`XeW��Gz�>��,�N�d���tMA Lb܃��Gw��/F�7Sa}#��lz����O#+���~'ph� -���5bCMkrs`h�y{����V[��N��/�L�`e(Ɗ���Z���'�KU�2�qaO3��r,���
�;����?��?u�b��=���s]$�����*8�zRwT^{�GY�z���]�?©v7NM�௞z�&��N� ?4u^�3���u���A��=ٞ�KU
���L��XW�.4H���z�3��@�s�1��n��pm���2t�v�ѱ�� �P�T� ��-�eS+�Av�#����]#��<wt �9�>��r[y!d�Ҽ�M6�3�߈��2(��i��2�qD�+��=�\��mUV������9�@�:v�E��n`֯_�+ݾK u�����j�}�U ��
��)KIȔ�����W�I�&p�G�Zx��5�l������R9�i��$��.�mNB,aow&OI(���i��j�F><��@�Dq�K��T��<��P(�.p{l��4�q�e��m�)�@���v\�#HQ
�a��ĉ&�M�Ӿ�=��� E��s�{&9[�!_6f6�kry���)_!��h�hw�ZX�Q����e�	�-�=сܮ�M�}�źb����/j��@9�(��v��P"`Ğ��F-p�n��ې�������(J�7��9 ���@NF�5��i�кT"�J�OM��ʏ��C�{�L��!�����V�����j��~]~O���y�b��3d��q^ף�ëAˆПd��R����5�9�:i��)l�3���*tR��m/�ι!�{�8���D�4c�h�E��g6��Yl����/sx%0�P
�̭���5��B�Ħ�yB�U���{�V�DοM�s��M�+~mV���%�h��<ӦT��<A�GJȮ �ti�ٹE��cF�aW�ς�)&z��%Q���:��C��n��҆��u{M0��,��Q{_s:	�.{D�q���ijL>7u2%��~|1�U�B����	Kea���O.j1�2'��rh ͳ�v��C¥�F�_����Y�Q��V�!�����98���y�a��-v�n\�m~�|�w)p81�� �|i�PA��t�M�a�<>c���E9�X��Y�HʯӒTsI�c�5�TB�"d6�OJ��M��p[�B_�
��T�ya#��+��u�~���OdBҝ"���%��PM��[Bt�AE
c� �b̄I�O'��)��&���톇y\B�P�2�:Ier뺊�6ħ���n��T��D��o��7E�'��@ð��0�$��R[b��W�ڶ��,5��d/�)B��S(a(� !p�������}7��L&�BG��vo������0
=��N-`]ͶO��]ܭ@� ���zj�W��$����ehS�Ć�P���DӅE�� �NT \p���J̈́w�\Y��嚰\.�5�Y1F<⎕�� ���D�[��'a4Ύ�s�|et' u�3G�G��I DܽT�O�8c�=�yEZy��O�3e��F��bP���솢��z�~v��.��l�0����din�1��}�ɤ��;*���wXߝa a�����^1�w�0�h"�]L_����R~wEjD�6�����M���z����q��XM
n����pSf���4y����[1�ի�wb�v�M�Ѵ�,��E�,�3�m�||�c��V�����3��2-o�KJ��8�ݽŊ[8��ɒ`dW�=$�0Y{����X@'NGa&�������ә�T1��ٳ���!ׁ�B;�9�]-�
Ʈ��&�w]Ǖ�q@)?2��.dߓހ��wӊ��d(����7ȗ:�C{I�f�oN�>�u<I��6��r�%En����u���VT�|��Z4���d���rh�|h��@�<�����c:_ZGn�t�����s;��T޽o3y�|�}�f .z��_	d\�P��+����Y��Lǟ�kAU}�M�4�d�{�˰P�6:�y�{��[�Ey�Ʈ��!h:+�6�t^P�U]^�Eu���5\�套P�����7�T�zCQ��u2�q��B�|�O3
�En_�!.�5�c�˜Xl��u�έ3ʂZb<�	E��W�M�r �*�l֞;aBJjm&!�
��Ut��������m��5�`
��=<�&��Q7/f�s�=%�1�����6t ����e::rIr>�,Ζ��1�ԃ�{Ru����`~[Z�Qt#�(���d8ZMI���F�6���/��=.��г҈$�TӴ���D1�M��<j��ٶ��
�)1��eL�{�V�Ǘ5@|����_�S0�$ؔk���P�;s�Z��9��ڙ�����<���[������@hi��(��<2ؽ�owa�b�����~��~��ҥ]d8Ȗ%���	Lq����;�18������8�*�-IM�p��5������{�{���aU�Xd �ځ��1����xiŤ|������V�|��?P�>2���#�2�M�%�7���XVD���n�]Ⱐ)����{}�~��UD�<Jvs�?�a�4kPc.�H��A �kE��_�-
K��lv];.��}���5M{Cώ}%��q�d�Ћ�mT�S/��2 ���D��aeӯ �����1qc��x�%�U�)� <���`�����쪥i���~�����|M��6��,���c��_,��}����i��橯ɒ�п^QS0������&u���k��v��c���\�i���J���[�,�śdYz�\E����?u(�eĉ����!�2�I����LR����J�����k��	p}0�I���� �'�V+n0��/�X�T�"L~/4�`���*;��gH�7;�_J)����h�{�����<�搰�㕢�D>?(��Lt��2!K}����{o U�uf�����*���coJ4��߁u��NL�h��!^�-3�oz�<
�d����(����B|����qްb
��p�?I����N��"8#N���4 ��g�j�;B��Ӽ�uf����@�J`:��T�6�g3�,r|�ܲ����E��@�NŰ�{���VX3s��qC�b?�2k�
��>����|��ZF�
��.��S��!�T?`����[�D�J�Cc��w���f1'��dV|G]�Ζٸ�@>�M�1�|M�Ex�̇�C��|N��[6��3}`1r�!ɔ�X·υ�?x�d��a��?&��8��!��=�C�;����o���t'컽�rW�Zx�ci��ϕ��ց�oom��l=+t8�S����m��:���RH=��v��d0�xͻ�ˋ��G��&��@N�B�+_��O���Fr3������O�/�=��k�E��H9pr�'r�7�8vgmy�
Q��Y@�S0��	fVe��!�+'9�]f,��#^�]t�o;lp�F�B:D��Q�[�^�+-����Ȁe/���cQ����fq�N��e8�'��g�U	sG�	v��}`5e�����E����u5�����7�Faw}ifb5�>�䆃���[\�o}��Qz��h�j+�����Eg4�u���C�s���P3��|�<J�Ʒ匝+�T�#Y�����'B�M�P%R��T��9�"��+��PE�\�f����u�1��J�~�U$v��Iq[�ձ�e=
qcf�Y��<������<E�2v������3L:hA1w�y�0wɹ���fz^G�r�yv�=jB�fg��K�`�f$���_��qp���p�)U��G��w�
L�E�NC{|c ѓ�^��ϧ�v녑8��B�q�k�h+��m�d��l]t�
��+���G�l**i^i1��_�řV?��"�����Hɥr�1t7�Nu	�K�
L��aw!V�JeFͭjT[�B��(Ţ�P~u&�G�K�@s�F���|�?�4�,�6�������\�yg�hj5���f�r�nԑ�0s-�xːNp�L�M�H]��C���ٝi������Ar�"_y����<��#י�A%��H]"(�(#�Xv|i\O� }R��]i�MlE�Š�VoY��I"R�ٍ��M �
���nПZMC��d�-�ϕ���kz���LwLe�$	h.�̵0D��D�H�W�5�\w,�/�,V�Y�/��p�ܵv��h�a!��ZF{��]�e)�p̦#<�+��v��>�ȸoj�'���e���[cؗ(�Y[M����<�_Y_s������m�."��׾���+ WW�`£�kIk�\Ju)��d�Y���"&� ���V�e� ���m�3u/pk�}��<��S��9t�*:_ԘxY��P���s��8	n������ԏ�!F5��P�UBy��,���p7ξ�/8�(��q�T!*P0?�E��3.1��&V��W2��ʋğ� I�
F*A�ٻ2*��`|&�:��Z���<h���Hi����_!��&�8nj�;�!��:{���4EFt���6|�s6)��1N2�T��8��o��A�s�%��(Ap^�v��*��w�裟J�U��ϒ[	�	����]��}��f�}0q��;w`�M�]��[��ퟮ���ê�:�[&�Ĥ�Q���/m~YJ�^�I^U��71(�cS��"P��F�8)�OԔ[2�����%p�o`���a�^"������HA�y���w���G_��.�9i`��,R&��Rp�wO����gG�"#:���jU�d5�r�(�ٟ�2�ŵ�|���EL�<�n��(2�6�P�A����U�g^����!�D�f���I��Ӟ��Z|��A�9�uM�w�Q�G��˔N'�Vv]6��Z5�˅�-ts��|LӬ�A���`�%4��li���*R�JKT)2�~��ڼ��O�V\Vl+�
h\e����#؟@��ܞc�r�O�8�ήdWQ �i�Q^[�#�P�@=��1"w+�ղ.�b��E���LBH�V��:$�.�2=��݋�m�&P����h;b+bpiiN��6H�A� {�ˎG�����`F���hKe�)�Aeۚ*��x��I+k�V-a�W��5����ṹ#��C	{"�Z�o�F�jJ������V ���1nګ���:(5V	J�tJ_��g<]L=Pb� t.����(�f��]� 	��f2ـ�Ax��En�����J�E��e��pH�
���px�8�������H3c&�W���63? ��ؿ�R�ﶴ�'^���ۺ;�p:���kc��׆���M��Չ��P��ea�~�����	�O��_�� ©��?IFi��P翐h��%s�Rq�'�#���*��3�N���/�a^Y���*�@��7:��H��<+> �O����Z�ت�2�[���a7�6�>=E*��[��C.�:@�@t��q���ew�d�d�s�(��8M�?�u�o�]%V���$G���ԡw��u9m>�`q�9?8��(q��(	=dG�\�� cy��DIt����B�����R��Y��?q+�?�9;)?7��J���IY�Ȉ��&��؆���)��]��`xd����re�0$���7g?��<��7y�+aG�ا�'-�+������1���b-�>X��>�dd4T��ũ�-��m&#������rqdb{����'���Ѝf���<[�H� �'�:�n���t0.tg���jb/�����ʧ+_m�+�#}��"S ��&�/>�Y�2�=�>c��l�RC6͙�����Np'���Kh��@�~C�-�� ݲL��a򆅻��o�z(M��
删$,JJ�9���n��$�C&?r�p?��/�UW��c�<��Ӫ��O�G|Ϋ�g��^*Uze��|�7�'�E������Ė\��_9�-�vQ��F��9���)��c��4�=d�z �~��'&J'Z{ o���WK�w$faL�d�d�t�L�������ʖtLi��㔜��\>��p��gR?.3�owu�Zƿ�Bgs+ac�Y[C�4�i��ޒ��:�y@l�����;��ݱ�\t���f��ŭ�/��n��^�=�ZT�s�h�|�k z<�g9�bv}!2�f���~���nZ{��R��l,악��qX&�4�4�ta���"S]$c>�`ĳ����17~`���xF̪��ұ�E	�f߷ْ-�YB1�]�f�D&�5'�9qz�^H����!\���u�@(�R���r&e*a9�ܪ�f��On���cۇ��M��+k&������� / �Ũ������.�"sH]\�īP��s S�B/}�Z�C�/(�O�J��(R����)sNH�
���BSʉ�%b���%8��7�Ɓ�� �z�6�)_8�������c�����EE�UZ�
��`y�K��;�vb��R7�իYjh�5�.���1�,yH���7`_�tS>�3l��]�ѽ~
�L%*�Y�6�(���?X���P8��4�
8p�WQ#���[��j�l�B��\��p"��W'p��?PJ*G���b�&X|)������TW���RliR�!���>�(���w03t?�p���~�kzZ���n"м�Ȁ�NM�:_������a�!�G�pT<Ƹ&v�Gw����;'���p�.��(R�-�������
�U��&[ۭ�P=������2Ь����(���S,��-	�t���xEՌ戀/?�Z8e�"z�4�!�T3R	.�Zc�6�r�SX¿Y,���Vh-�4�6�kգA���ܝ8Z�#�P��B�6�1 ��У�2�5�p�W��R֏Y�f_�w��Sr8f��5ɻ<�����Γ'h�is��X���dB�e�B+??�;�v!�.>`A����%��Q�[Qc�����(��������Y�����̽.��]���iKHl�Е��OC_{8Y�)@;�z��
�� ��t�n\KT�qZxꊡ�;�nz`�<�+��v��E�VDZ��������D2��*xt@M
u��m���y`���f���M|O0�̓�t�E�0��B�P1����1�ӥ��s���ŕ�QH�����-Y�?X�ߤ���lݑ�n5.���p$���ɖai��"1c�v�8��p��4&[���e���f�۞1��Z�J���,�ɳ����!"zp���=�	I�g�ݑ��j���<��P�t�R$��0m"LX8W�\* $y���w�1(���o)N��]f�;��QP Lĺt�0��i�rN�9��5"�9g���֜�^(29�]]��+ި]ﲽU6?w���x�t��HίR��9u�ԁ��{�R���ED[����Q#���l�2��g=�J��8�/��8�"���p\"2���4�p�&��r�<4p0�����?�p�q{_���!�ˈ���e�0�� L,�=��}R ��X=c^nc�p�o޾Du+|p�/R�e劅���
-�^����L��G4�`�u�wր�C��j��ůR�h*����юrdP��Ha�X��O�2��2J�`&.�}��w�k	�%(#��������dx�r��fm/v#��6����Ih\��F1$\��IDk@��R���3�r����2ƑPy���;��-qq�I�ˮ���V��-B��LQ�5nE��^xq/�r�ud�T��E>6�	,q�_C�nqN�Ehq!��6��������8d%���@��D�ޣ���~���	�q_���@ob���\�����[���� f�K����q��� ̥��KȤ��U��X�dFY�����=�u�m�ѩ]��B*D���*J�u�M+��E�������2��FѤ�Ó��
��3��y�A�7�{��X���Ӑ�U�'SY��1���
�ʔO���*���J_l�eb>��jx�B�U{]�܆	[h��QkT֋�m։�`�+���Y���`ڈ���4C�#sU�&+i0��,��6��9D��K�q��T_�t3��ӳɫUl��i'^����s����<�PM�N�߅ݕ�[~��kn��?)��Qaq�KY�j��)�"�iP��������e��!@�"H�Ns�O�LGNdN���zW<����h������}�]�s+%Yt� 'of�\�;����o�s���Dqu� 3\�۴>z���4V:��0>��lz��`L%��"Q�bN�P�-\�gT3YBW�&lK���"��;��#1"��l��L���G	��!�:�_����'(�g|,�Uc���r,��@m�^�Yt�P����(���٭z��i�t�`�Q^ļ�%�V�ە��н�G.��M�艐�p�c�v�jB���`2�k���^�l����`U�` �9P9��V�yG�m3�z�.��|�)O��2�=�𺫄�.b�<��o�!U��c�.��#�Z��x�/�hvVW�1�����/_��;�x�R�7$��5�H���p$h��N�����V!vގ��l�,O��ͨF^l��P��s��j��{��[��ch_k�'��=��nL(HN1>�&�?my��=��p��p��{�����#ݝ+Q�Q���e�3�4A$�夛q!YE�9d"vܗ|ByǬ�tLU}�V�됄u�
YB��B�J�E�BuG�i`S���wD���K���c�����&0\zk�B�[��Ć�x���mY]�`uPh��:6 �`�q�:���7����LG&�5i��F�+.��a)�C�	n�jB
!�h���(�4z��؅���c|~�)�0����c>b*����%��%��<S�,�so����Y��BE���ЄյUi7r�YV��]��?"����eD��u+�;_�c�m��-6iGHd�~�r�XZ����SL�#�IR:-�#K5��ՖMAلjkE��l7]���� �|����pL
3���|qB�Y3��(cw�w+#�<Up �_�rm�]q\k�ǅ���1�Z��e�'
�w���zT�R,�
�m-��g��"�3�=�?K��!�5.d����]�8"�y���>(�\Z��,�����߫���p��5����w����Ш~w,�i��K��
T<{�c��6�^볪��B}e�8'1���}��j
�Ȯ�,'��X�6��j`��ۖr��|C���@5w����^ ��r~�2�>1���Xّ�V�^�c�� �'i��V Ȣ�4Ihަc(V?D�ET�Qx�
�c��^F!ȥ���,��ȅ;��U��u8��C�=M�|���I�aV�)*��̤����M���Vl��TID��-"�Ą�*Q��F���}`���������u����O8���4O�����<���3ֺx�)~��ohRw~]{�u�J9v��c����{�'z��N�Tde�2� a��^����sTm��X�QV�˅��kg�t3�_c�ɿI�^�*���_%�䬔P|��92��a͐���
�x!�PS��qt���:
c@���e�����_����	��#�(c4�$��i�M��R=�רx�	�Ev�Cr=�SDB�����^0,9�� >ě���̓XrNH����-T��>gB8@�P�
�^,��l���Y�
\t��������Xz"Sc����;s�-U�+��L��Y��0�--�n�>��]�.hpr��R��G�7 u��R7��(��[�ڇ��p{��D��W:1�r|��7��ʶ��C+�����+������J�Hf�{ԾT�SW�(�k���?�iQɺ&��b*�Q^�m�����0S��.�)�t����H���(�	��p�rKdZoY-�o(ө��Ef�HY ����'��]3�)MM�u>�/]���y.�zNN��A��/� �D�u�j_�xD��R}�L�!��������ur�HU@p,|�k�ʒ������l:#��u�.����g�6?*=������T����x� �3�B!��G��_ok��C�L�Wf�V���g]�R��e@f�&�{�5S.�����M�R9�����ͨ;���<����d\��)f��o�v�|2�`�NZ�_�'(`�c鎸ۛu�V�b66|���z��.��":쾙�*slgy?5� ��!�=��
(���>�}���듒�Y�/J����"+�b~�