��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ���������	���u�h�z�ו]%M��i�qw��lY�(�)�k�ֺ	�ҝ��r4F.`�|�lM{`�!�:�z�f,^�>
�S��G���y��Fl�{wLb%�J�����x{E^?�׿{�^G�k\�~�嫌�G�3~�{����x���gj=���8�:$Sq�%�����(3�c˲c�7�e��)��s葖R"x|�͊4v뉑�]��b���?Oڐ�Sr�#���� Cl�-�3��*3�O�dY��
8�E� -�j�خ��d�/�R�8迏�<S%���SP_�C���n��6)���x8޽��z�W�6}��Px��^�h[����?�K�u�-ZZA^�/�"hu<?�LVj%E���8Z��,}�l^��)�Q~�1lk��3�F�7����;��@5)��N9o�)�)�T_v��A�B�!�W�Z���G��0��3 ��Uj~�pZ�#Ib�L �挦99Z7Ƚj*%���r~��"�xQߤ��Q�!�͝U#�Q(ӱk�C��p��
�w���`{U�q����J4qv��w���T���H;h	�%��Ł|����iZ�(�d�v=�_�
�a1���z�z$m�*ash-�Fwj\�J /�헬Ä���_���>�=����	ì&�'l�oG�@'>ܞ�!2��L��e!�n�H�Y��/K�;X�N�A\؜_7J�zM���F�\��Q��_K>D���WG�"��s$&�b�GOB�d��=j7�tV�����\a��8Ic�0�',���kv�ǋ��*Ŀ��Ҡ*h�ۆ���U�|(N�6=�H����+Y�MC�*L�&KK6<I}^��!C|��~s�U���bTb����ѐ�p�vp�6*��v�g�n��S;\L2l�~a�F4�L����!vf&ݠ�F���. ��	ѭe�kՍ-�R��䢦���n���w�[Pnب(���z��2?&+ƪ0�R���v�%
���l�ِ��_|�gd�8�d}@#������G�'�ؗ]~�wQ�s���d���#tcS�����u�me�̛<�-֮���L���"�n���/���c#54od�k���!W�(�S�0]�mku�$\O�]����Mf!�<.7U�bU�����$�1��7��|8�罧��D�kO�J��_}��o�7\y\���0A/J/+��'ȽXS�@���q�����-�|������~P���*����-�
_��,�]ۂ�� �4I@n���C3��J�w�S"֔o+��qVLt��د[�s��? ��`% ��	�P���J���������X� ����
�V/��Ρ����g��")�MkS	���n(Z����vi5�8Hf�'�Ej���/l��W�o��.��dCDT���f�H x�����~����%�����#�WEqI�Dy4��^��C�JC�S��z��*�-�I�;%p=b�����b��T�F�lF!��Ï�W���6���+�������l�>P�sʸ؞�$���Q���W9�W�"��m����4��?+�d���	�p���fl83�3<_w����?9�wz�ʺ��vT����.Ċ�[l�޹�8j�Ǵ>��j-T7Gn��(�bh�Z��x��ߠ�ܗ�3��w|�O=��k+&���x4n&����B�Ś �|2�py/��%ۛ���8�nP����)��Fe	N׮�x��D)��{��ߒ��|#a���5Й�����H74��.};�SQd#�NL�m�F2���7�����XH�	>��$b?qI�$b c%��9�����A4��mN��,tR����C,�@j�u��v��,����!�Rb7lkHi5����l8���u���X�m"�sj�	�<�r�!���&���-��\�a~�dQǯP���2��m~�Ĉ(��Web?f��K���q��	-��{{_y��F$��I�F��r�x�i���
y&��a�+k$�<d�J�N:��v(�{��z�:��B�L5���7qC���vјc�g�����DI^Z^�ל�ds\���Nc�;3����� �3(A�B�Im��Y�]͏YM9=�im|� {�'�I�S���0~�&Y�)����U&GX�_.��C�]��a+��UI̷x�^M��9)�5�.8pⅷ^*��N�&�	�r<�GL֍���3�ݚU��	�-^��v��|��P�O$�)j�y{T<F:�E����UV�7떚n��l��V�0�����7L���PIx �5o]�L��h�P��6��G_��$�.���@�P�_ETx�o5�Q�ALD4/��,�M�a�Ԗb�߲�w�:��[�^��v��6�7��v�z����0��M��H��&�_.�-HǚH~�A@__�lQ��d�`���vt �� �z�?nZ%�g�	�3sfq]�$	c����8T��Sn ���0��%�-���@����,$r��9�3F2Ds�,{8����|R9w���A,&�~$f�h~��))�ȍ�`*�g��������(i)RU���:D,��K�1��}33z������*p�)|���տ�B��۳ې֓�;E&D#���9�k^���_p�*L h
� E\@�T�`$I( �=�$��v~�F?a�	��,H��ٳ�Zbo�y��EMC��򩢬.JW�yē� VSSb��KX��In\�%��,��66]BO�$��>��k+�-�1H���N(�N�X� �B����V>�1�%���lI7Q�O�z�f������$y���[n��=w�mʓ��RΛ�e���<h=2�=��C��+S �uM���1'�~�����
�(Sm��#�qfv�,s�G2��e[JdVbڏsn1�B��ά�B��eM��V<�#��S���Wm�Z]��*��9t�Vc(�5L���ʋ%�}摌1�x���y��ՠE��P>�Jpv~�	�.ff�A$��=���΋��6�V/%?�!�㝞:o;�K��IO��g�,�d���'�d��}�����#�1�����3��"��T���5����v�k�3m�3�5;���'H|IO!��Ἶ%�O?�����e.f�����sl���V�~�v5���W����:�oE�����]j�������-�'���v��؄�ӦlkaAQR>�9����8>q$���6�A��oz+[�;���&c2�5�qhz�ڲ�F��j��S��LI.0��0�@�	���M�_�+�OtuC��4c4��\���^��4�7aB��_82&TH�k)�	x�c�ꃢ��=�z	�)#�
�4�ʎ�b|'�]
�~ӛ�y(�{䯛!���xF=	��!���&d����Ѝ���$��aЩ|�tL�"�w�(F��٪u�01=�^����1��[��;��>�멒�g����%���7��'�Z�6��)b\ �FpGN\P�0� V~�z�v������;��y�N��|��������rN	~`��0,��la��
:���~m��%�EC�=�����h۷���݇��ĆG9,W/&'�Q�"8g���#1�&,?9���]0#�]���I)U�V-f�%��@��f�0l��݋5��=�Opz�%cx��kp��T�[6+��6Z<�	�7��J�d�9[��5�`�htl9T�:=�*ԙ���!���ʱ��t���V\X����};�{nK��ϫ��4�}X�w% c��/���x�d�X�������nW�%�C�$�'tP4	�~��CʾS�p'��@a��0+X��p�Uڿ�0��+���ձEي_�"f%T�l�v�j*߲���(���9�wmi?��>��2��W��=�!���F�uo�A�o��?��]N�؛��Eu��F`uꗖ>��� �����ث ��3��́����A��ah�mx�q�N�A�I)|�X��>� +7� 6�*ؾ'�P�?�r����T�1)T`+�m���ө������H�(� g"#,�+��5�y��.H�;���_�a�����Y3�������.���.���)��vc�?΄�T�Ŧ ����!c�h�2���t@N0|_Q}$���<��֏U�X��KTS���&�1 aC��h��?A�Bd�n������t�5�FF�N���ת<�-�Y@}��F1ws!&��:�!&����b�eB�*�Ҥ�AB��*S�m$��42��K��ᱟ��ʗ<	�v$�2aysCl)�j�p�2��J)V`��S�fxL��E@�g
'J�bi�	��Q���j���P��Cn�	��᪾#�M�3�lL���:��$�F�Q�6�������Pv@A��IaU"�n��Q�(;K#���z�B[�0�rO��AU�kv`���7�W��,F��7Ƥ,o�%��z�X�19�`e'�W�/�+�2d�H���?�J��R�|�$�~C���1޽�B�.��k(��O��˴%:`v�d�j�D(�S�T��6���A֢��ʓ���H-V�|Ӹ?���� ���	�[HI�Y�K��k�!Q�����*b�D.�#�����:�5Z�v��=@����$h�ihl�_�A��'�+5&׷���˿�3�E����z���ӵE;УɏL��k����wKԽ��2J{�S��M��$։��D��b8�J�C�Q����[�=Xv���z���`h�*����<)����ws��;\���3ǚ��c�lʔ~*߸����!���Vp���>�ȅ���|��4k&���QnS������*MD�rh{��� c&~*Ik��Q�HJ��(8ˢj�!5@.�/H�A2�=�����4Ȫ�k�����O%:�TNMg�>)���u���x��ׁ]6�E����nK����EkO�F�)8�G<yHp�9ɷ�U���f�|ꆤ���w	L�����R�(�[4c�|�u�-�n���F��vvJ�A�� 	H�$}�)gf�K�A0,y@J�~4Q1�@�G߇�(�B؅0�*�q�S�����j�s���ŭZ����~�R��'�����0�k�Ϫ<I���AO����j��@�3�F���[�����w�!+�N����.u�/q��8�����ξ ̖k���Ki-"`�a���<����1e+�x���K�b�=}���T x���Dx}���
6 �=���q�����~��d�U>������N�R��	_����7)t^˧�yJsV�%㰦��4�0������Uu�!!u���Uc�ƌ��e �ͭ�ĺ3`�� f���r����&���m�TW{I�*��-��K#~j4�~:�.����m6�tu��jn5��~8I��=2�$;r�8��X��-����s:��cg���\G�`�������p$|�����=]�A�3��*,���{-T�#m���"�|;i4��ˌݙ��۳��֨�+���1�
�˶	����@�I%�@�;�(����]<�'{/�	
b�M@����7�@���pB[[aQ�"�h6-$8K<�D�m�J=��������d�ʮ�ɳ��`�	�=��͛�t�Un�k��Y4E7��d�Φ��E��h�Q�Tˡ�ՆON/��[��5��y#}��9 ?�SV�"C9�$������s)�k_��xព���'�S��f��۴ct\2���wڅ_��C��Bme���������yq����mRo�]�c��7��IYs�96l�����D��+�W�k�w�\��*R3_Q|� ����H��|H���J4�\a���C..s��m�څ�s���˛s�R�7�TGT����5J
Ǜ�6g��ۧ��y��Ɔ�~I�Ij@T���NI���EU�����TC���	�)� ��r�^�0y6oeJ��"��Ec	
�4Pcm��=�4�"�������ݎ���z���_�c��M�IhM�VI�O4�y9)o�>>ᙘ�sVМ�'o��Y���p<`@O~݈z��/� 7Z%�/5IӸh^&�
�d�r�Z���!!⊐� ��=�jH�@�=�v!tt�P�谹��e����R�"�����q��Qۿ2ݺjA9�*L��w;�<NC1|"E!����G�_�ɥ��)4���iq`�tsj�����	�6�L�TLY��vq��DЉ�e��g(���rm��jV�Z�9�"�p�$V�,�[ `����+�?v�Y�Ԛ�h0)U� �i�&D-���՜F�Mǜ� ��uJE�'� %y-pKOT �3���p�nեѓ�o�ˋ]��)�W���&S'���`pT8��͋1Էa��)U��9翖&�N���:�{"�(�ތ��w�_q�<9�TS�R�֏@3���[������H��?B�5N�[1����%^�QS{�|;uU�Ы��^���b�-�55-��"�#�:Tv�)�f���M�k�[�$4~�A�$�>Fei�z�rk��L��`*���x�<��={^���фwL�k�[���f��6��J9�C�	%��!	��,x~����oi8{J&�y�E0Liֹw��e����vi��4����LhP�닼ޮ�5���F�S.�Ź���qb<Yml�R@���B�J?��3m{�����xD��~�_N��.��l-��� �n���SL�����A�f�9���e�$�/�d0���Ȇ�v��q)U!��+���Y._�Ee���~����mn�=���"8�޻�=f�m��Ȍ��E!��ӊzB��nT�%���9(1pܠ�	8czv-�]�.&�ي7�um���GJ�_Pp��;��H%�U���5���)r�.�N�/C��6~i4z˻+q��:CGr�����!0+?���g�z���T�e�+1���G�����(�G݅$"��R��9/�r��[`��|�2? ��'�z�҅2AP⒓�=���v�<E��,	!�*�LF%w�C=_6�Q5��a�"H�d�ӥ"�Lӡ"�j��r�h��"kWgwJ�p�V��N�Lպ�w�����|�N=�:.�׍�v_	?�T-ws̾�V��^4>�a��|����?Ryӆi�r90ܙ8i���#�����g�'<�}�N��[��[1gds��*��co�'0)��d�a������Q)��(8)��{XeqZ=1sd�_�9�=������G�M^�7��2��0�Ŀ���f�[R�?�z�a��m��W�l�z�c��4C������k3����G�"��=2��0����[�D�X|v������<�����A���e�K�+0�:�U	��о���C�9�?�d��8��By���;��*[��'x����r%ci�J���šy�9'n\�g(U܃*�
$i���6��]7����ʗ�U�e���,��hq:��|{�)��G쎗�	�ePvK<��/�Rr�rT
�H�^XɘÚ]d��O[��Y2� �ն��)i����K"�V�7~Yz�U85u�����3m��֗�-D�5�%��y�c�����x��Y��~5�!^z_�;�S{��_���a=(v-�<S���w^�\��3~��M�[8b;��oa�%��N1C�Hr,��8���ٸ�!��2�O&`���	�.O��s���{ݍ�K�����o�YvK���Q�}�������nGw*��}d�����j��!FP 7l�@��n����K�	��c��#�y�H{�
U�*�@(���F�E9����n�%;C(�����w
��*�|�-?����@��s�H3OZ_� ��yڽǂ�Yz�����X��%A�@V�����5zX��Kq�GB׻��{Z^%�zw�Ey&���@)I��������%�[<��b�����HkA��ӎ�ܙ�e�4Z���@V ��ng<�T�ky9���G�o�<pBe���7��a��s��%nJȿ*U��ԉ��XO��J3�I�ώ�s�ႅ2��*;c_n�{@$�_�3�Z�����<�6'0�
Ú�&��p6�~̈_�?��뼋	Rߥ��g�Zʰ&�,0-����dRK�,{Q�q9�g)�t[�7�~��94�A?�'n.h�#T �;n���%㔨�ƾK�q
����]���"+:y|��N�~���$uN_�ͨM�>p��h�/���`a�8�*{a'���c��A���ut�6�։����FC�:�GK�í*�*ݧ� ��Y��,��`�=�b�:0�c�x��Ȧ�TO^ɂ�'U#�<K��>PT�H�3J�Q��!*�*;��aӣ�B���`�8e��[p�^�BW|�2+���W��ň������A��.Y��I���Dv�P��⬔^��D��F�������Z�D�1H�Hx��eI�����tl��{*X���M����]0�Ƣ���\A"b�����ҿ�V�ϓ4�R7��7\N�l!Nq.�@f��),���g}7KhC6r��X��8֡�[�n�in7z�Y�c�'`�'RC)2K9���X��U��X ̇�1��ImǕ��A�tc���l�d���!O�)�xJ�y��ہ&k�)���E���M&p��c���ꚯ<��":�M���Z����-O;6МsO$\�~	��)Y��hvA�D�� �Y���Z�s�L�3�R�R��#cjM�t�b�������\�#���L�,��/�{h���K5�q~�?F�%��$�.���W�?C��zEk�@�V��*�t��i)�NF٥Ӳ�-���7�6((H�i��&Zc^���z����Y��:�p-��!�F�FT̪�Nhrʽ@
����m�G^���C3 x=a 3�#�e�%��Ɋb��Ϣ�ٿ<1��A�B\��L���a�.�;�b���Ӣ������Ƚ��2C9�N���ܫ�48CM�/�q!�l�/���.S��fFB��<�O�����3@L�q�7�Ib�Z�bȰJ��c�݆.?G�F~x��s�VA�I���\�����srV����1k?�l~�������OJ�/Q�؍A&�^���*u #?+���y���p�U��|�T��b
v��"���
��S:�;�n:�tK�Fၨ�i���Sd��HY�/�sI�4�P8����C6=��9��M܍����颽�ȡ�V�����fϾ�*��U`�������%JI�ix$��~D�O�y񝾙�3yD*�ޏ�	��@�N��#��"pV�y=��<nm*���U5�����*R�)���'Մ�|!6D��3I���	/���J��9�l�MAR8��znU��bL���/7�?��ۤ�5pAV�1 Z���ZF�������UL���'�%�r�{
r��El@tX�Ӱ&�w�X8���1Ng�z�s����Fp=S`��<U��0�b��"[ٍ@��I`/�e1f�Q=�c-��Of���؊˴��-���S�b@��p �]7�J&�)c~���m�7�������4WuW��O���K<F�*��Z���S|;{�����KB�^����Ȩ�:�Ur+��
	\}�I�N+w���{��CS8^��F�f�����g��W�����ee��)gɝ��n�֝��h�	�b��R�!�w��C,�[�"����:��U�+���R�N����vj�l�-���!��ǆK`0`���� ��IQ�����{C#K&�;
�����C�% �ߊV0F�^��ޔX�Ț���6O�B<�u@7�Y]-QX@�<�M�cYc��xFN�� /�S�p/�����>?I���a%4����xǲ��R�ȫf��`y���&��%bQ������N��CEj��m�f����aXM�S�_f����Dnk���.T������LOy�c���-�<!NQ6~���	d��>�c��XC�#XXgL�/�#@P}���=��h�m/��O����(��/`�qKyT�ҳz�ϼč�k��D����z�뵔��٥�:/[��F�^8�j 6Gm�=9��Q�xt>�ΰM�0�Fd�	�r@?]�Cy��%��h��0#�)�� �� m4O�>�`<���Ύ�&�a�)<�`�e)6�G��47��3�N!7cn9S��Ot_eE.��@%�v�n�`A���l�̭B`�X�*r�Ƞr���^�
@��v�F�uw	kYB�V���D�ݮ׭����*�Q��,�կy������s�W4*!��Q�֫ e�b?z�O.�[�����(�9Z�@�!���c��{�:�U�7��?is3´�q�uj�}_��v���	��@���kT���d���0>�\x��%�&�'3e��n2�1m���N-�X���3	����/������ZRFvfԮ��(݉���"ś�C`��E���6^�ĈGk�%Ŗ!��y��1�>v�^���ϡ��?�ZN~qհ0�����r� �9���x;��p��uv��p��[lx>��t]c��0s^Otr�.�,_Q��[���\���$?F�f�4�����p _���H����G����,F����[%�d]�c���R<5p��! �*��G�)5Y��j ���9���ȋJ�vT���%dʤ�1�'�4��C�z��b�%��ޡ�ˮE�Kg�hX!?#��Z#|�1h�a@������mf�6t�'�y���EKC/��
;�y�c��sеx""���ǟz�t	�`�m������s}��
��x ^�㐭`�z�<&���)F��&Z���_�G�+:��e���< �9ץ��k��͏��Yf�!�.0�%c|v���@�d�Z�㖷{���m��(k�M��t��7 ��Ls����߀te�9���7�|�P� �۠kq]v!��?�#[��S��P��\E0��ֿ!G\����cro�����/�m���WE�`� h��z:��W��FG�t8�&��1�=�ܾƊ�� g�<�1�����Q�EH�0�4�f�B%?L�a� �o��$LV�����0#cs�����\0��n���~�� �E���߁�>�Y�ڂ��[
 /�c)/�.�����K9�hÌ�u[m����)��B���"���X� (ǌL��}X��=j�j��#r��}IL����؊oq���nMs���f'�Gn���S���o�b��it9
��kثE�#�\=;^ܧ*?�j��IC[8���3s �ue�/���C���pw�e���W�jD!&�\�e�B��;���?꤀��CmS�p�4�BK��4(�ԉ>�����|��UjO{E�SHXF��s��P��e���J�TQ��DU/.�H�fA���u�<��|�kk�̢T�%\����=7]�<�������kP�z�CYb�h��(]Y�\�̯̌J�
36}�[<2�!����P��t����P鱋cn(?p����Y�c4P�_����E��i�p���r�Z�ܵu�z%��3 �Å��V= ݧ�����m4�S�	�m��%e�[�4�{�mŶ��̦�� q��f�kk#��^��X��x���.I(���>?�@������D{o(5�Y.�+?�`�9�e�_�!���[�'�>��Ֆ�$a8�IT�M�n����N׼lL_����XXt]W�i?8ׇ�F���#Tp.����} �ϛ̰{��'�ڕoH�ob�@	�,�ݵ0�XQ�8f��=�ٚ�^,Q/.��Y,j����%R#n��.�.��φ�4����2��u*[y�ylƝ� �8��ᴬEO';��dܲ�1W�)Rŉ�F�:��À D��*��9���"`V����*�G�bJ��6&���7r��
xͶ���
�Q�OG��?��2�Z?C��cTeEw�6���laҐzU׵L�4�+T��!w��	;9`\2jZ��^l9{��Ǻ�-��$`�B��`�0���� `d�Ƴ�S����{ż���J����m�T:*���e��3�z��PI��yx� �:Va�$nR�D�M<�鯸1*E�\c��ϙ8�r��D�rS�'@yQu	�~��<�W��?.��Ct��P{�
����/�P��3���ۮYC#�K�y�9q���/��E8�:0��,U��F�P�8�ϯ�`��U�R�����8�����xI�2�[�ިY��74����;ʸ��-�@�۽��<��;��T���
=��G��.���愲;U�&�v�F��}�ܗT!K�#��f�.�W%�z���n�_G�[<��K��k��Es�䇔ul��6�&��7J���Y=�0f�����(����D�|�f�P���,�r�)��\f�?���#c���Oӥ<e��>if��D��}���G���uj!.���Xpn���}�K�0�4�)e!��uʦ	1�����4N���=hΊ$�Hp_���=	DKv�NG8��GdL/2] �ǭ��uh�:C�.��h�s�SF��3ٌ��M�?*��(oϞ�t�W�պ<��Iw��[�j��EWtNqj�[0�D^�2��;�N�qG��*�t��
���J�C��e vơ��S\l���2���Nᬉ��*���=�9��ǂB�>	�`�o7�r��mHIN@�D4�Tee���f�,%Ė�F>��4��L`�|6r�6����8���\g��j���DB>�)^���d��}O�NkD�$\���z#?Qph���TB�7�7*U�E������D+Df˴�#w�͸�A+^�ux WP�B	�]��m��0��%^��=t#Sdb�;��|��p�̃۾�"QRZ${�A�ua����N�pM�fc�;����dC볷�7��&B/�~.-�^��}�Y���
�搳)1��ެ��K^V��!^���;�\i釲��m��K�#W�����?���;���Q�R� ��� Yj�=J`@$y��B:b��$�Z�i��S�wC�U�`_��S�1'_Y��t�z;�B�W��g�\�h�z��byB=8����p������5A�aBsF4$��K��8�]'�Ȍ��|��?@���5F��5�5V�ghO�"�j�@��Kj;�R�m�u�0;[GcI�nm��O*O�ԏV�i��/�Ą}z�X!����}?ĭ�`��W���,C+�~ f3�C�0�(3Z�s�jS�&�Z����HU�V�h��zy
�_��EY/R�2�J\u7��n�7�h_�����
GJ�(�K�Ӹ�U���	!�?��,��ph�y�	"��oiJP�[8>�9��U٬�&���^X��b���UF��s�L�����g�d�}xj���t���a�fPGv�z�-�O>��m(�~�s
�-��i:Q�j�u��$���i�����g�DuYY���tj��Pa�(��Ĳ)�e�8{:�Ma�a�5M�ʑ�T6��WsG�����0{�4J�h�L��rk��`�4�(��k�T�Ce��%t({wN���韔������f�q�5�]%9�oV☟o$-���"�����|�2��`��^zӺ(�\D>�h+��st�Ч�u�b$ޅJ�3��s����~��yog�f�ŏ�;�v�2��޹��t�~�{��N�!�|�R�x�J�*=�8m�4��R�9K������f���'[�@�⩘6I���'Y1�9��5�%N�a��	\��F�����f�� o�w�gniwx���E*C���YN���9�Ȍ#���IDT�:Ux��^Pw�MB:JX}��/� ��u�-=����cE��l`�S�J�C!9���I�эvi�9��	]}2n�Y��՜>2�����h*�F*��E%�wh/v[��9�+���x��륔n��b��,��TpΗ	x�^�7U1�Kp�lh�!�z������6<��|,|T��&�
���2�?�*�] &�ʥ"G��T�l���j��O��d�}ʥ������Yw����*�紽�`����>�������ј�����'��/W��i���*Z<�N�����|�DuP����f'�ܾ������v��x��7�[+9+�;\wQN�S'�����9}~� ��F���㎅=�y~F��q��/M�o5�A��-P4g�WժQ1�~��Ğ�X~CS=�?���t� �XH���O���y��f�I��t���w�o�'2�������UY���W旦Y �5��@� hD��1�d�s��h��OC*��Ve/�"��&�J���dC����hs�	?q!�����l#��L��!'x��
{&��eH�g,můQ��޹���O	z�7���Ӊk5E�	/� K.�o� �V�1�_Z�s�t0����]�O��d) 󃠠{>E�^�uc .R��Fk�ρO١��rERXhl�H��)�2ªj�V�'ƿ��Q��PUSX)�+j��k$9߰�\����`����[�g�|o�Wt���w	�h>yk}:�?]\�K����IJ��e���Ar�a�[���2�ک�80gV�e7_��1�eҾ�U $)�����f��P�A>�^����8F�-3W-!8+�3C��E+�Z���g����\1��Z�h6���C���u�&"	����
�kj�Z��FN(������u�av��ڴ���DV�to2rf��}����":�5�M�����h��)~%��5(D�WI�
'S~ ��1�_Eq05�,�������y�!j��ϊHYk�T3���
5�~��9�vd��V(�kuMI���_�v��~Z~A�<��0������F&!Cq�/@�����Y'�����`A�z�� ;W�2�Ho��(u�t�BCKt	M]w�.o�����LhSjl����"�F �����Ǘ)f�TMR��6Q6$��w�g]���H˲k!�6.E�~�1�-��7�LFm^z8o��[K���;�/
�9�~�[m���_�Үs#+��>�V�o��14����bL��!�Q$���UfV9��@��*�@�*B���ڭm��,�tʈ2�* ��^(�����_���$6`1~�����8y���a�*����l�Q``a�z����/m"�HZ(&;��\��R@k� ��u~�������i�{��DI��$�p�"����aF�ƹzb�������j�rLڢ�ńH^�t����0�W�Xe�J�,�а��]�&�6p�8!SE��̙�2�4�6"�_=��+�o�z|�Q�s�č�poRfF��b}����%�9�3�����;
d� ㈠+�o�>(�e����D�Q����6�WI�T��Q��O���
�� ����H�`m2Λ64L�� ˖椾�e�2c�z�v��Dj�� ����f|�6�ؾpF��a��ߢ�Mf�L�Y�,v?Cr�I��H�pFྎV�?Q�Dc�+b��~o���þ�[Y�9O�x�����Qꩽ�w e�S/�%a�j��l\,��òJ��Ie�xҫQ��U�S��aR��ގC:��֓�r��ͽ��vs�w���k�D���M-V#���C����Q	m�o葷���d��2#R<�ᴻ�uX�ؘ�$a;j\��CW;!r�������b���0�`�m�$��Nm���RЭ��y��)��yh<F�Dif��C�7��K�4,w(�Q�d����t����f��]`�����'|�i����D+pt���v�ϝ�Q҄O�pX�z�;X�i �A���n��'�ǀ>Ш�{'��Dz��L/�S���K��2>R��$�x���I�	
��҉?Le��]�|�Y�����b�Up��gM�Ejj�A���.�m,t���D�ۓ��/$��;��N�������H�k*oq��]1���0���ڧ5��_�UtН$^���ʴs�����͓]JWn�Q���~���\S`2u�u�����"+�
�e��ft{�����18��r��Е/������@��6jZ>@���No���KW�M�8���gtJ(��xtRBUn�{��}���ktQ�!G���"���GO��KM������z�;��7���a��w�P��N�/��
������#������u�p9�"�(���_]��"�ށ]&�P�=]�'��}fǜ�{�P	��ǻ9�J��=g�z�d�H!�7�6}���ɉq�ȩ��}pw@Fs��&��k���o�	A��9_)�ĮtV�e�Z�����.�QxȀK@f��Q�%�
6����s���D�����,�,	��2*��jZ��H}Y��:7*�o�� ��%}҉��V=�7z�t]�M�o��X*3D͡�S���w���cq���*aC��\�]"?�ܫ������{*0qR�B���y��:"���v���PJ)/��ġ��Q�JS��7g����)5]}�Ph_��l�M?�dn��b�(^t�ҭo���エ����{�%�Lm\x�D��<@�}���-s���k'�1��֌[��١����^�C���Q΂�L�1)�M�d�:��X�tk��P����<�P�W�r�ҴC�r�}u3u�9,Z��S���/N�Ɇ
�m7��O�ՏQ&�:Vw��W�����.��-�#:Y�]	s�+!X3��gҺ��*�L�8��:z��3����v����®יZ-�D���mҘ߯^� � 5z�t/��W8��ggzKB.� k�9��!�h\��J��"���e�c^Pw��s����%K*F]%�s�Ϲ>��<��i�����<��6
	�=y���m�����PB����ǋG���7�*��~Y�E��
m���1M֊b�c�U���PM��潺*�z�ɬ�Shli>����)2�����!�������=ҿ���ףd#���3؊~���5$��KO;�z�)LQ�����U��)��ֳЮ|�y�u����
�O��`F��]����sC�O�}��lB��Dàv{ ��*)�]�3��pt��i:Sy�9+r!T���0�����h��ڴ0^�qct(8/'$���M���.P_n��M�=D/M]��TR]��$��V�|V�H�ÂE�"�#fU��hEv�5�x1K�K�u�~3��^�J��kU�>�*�*#K?$�&��tB'�WcU�"�}���ñ�aq0�X������;�˕��'�n�:?�JQ�L�Jߍkb��Q �9�	wYR���3��`,���pׇ&<�t ��Z��0�F}u�{�v�)�Rm(cgCA'̄�P�-��4.�Z��^��$G�)��G����S.�4��\�l���Ԩ�`^�'q��)jQwl�e�*гg�pӫ`�!$\��$���G&�G�er��q��/D�^7lN��i\c�xGo!�c����9�U_ӈ'��6��=�Q��]z`�t��X��{xm�zk�C ��ݱ�}����S�G��&��6Bx���R�퍌��R��+��E���V��D,b�`W��Pk!�A���ϡ�uޓs���^}�LѯK��Z0�@��|qm���͵^�PA-I��76�Ȥ3��&�b?���k��+�נ��U\K!Bb��jEW�=�ȇ�����,4e��������ܖ������O�޼�7�'��+nF!�[!)�H�Ё��!}YQu��_���dA�L
)��ΥV�6섷���7�
=J���� fE�K�C��qW䎳���G�q1
���b��}F�'E���͡s�ݺzg'��80��'�_���؞�����.7��_��tn	ϣ�yf�499gp:`��}�k/��p�愜ck+\��k@�����Z�:8J�~|�Œ��
lI�~IF�K8w�X�Z��У��d��I����c�%������{B��L��y��H(;����Г�T[d��~�����V������'#賩a�i�kg&�/h�Juk����������i����<Y,�u�Hn������l1P���* 9�JK!�3o�%�7�FP�'�A� ��="<u&�P�Q%���Ny�r�HF��l��k7w�bB�ㄒ+)ou@L����ރ�wʑV|p�U.�Kot֔?_���3H�[�Q�r\sO4��W�P�e���n��>�_�Dc��ʷ�"���ws���j���;�׶3�(�� �$�-2�]	~�B|�)���_���Zh�}��p�F���7��
�Ro�i��y��͹�l�
n ��?W�X>�P�I�ųV��)�h!an�E��NY�	Ӆp&���hC�YiE#��EDI�bm0�}�UI�6��|րp���6��{'��,����΃�S��z�P�e�%4��P���w	72yP����F5�(ܒ�I��a?�	C�(}mHL���@|�&qC���5�dF���a�{�z�(&��֯���S�O5�c(�V܃���
��ѸXG�"�e�="y���Z?��4����f�3;�|%w����9��OW�������5�Kc��M��"-��?�e�z�Cd�p2����ғӰ%�����f'F������
 )��>�!���MёQɧ���Ab]�;��#m%�*�J���Z��"il~9�5�gv$�t��Lk6�A-�xe���H����jg.	���I�XYP~`ũ;�����P����������
8O��
��AIq;*M���)i�i�v��X�d�"E�*U��r0$��Y1/_NA'����N6L�]�F�.�3��ŁQ2Q	ᕘh���Tv&�ꏃ�g&DB�1�sS`g;Ng�"�z���-�\	hdl�ד�s�Q�.��4��Y���~E����?'�|���>!}v&��s��@<�2)�a=�uq�{c\���2�2�pa���0�<LB}�5%\2�-H�����ӸB�����Kq�P�xܶ0��/W���LiPL�>tΜ�V��vZ�4^=I��Y�9n5\�z��������l���r���V�X��ʪP��>��P�|���.�5��ڢm�39����7��0Ot�Q"&�nd���t%E�_��_,s��i9������Jg��N1��u�8�<B|ģ� ���#�v������g�۸�a��L?J��so��+	��+����t��xÿ{֗X<�-�ȃ� �XQ������KFq<��̓�U�C5%��za=��6��
��i��6�dz*�߂�'�1��(h/�%�c*}���l����6��?�Tյ��|i�Q�gK�un #�.�Lee�1�L��s��ad�Ī.!�B
�\}���T���!E��MK�j��+y� ʳ�66���A~��ػ��xxz���$�~B=���ym�he* �"����v����(oL8,
n�cR��o��L�|����¸���,��i\<}�
ZT������c>B"01�3���jr�P9��F,E8�	S���5�`t��6�HE��;�Y۬�mi�)y�c_2ܲ/�`\�\�N.�@�f:�"a*r��|�߁�c�U$�3T���M�Mp�wU�m��42�����H��$�,�i%NH�	���%.wAP��mg�n��~a`��IW�ӌ%y�<�y��ƛ�ϼ�Ѿ��ef���x����E5�H������o�@v�te�&�r��I�(UҸT!K�����aIb-q}�(0 'Lo��DZ��b�KQ3���h|�/YEw�L{GR2BޢQ��0�E�q�%a�,G&���|=^=l*M��J�[p"��P�O�b'�ܥ]�"�Gj+.���ִ�������q̸ȩ�$���K��U=���+l�4R�8�e�/�U����A�i�1Q�y���!�=�?��1��B/��DwMw����*��_�e|`�����A]H
:%�A!��s�Wal�b����"��p�D�'aqW�y���ɉ���%*W�d���M�$Z�*E�6���}N�/\��ճ�U������Dn��nE�񹢙e),������ �x����"��u�#�gxܩ�2$��+~|K
	FP�o�2.>k�/l,�>R�l6����&K�����5����★8T�
W8z�!�"�����s�(�8}�#.����/zBqj,A)�u�.��N\�h�a��E�|-������,��'�)ե�?\��[į>yht|Gs����Βh��s������3f���|Ԫ�f�~�nX�AT�e��}���P� HJk͐5�o��*:S�pt/=AѢ]/�ݠ��^�v� -t�RP��䯡r�`�f�q�O@�_���Uz���0N±�V}x�R����\�:�[?�=���C�dB"���+'�s��ɨd@���T|�d����<�R�CȎ�2�O>J��:Xr��7�,�8�����}6���b� t@�'�z%5X�_��vm�P�q|�I�C�Zʊ��@P���"�p�պ�:�ms[��-X
c�d4ǁ��,$U~�A(7�����@p����?�&�G@���]�R��[�Bc�p� �ZQ!����ș%��R����W�ꏉw"��4��(�^�0���ܝ���6�}�_P�����6��L� �Z7$8���K��v;�_t*�p�ED
���B��w@V��M����ˠ�+�~�Il�v�����E�a�=~�X��Gb�7�V^\�K�v���V���(9�s)ZX�O����%�jD�or�F����D��q���I|I¹��qX��~y�Z뼩�ĳ��_���e%��#޲SM��	U�ξ��ĳ���-[�>N�%�>�h����j�Ԙ>�d�=g�G��6+�|��6����֥�g�HvSaX��:�uw��c-vR&�̤ao��1n�I����-���H�x �9K6�������<�N< |�����M���p����+M��NVZ<b�XLB�pu�}A��-Ͳ������k`��IĚ�����
Y	��!���J�`���i�E8�ί�Yi8Nh>������_D��bW\"���G��Ӄ�a�9�VJ�����b�1�wH��7���*��e9P["rN�Y��Y.���|�5�h3;��)������#���k���o�n_A)o.�ظ����y��fӒ�R.̴l3���޺F��6�R��(I��l�s Mkx��5�m*@������zI�.y�Ƹ��
�P%S��VI7�}#�&���c�L���H*2%��hw��	(덃��1!�uҐ�O�T���1���23��% �e��H�8u����P4�E>
�E��OΔ���/�Nf���)���19�>
�t���W0�H&\T�-�!�[��0T�'��c�Ls�����S���ݡ���{U����
�(�:�/��YY�����D�f�l ��şq^�z�}���:l�x��B�)���:���Q㭌+�@�>�d���m�$�v�Р�v��c�ʀ��B������.�tvN;�NFR����G���L3��k�Ha���Q���hn[������[������n�/{�:�Ɲ�h�P��P�^b���S}T/�dS��g�Ǳ+��N�D`[���V��t������ � j��±Y��Pp��KHVKjZ������	��L�| ��Gq��e�p�N,Phf�&�WZ�WG#�+�×��Ah4��L�L�Xr�B�)_�̣�ې�uP�A� �C��(�4��FK���!�s؄l�1��h~��j�0�R�oB �����Y��ߎ+ �p��RF�K�i����W��ur��Tc�T;uph�!�/���aV)�A�|�1`D�� ����Ixi@u��8L�P����s����lL��-�Ĵ��}[�	���VE;�(ަd�^��X|3  3]ږ.^���_��c֯�,�����lȑ�LO�XV�/^m4�:J�<�����t!�O<YOw�-�D��k����nh�m��͜>6�'�����byn:����/'0J�d]U#��F�T����[�![m�Mi��NHM���ci�D��K��Dfj�uee���K��a���] �j���,R�D�)������ ���%�̈́�E~K���gmk���ܯ�Af4�v=`��+��+���2V��(V�߂�s��/��L�7�؋���]��d)�r4;��@93�H~�H�;_�lR����zD�PBU�[s�U��As���HΊs��
�{�8���#Q�r����bht�^�`��$��(oɊ���N�Ŵ�-}����:�W@\�+n�(H�Ĝ��W���(��h[W���K�6�F�n�r�՜bJ�!���rG��沨;���w�I׫r����N�^�� "/"S��tf	E��@!<coF&��x���Y��<� �����Bh��^�L��5j�Z�b�n�<�>���0��|��.Qq�E`�ʂ
{��-�.0j�󊤛��9i��b��� X��.�
/V\*@�se�%��]y���F��L��w܌��UM�j�M-C_����.����V�gn��gjQ��ρ�w|PY���:L����2��*��v-�k.���Pd�ٍԮ���ϦbڿU����ު�R��4��뺏�	�WJ�Yx����wLA'O2������W[_�6y�����s� a����gO/�`Q^��X��ýUS@����@-�D��B9Ș��;�*}�:4�6+y�8�X�DöRR����tk��ظ&�.��_ z�h�L�P'4J�!�������@���a>���.K����{p����A�Ըv��#����r�H?�9Sȇ}�%��M,g����	����v��V�mG�lÈ�r��vu�q˵0Y�b�FM�ך�E-+gL&x�qA,	��UhS5���h��/z���Z'/*��_'�0������M'�@t�����z!��O[j��vo��P~a;,h�O�ֵ�d���B��&X�WhϾ�����.�܍qb�Ԯ�Lҡnjg],��?�4�s!m5�\E_��5�8Დ�^��o�Zh_���3w��#��+�xUc��M�ߺ�z�D�e�h��M��~�F� �x���� �m�tV�@ā��?��5���!�] a��L�W�ƞ'0b��T�g`�hY�x`�u.M�! v�����nw�2��$����L=M>�~��2�qo�HV� �#�����"W��CE�˅BJ�9v��˧==W��/k<�����:�Ҍ������M�`�_��:�=u������ܢ���3�H���5�(��u��0U�.�^���I�/D�s�5s=r���x��.��T�\���q���8�2|o��z��77E�A7�mH2�Y�x�J�v4ǐ�;�X��ZJ�9���%���ͯ��t��U:$��ٖ�V�Rf��p�MK��5+E`��<�)�F���u����U��!F&؛����{��< v������u�w�{��^�3�]l��	T�<�	�繫(^�c�z�ʿ� �+��^��Q�.1��ΚHшjkTk9K�$쵉IW�?���w]��I�sų���7�sJE$�ǧ�-���q�\6��R��][[���n�
���y��Y��yX-�jgL�ئ�a���D(7�n�B�ӤX47�D>J.��8�f��i.�'��r✊��n�ԾI�;�3�,	V�2��J*�O��B>q�}NL���yҝ|,`�=��ͩ�'�ӗ��%�IXB��2��5�j��"<ҫZ��0Xju���Qeyy_�d��{B���{�N:�Ѻ�X�s�Q����K1M[��0˂�?�������XY<D��K^|E��!�肃���^Y!6�cw�]�0�V��"*�����!������jʃ��ͭ�#�k�d�?#G�u�[U�p#U�P���	�oB(�\���6�^R��&�Q� 
={	�o#��f��0���Vq<#<�x8D5�s�\��S��.f�b�~Ge#�4�Oz����ѦEJp��ڠu!]>T��"����Qo��o�~�Hd�O�!�=I�Z�r?E��,�?-h2M�!%q戛��.a	ό�>�x��2jKb�2�Z>��f��R<�^�J%o����
'v�.u	l�\������}��L���UF�ݔ�Ũs��M_�_��ʴA���,"��'OX�X[7jT��V��=�c��J���f���m��й|��
E��˷`���7���We Ew�χ�:�>�ڑ�&n���� ��fh�����[�"�ntܬa/�_�e��w��.QXrH��Z �v�5�[X�����o����'�JZ�k�����:_�tn�<�@y�����DW��j���Zyz�FU���p��E>�A�W}lܹ��jw��l��>E��"�4As��n�8�猇�8K��#b ���r�l1���x�-4ˤ����gp��fZ!=\T���z�0w�n�$�a�?7�]�I���:U>刕:]Os=�evt��^��J�2ڹ>�Ț>}[�u� ���,Gd�n�6�b�=�ʟM���,���g�h��T���-LL�*�)���	,J��!zi�O��ԑ��b���ɵ�ܕ`R=�;!��`/�#��z�5��i	�q�ʋ;_ĩ����D�����`a~�Ug��>��t�2q�0���W��ɛHhw�߿��ʡG�}���;�9\l[���K�<?1�8Et��R)��_�Ԁ3�Y��H�h��i�e�f����T��a�0n35�S�*��:�ٱ�w4��kD]
���#p
��Q��	;MJHO�x�z
<���&ߍ�Ǖǩ_�cT%�ċ���x��ƛ��E�FJ\���ý'>��[�Ļ��½z7�PJ^'Ӽ��5��u�)��*
;�t�9��짡���z����V�`I9Q��X/W��Xv�	�9W0H��t����O64�����ի��VCB{`i�_������T��M9�.�G(�F:�MB�N�k�4�ϻa�+<uj�݉��v��@��C�v�[=�ޣ2}�����DZV�բ2��Պ�kBx�̍@��v5i��)C��0s#E��"��	s�g�?R/�^���+	􅣓�f�F�K�����p�f��N%Zs�sx)=K}�����,"����U~:X{)n6���HLaV�@1�U��T������.E�<H�s��C�p�����V-;����i��;ɟJ�S�R�rtL:�\�sXP�)B��-���0�A�w��#���_���G�5���Gѥ$����:Y~|1Q-�2�*��ME!���6���@��X�X��&L�C,��K��#v
S�`�&T}��?��H�x��]��m�v�)Jj�0�xK��f[ �Do �ߜ�j�mc�T��I/��b�놌�0�VE��X��тqGf���e����؋h$�ٮۙm����Q���t�5_�φ��ЉY�ҩ��[۰�̤�5�L�0_M�'���C1B�� �8�>�C�q��۩��!QSR@,c ��g7�z�j��Te]Q��|�e�p1�������h��4Ju���i"oD�f$2y2�w]2�x�����f1���~w)L��w��[��4��fҷt�-{����4�"�����s���M�>�P-�0��0RM�cv��,�>��*�� HdV(������eٶ�j�8 �O �8cV��PIv��8�`�?�R�m�h�hU̏Գ��=�
	���{��%.,�֞�T����5�a�\&A�@+?�Ey2�TwZ��P)�� ���|!���Oi?R$��ϴK�qZ9A
�e	�Ou�~�`�$�u9�BNS1r�8G+%�7e�ֲX1�����F
c�����#TQ<��; "x[3���7��y�Ux@u�0�uLc��c�e��2&���u�R���ô���w|��>Pk����M��H̃)�`�7�6S��9o�=|�ݴ�t���+�K����`Ř?s-~����L^���{j�0�bѕ*���%��A�E /����{3���>�,s�f!�c¢լ Q�rRb4���7o"���y��XT�_�%� �(��
�(���+����w�1��z���ed��?~�n�Į�|u����
�z��d��9=d�&�+-�L�ڻ67�tõ�Y�`���b��08�O޲��s����G��X��*��2QM	�J5"�Wb�㐤�@_
><���RJ�D|���%e8��)>�qS���v���(�%s���T8��Bx_`[�2C�<)hH��3#��4�o��� �L��H[ʅ0!uR5���y���J�&�!��1�n$�>m[T����~���_o��=r���Ʀ�>a?f��H�����sX��]�!'�B�6 ��br�K��"7Xa�dk�<-;ѩ�F���J���-�5�֭:�~n˳l�M����g��Z��&�I�6����%�r���x�"�x�)1t��V����E���q�^�i���7��if�R��%���7��ouW��hK����Br]Z8,��Y�^PG�2M�NZW?�v�+�Ѥi]���Bw����8�q*��M���Yq���e�(����L����$zJ�l����^OʜG%) Vu�C|����I$ٿ��s�����b�z�
-�H~:B�z�:Ɋ&#�@���3�5(#�O���Yڜ��V�W��j�>z�x���Pw~�R�Gؽ.�Y��~�C�io�b�8U�Wq�3u���q6 m�y8�� ��QZ<�ի^r�YAR���M�tr~���Nn7A(hT]b34
%��?1w*x]�����!��ϲ[S9]�^��#,?�ԓ?E�m��˾�W��h�"�t�ٲ;yr�#B��R�q���g�y� V��w�Q��'�⩺'�U(��ժ��a_��n�æb�Z��]�kvYd#���3#��8_B;����P���
��i�[��jZs�R��Er�!���e�\��.��ٗ��$�� oT����h���0պS�L��X�H�:����%��d�x���y��B�� ����v�٦�,BέF�B�m�L�O���rh~yJƟt4r�	|��a��Q����a��ꞧj��|b��60Z5�^v�eq�=��$�ۂ���bH%��I�<���<:;{Nml)Ap~#Q�����ۃf�ٶ�F�#�c�ɠ[��ip�����PVիxN]ŽE^��'e����=&��P��-�P��J>|��L�ϙ�:|D�����y���k����,��>u�Ä�:�/{Î�j/��.4��1��4�B�g��ҒU�v�1�����%�lڄ�_y� گN�DG�7�8a�ak�ic?��Mc�6��C������,�>OK�%60���z�I�<��[�tȥf�e���R��y��m����4T�9Be��ط/"�'� /M���wFĴ��Z�i��	���q��m(P1q�j���^<f*��ceT	Ǩuz��i�����̕X�p�$ ��My�_
��pi�B*x�k��_t��Ы��.��1΁�SU�/?B.�S~���-ߥ���K�b
���fy��'J����w�e�֒���a�e���~���Qn0�e7��c
���������	�?��&o(�����pC@f^4����p'��qQ].�d�6����R-�t�g�F�C%�����.��3���U����e�9P�b�h;!��$S��dف#$X��'9�V�D�Vc�����y�+��Mi�٭W��c�)�S
T��My)jg��;m���C���x�l7))"[�:�Ҍ�#��"Ε��ߧB�F)~<ZO���M���i�4�ÐPvG�T?X\p�';e�M�]����L�:ڣj1���q��I�m��^� 0%Y2��7 ir�J