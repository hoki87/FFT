��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#�����a�qbZ�dS��dW�����&�jӅ�Y�j=���H������]�����X��S��=��rZǳy�y9[V��9 ��B)�����8������#���ٶq�]�����"�����I��p>Fs�C��w9�A}�9�Y��.c� &���~�0y�ېSս�x��.V��<�TV{	.��/,����K�,��@���
�����Ѭ�,E�BQ��9} O⫝�D�}{����C�o;x�9n�p0u/���W�u�HqjɃ�o��X�6�7}˖A��!�ܓٿ2:��k���N�"zywB}p���2]�I< �J��,���/����c�$�)�KuNZ�Ţ4
\�8+���$'G 5&@��YH��X�|���Bt2B-�n�D$E(;�|U� ��і��A9b>�_�㹎Դz�&�kc��?`
@wO/[�
�f�@��z������G�|,R�'�d���c�,KM3���4\�1�7�ly:?yH*�D�a@��hN|vI��<(�I�8@`ԗ��g�k�����4��N{�0P'/� P�C#���?����{���}��S��x;�Z��i?���^'�׬���E!��a�����u��߂/Z����V�7v��E���|�um�[�I���}$;+�~�~l'Yp�v�#a�^��Җ�w ��}��c԰a����Y�~�:�P��[��}�$�*��h��%Ң|������t�8uJ5M����PPH��Q/�ؘ�O�0�w+Q���:���d:�XH@ՠ�0�����ޒ���	��j8 ��Չ���)b}��8���}haE�PV�*L��r���<���'2y]�D�L_��hl��8��&�/�D�[����,_A�}���e:�� [[�i{����0�ʆ�>��t���1����e���D5�<�v�I��?��M4�&w��U]øK���;���r��ӂy7���QH�twh�nk�Dޝ�Z�YwTL#=����
�~ ��3�R9�7U��N��1LS�Tw��oS�^m��B��ѐ���Z��k3G���e_2���G�h �Rt��X'�#�sR�� w��Ldn"�,�� �>H�Yn���/[�Ó�K������dwd(JᢤC�3����ӥ�}�;�W�E5����P\Mԇ�{{Eeg��x��������^��<�(R��D�����^��c�t�7\��5����g#���|�6\eg$��n����;>A�MIt���8����2vz���ƱQ�\CM�$[�Ó#D�ǃ�1��	�����- ��ׅ����<�R�FL�,��U� "��8�h^��P���U�ڽ��G]��Ew�_��7pJ�oէ��z}�D+,�["�������Ǻ(�jn'���N�$�4&}��"�q�r*��h��`��#�+����O����|�{�%2Ky��<e��ؔ�b��z���nd��Jn�c���b�˓/ �d����)k!�ފM!߱1�f��z�8t���yU	:��P,�a䗐}��!� ����@	|�_	�Ъ>n�&�/��
����hR�{��%k���
�SC���Ja᧶�(]�~ū��M����'Ǝ݉�dW�+@��D�<�Ԝ��^9��]^q0���͕u8��C�D����4r�ЖPA���_�n<ҭ�!����ho�B\�s�������b��/G����Gw��� �(���;C����͒�Q�����i��X���&�{��f3��OqG�Z�hN�ۤ�A�s�h[�(+�(!Ƣ	w¬�L*� �-!�^�
�Y ���Ї)Q�\��,��>� m�;ؿ�}�J�;Iv�F�׫Y:Ơ��+��	�d�dCB��ۭ�c�����LQ�y@�FEz�}��B@�-����s3ͪa厚�?�P̓�G��5u�',�3Cǋ�W�-�h��w�ٽ�L5~.�66�J儣{ٍZ��z�xӱ
��C̱�2gr/:�B[�����V����^��lV�Y�����)��~�i͡����ݨ`W�~/��ᓩ�Q���ۼ��x$j�Lo9��(X9�ޒi!x-�p�|�G,9�8�=	���	����2�"���\ K�[oڕ�4�{�Um~��'X- �#1�~}�Tְ��*�Ok�Jc��ލ��sa2m�\VbT�Y�Y��]^l����N�����e*��~�u�l#�Fw���'�������R��Ԭ�������Lc�ϖ��y��E��}����%YzQ���w+����i���5���@m 	�II],���X��.@ϝ!��	Y��o��L�1����_�9�ܖ�#ؼ7
�#���`(����3��63u:��RC�y�]� ( �R���"�,�Y�-BB��3v�~�ah��a��@5�r�\f�~�M+R��?��˵����߅f�{������O(��K�Up� ]Q�%+,K�'�UT���`Hȧ$Z�}����4�j�J�Bh�srb48k6�cgRrd���{,�`�6��|w��iKm�Q��V/ue�*ȝ�T�8%̪[L�y�u�V;��x��^p