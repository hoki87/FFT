��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ���������lLL�hP~d����Qi�z�;�hN��� )��.3��Dx�D\���rg���nE.z�6":���yq�O�]D��9� ���U�[��T�q<�A�����+���@�7�;#�v�P4N�b=d�@�e}���4�^����
_-�9b������}�)�Yk�P�*Ǩ;3iI��(T��ɟM�(�4� �!����$놏 W&Z�+�fpeK�""�4(�x��&1>"Ҥ�ͷ�HYkG�7ۻ��z��m��(ؽlx I�t.Z��mr?�O&Lp����G�:�B|���p��I���vi���+poY����z�����U���A��Uy�y����6l-V�?�u��Da=�H���Z��_ȸ��͝ QHކ�����P��
va !aϋA.�&(Qo,yr;��f��~��'d�h�:S�t��~hJ���R�s�}�J�Gm����JT]b���˽�[TZt�\S�����&/ Q\��+2|�6k��VE��h��y۠�S�G�}��-Z�}��W�0��	Em��I�q�5��gNtB�1|j���c׬�6\�6AG��1������ĥ��lV�Ͷ�%b�=�PbA�sh<���7���#�hg�oeE}�� ��o��H,�߶�����TǊBgݹ�R6<��8tB6���^</%�������d;e<��A��[g��7��Nߺ�B3@���(7#@���FFY.�[r�M�Y���ǿ�����JB��iy
�YT����������4@v�bh����:���_�x峦�Q���k�������>M��8د@8��� K�CY!�B5��ÁB��^@��#+Q�_��{�k���2�6�H�:�D�i�и*����/W�|���:�_Or��r�6�uے���3�U)p73�蝲��;�zܷ���Y ��%�q�>�w\����	�m ��1.������L^���5��|7�V1k��n��$���mT���wYA[{�3�is��佼��}S�`���l�����g��9��O'f2�F[�(I�5E��|V��i`}q�j���!���\� Ю�uB9��JzyR��/ �㒗/�5�.���?QDOqT�Pj������v�)��K���'R�2�˛ޑ5G�*�U�}�pCi��z�p���î`��?�K��A����\�*#�(Q7K%�/f�#@��N�|��df�v�הƭQ�`�.�냙����:��G��1%�L��kt|�L'�.�Y�@�z*'ˁ��JV�(�~p�K=z�(>�hSM�<<����"�bpe��G7*��ͳ4�0�E_*��S'"�~�.^�=��*JDzz�]3]Ԭ�Y�4������IV��n�ݼ�Ux�\:U�P��g��|��F��YG6����7w�Z�dǙz�k/œD����h� i�y:?�?�V�[��ue꛺��6i*љ�pUBW�j���Al��GW�!KRiv�x��I�sĨĝq_h7=���_D�� �:	���pH�s��#�==J���*�B-�}��xh0�j��a-?Jڍ��(\:1�#����As�m޻��Aܵ���:��xe:�5�]=o�ެ��yM�o�蔑�F���bd�U1)��w�=��Jk=1��~��[��1������DRj4m@���q",���@45�ւ(�)������I,"�Ʉ�OR���h��� ����P]X�V����Fp�T��~��1Y�1��)��4��GqbG�C��&�Ȁ,�|*\��8��
���E��+<�(�
x��5�������]
Ŏ'wu@9Nf:0z8��//T��I��ĤF�h$D����I�D���2&�jR��;\�,(,���R�I_*:��MaX�NBOi$mxSg]�0���������9��%�t+�$��ZjB!����w���]B�:h'	���i �c�Mr���z���P5�׭��feis������3ɯb�?�(L?�QY$��h0G���<�U�<=�ģ�����_u���w�s�:O�5�w��A�a�ٸ*��m���c�	���X�I���Hq�)���X��h�Ą�a���s.Q�
�L�Jj(yP�/�|������/2�9�G������̀:�-����@F�U�4?�u��F�Bl/��QAe
�j�^��I��l�&!����y,���2�U1�@,t�FR��i~j�9�����,�����o�m:˅���*�b\?�AI_����/�F�!�8;�V� D��}l�<���	"[��~w��\r9�~1^A[�?ĿP��I6Oԯm���Com�;�k(p�����h\'7���а��u���9ߥ`$;N��IY3�5���5�Α1M̟���J*0��_D���Z�a
��c5�7�)+�v���Ss��%���D~�Dag?l=m
�q�+�9���W�߳��t����"i?"����O��/��uin3u[��{���M�����Q�&@,�qU�;z*�â	����*Y2�'���lЄ%��H�d�|SAE���u�Wo����ŕV]Ni�?-��<hז�_<Y���1qC��:�r������ePM�9���;# .7t��/����<�t�D��ڽ�$�Kv�0��7[�ҷy^��Id��ѻ�6��8��Ǖ���Ƞ ���-���S8B�W�F\~T?�➧	�O�8
{^� �I?�x����g��,�눀��_d�Ȫz&��my�Ə)*�TB�tJ��p`DR��iWܳ��L�;2;ݏY��1{����A�PLD���� /�%�+ G)�d�ko���U���}����_-ʎ_���,b5/�Z��ZAh[����_�(���[�Vӷ|�7˛�u	�I=7�D1����ҥg)�3qw3jR(�<zi�l��Sf[Hdܵ��ٵ�y����Q�O�.t�o� ���e@�eʋ�4S�Ż�Z�W�Rawdl��#O�<su����b�T�������}0�H�%��&�/6�3B�v���ԐT����:Sq�	�ilcQa+:k>g珘��`��&��s0,b͸��*�V��fwZLB�K�b�:��/Yvi�w�m�F!�Yl��֍�EI.RzLſ�w�#�vC\�9W�+II��4?6:5;g��iq��zj����V� ��?TK�a����URņ��f�A���v^������,�V�x)ETAk$�?��[�J�ة������릟j�uIh�JT?ЄG�~{i�]廽TMh�2aJ%����i3��Ml�e�Q�%��?~e�IU�t�� BX��Be�T���7�Ҵ}��
$
�F�_E ����N�g���0p\j�����#����:�H�e��?jd_���Q ���r:�'�PU���Lq�A�[龉��vv-ޜ�`n���w��l������I}�T��y�$x�%����q�1�K�úܚ$�����\S�o����e�W��·�+�P�>�0��W�U(�Efܻ�[���� ��ך	�Q�g��_VcιT�Q�����MEV �I�}�H����t�b��^�DF�oH�	;z�A
�h�<�@T�&��mf�J��_T����P�+�W�Hs���������YG���<�)o��Կ���{�h�:LQ�t��v&s�f	��v�����{E	��ݟ����D?s��RD���o'x��\�e.�	e�<�?m��Zİމ���7$�3Q��cDkЄt��VG� �H�5 1��i�*ue�{.�zh�SUÑ��$��tz�,���"�H|�ѩ�8��/��^ѓʜ�G�����o7����y��w���t�3��.x�8�aA5	pı,�wƳ��*)Y"���3t"��2(��ɕEJmF$��x�'6Y���l�*�	<@�#����Lw�- 6����-?������-$��m|�·���v�t{����c�i����ZȀ�EF[��U!�b�ōN���R4��/en��Ԝa	����ż���x��#�Nʹ����*�|ť¥��y���yM�3��֍T��֞]s��.�Uh����v;�s��<%+�U���7��G�jG���Q/Nɪa�>�g0m�p��g�nn�$M��.��;7u>�t�̉U&�o+�Se��x�|�S�1a���b�q�7�aɁGԦk��)���4v��9�Y����6(��}�]��	��\��RT��BJCk�ȱf% 2b@ac�w вQ~{]���s��
�a�G~~Vp`�V���EX��iy=ܷ����L�)x�i��]Qʏ=�~yS��q�����z^E���T}�am�k_��$Q�z��+��(��4���]�OP��3�b�Zy�8��5u(�]�s�����hR}(f2	M��
����L�SLOӶ7q����. ��:&�F�%FL,��(��oQ�
�^�6~�����������NP]>Z1���Ϧa~n�w�&kSgᣒ��-oL�_��l�܉6'�G�a���W��a	��r���8��Md�,�dLNzᅽh��:���A��!��Ϧ'���;(�U�&��b�_I��
��ŴG�I���d��.��*8�"r#wdI���J&n甑�?��9.�6W�-�I>�����@$2E����nG�/��i7q�[o����+O%q&�ތ�ϓ��)\�:�|U�;�;�/)4���14W�c�f/�=� �>7�ժ"��^f�ʕ,�Z��*.s:)�e	���œ�j�)�5\�([1�At���8tTpbL�����]`�-^�4(�9�b�w���O�v2�!���r�g�1m�e/�|�?���U�,�"!�0ɖ��z�:k��X�M���c1,e{�@*1��a�d,Nx��[��jc#�,���Ƚ{d���7*eh��Oq�K�6�C�9"�T#9�b}#)v���Va����,�˥z4�C����-SX��n�F�x�� �w$8��~H��I�jx�����j��세8��Xw��9o9�����V�cW�U\��47W�B�����q$}ЬG�=���� 9}��$%��G��cf�����n������(�.����4���'�3G4!Ė��m����Lcx��h�"����~B�5�? n/��>G��4�G��Y���8]*a1�%�h���u�zY�m� ��6�����y�툝������Qh�[=�����v�>�,`˰���"Vh����`=X"�׸��x�1a[s@����,ˆ���}#f�$�YY}�+[*�vZ0��\�����ɮ��+��D�.�̱�<⟝���i���I����Y��A����m�t���fl��a�>3��ArC�;��P��!�h����SgJG��km�n�0�G���N���C��8�}>���Ea�<��UE[_�A]��Ȝ��v�_��s�dysad36g�74'�Ⅷ��R�^�_t�,��!�G�~��	 �%��2R��!D��~س,�V�	��ݺ�%������t��[oCST�yш4�����D�]����+�-#^Z�J��y�m��
0U;䇕��Rψ���Az������p�P�[k7b�Y��\��:B���#��D�Sj��x;h��Wn?�J��.2�Sd\�Ӛ���Z����_E�>x��^��R��*�¶+��������*^L�ڝe��gup�p�	��T4T�Ֆ�T����A(�����Ҳ���y����uS�#\ ޓ�R�_�{:'�h��E�O��W@��L�T�����3�bғ�.j&ܖ⧢M���_Z5��ϟ��
��r�~�*�ޅ�]B��#���O�b��7����JA��,���7pЛ�S����g���Kە��p\�!��#�QMz�M�o�T_,,雷��V	�e|ٴ��ʅ�=yЎ�$���}�t�{�>Df�t���a��?Q��
F&N�DWO��u��ˆ�O#�������(�>�ex�n�UB�����=孕p�����C��Ƅb}@�>��4�0�[�qe5S�Q9�1@OU�]+wZn�X�=/Yl�c@�a1�W6D��(�5x+:�;<�$�el��(�n�nV������j;6Z��ĕo`2���� AQ�=*[�pY��3�[�դz^��'�tXK�Ղ8��IU���k;�o�1]]A�/�Z�e��4v�޲��S�\�L>'�}+��y���e]����8��/:�Z�����W�E����h���hi.cE�W��fI`�x�k9�����_.��U�<4�2�!ⵞ"�]��r�졬�]������)�]R˱�^��Ho~K���S�������0����ӝ��=Q�B|��q\��9�$z��쵅��B�:�^�e�^�?����,��
���|�eSݱkj[��koeִi|M3����QxB%����$eeRE���ۅ�K�uwp��4�D+ �ξ�I�
��+�H�3����M�/X	k����_<]<-�ҼZ'�ח��zd�Y��ĹFg<.U�|d�"b�����v����_8U������Dͤ�\��D��f���,��v�u8�9��K�B���_�
�s$�8�ۢ�ͭ�qy8�w$�_�[�9q8^��޵��9�	@���6}�V�֕�{N�v��ib��u�0+�jp��u1[�M�Dҋ��@wk$��}0j�@ꪖQ��3�w��GD��V��S��+_�	�vҖL7'!�t����KX�N��H6�4V
a��8��j	-�����M� �ꂃcd���Ý��4X�!��@�GFXР�<W͸��ٰ��2�\&��o�+���`x���ȏҕE/��Q��	i*��)�4�6�5��s�
��>Y%���4������C��:�