��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ���������w�Ȕ�Z��z]�.�V����G�D����e��&�l�Kɞ44��WB���N"O,�A���ū����kn��($;�)�M
��a�}ަQnc3�ʵ?����2֢2l�R^g|��t�`yN}�(�B���v�̳I�ވ����*���Q��|r�y�0�$>������\[8MI�v׭����2O�܋�u<a�� ��~�	~>��J�J\�o���s���۽7lT���i4�bH�I`Q��UC�N��j(w�@�X(%/�-��6�ܖ���隳^1��&ٝ����r�����&q#�^��;�r��f1/� �@[�^�oz�`q�:� -r({e_�y8�u�Vm]�R6&.y�m0���tn�i����H�	�?����A���7�NP�t�����6}�� ;(s�E{���� j�z�E���L9&_����ǀ���d�8;V���c��x-ZSMW��)��|���IO*�Z�M3r�SG\��m�u;�p�Y���Ǳ'��%�g����O̙f����ؚ��<�	vV6 ��9}8�Z*�Pi"�k1t*�Ēr�<�@���;��-���,q��!;!̅v9H��������<m�π1��~�Ik;���� �����&+Κ&&qw�L`DC��;�Sg�{'e�ƤW<���* g�Ȼ�����`=����!��*E����s��E��&�Љ1ps�SMG��}��70Ly����#��P��Z�n� O�����>��LI������[|�j�5A�P�����Ś�Lۮڝ�w28���KP�	�X���1��?�F����a>���F�>�,n��s��B�5�*���	�0B�e� 6��ev}H���e7��g�w%��֬��!oxT��/8��)��
U]���wIש����E��*��>X�Y}�'�*�G8��x#��V̽�U�U0pJ�\?��~O�p� �PA}T���n�vZ�mp(S"� dhI��s����ʆ!C����p\���f���=�ɫ�1Ꝼ���c��	�i����f�@�u7�+ ��,���=թ2��S��Lm�F�
M©�?��IN�b���ź�҂��Q���O	�z�]�� �7
�ϳ�3�
�;2b�}��P�/�m%B��/f��@�+�Pm����%��
�![�J�O������a(���F#�1Hu3��@%��h�Z�(�8��Hvr��������4gh���j���R�11	dX6�D����_���Y=r6�{�z=���LFK�����T��q<����~n.��zW���^Ĝ��0q4.�`�r�zB>^����,9s&�o�}�H��gZ����]����MEp�Q�͂��@�J=�N���r�����#�.�֓y%þ�k��MJ��kv����k��
��������QHe�4�UBe���A�%��f���V-wL< �z��*3�C}�t�öų�g�M�Q ��rS�@��
J�IZK�|kE�]��� ���n�6sb�p��?ꍘK�kJ3"�_3��͗va�z�]�m����V\yً��+o�z�%�4'�J9�6�s�u� �.�Nt���ak[-q�@��BF�A�ѳ����uT7tXN����`�NV��e�?⼕�e�C�i�RM�OTK+���1��� d&y��\i��B|������y��h�|V�&O���]��k�~���i%��EY�Y�+ۖ݁�ۃ��nE�C�֗2�v0�\�CߐHRI5d�oS�-��,J��ٺ��wd�@��O$m�v�� 9�
^����fɡ&��b9-�)��u��9��~D
�ŮS#1ab6q�c~�'��r�SO]��60>�,_�bb��@��4�1��æ�k�.p��"	���a}����o�cp��D�Jpj�R��' �Fp�}gC�����9���܀G����M3@���|�^�6ɜ������Z�T	<���=;��F������ي ���i�P7�+fIge���Q�y	%����UH�m'�Awi螼I^�{�����dh�0��dyӤ�� b����zrlx�Ŧ�7�+�00*Z�X=�	��;ʘJ����k���K�$�(q�f(湺��/�Q��Ͱ���M��\M���b�	<ǀ���I�����?����8�5��'���kgR��n+�tb`8��_��.-E-U��^8 )
"�&�+�V��q�(�VS�y]c�-�Հ�٫�Iit�xO��	$�'$����=���c�<�Uw,�:��֚H&Mg�.9������$Z$C�)�P���� �/}B�3���u���e1nŋ`L�$4�	���e����J���K��9��9��җ"���P��մ����D_�uD0OL����e���ȸq?B^�k4*��F"��?8X��m3�o�m�����&}��5�������3�oI�N~]�Yk]9@P���?;�ڡ��\������&HuSf�_B���aB�'�v���� ��!_���w�y��ї�b�2Qg>F��F�d�4�v]������*mrk���[�tx�Ex1�'q����q�3�\7>������[�V�ng	i���F:o�E���﷛7�aT�2�H����Q�V`)^�[\� !�G�л��p�t��Toa����m�9����y!a�ϬॅQ^By^���u����6�G��i�q<�,�0l��m�c�Ul�+f������Z��Zu<Y%���!h��0���*x�����g;'�c]�^�>������ks��"��z�`�a�>)�u,�t�a�ݬ�WF�ɏ6f���%H�o�@@{ي4�f5 Q�O�t�+��4�� ׌pA@=���q{�co��2af�v�ߦ�KscNU��HϧFQ�J�����$X�Qj\/8����D7Gn�̞	�
��a*��D�'"���>����N"l�teÙ�H�mbF��3/�>p��z�_LJ�a��a*�a�DM��Ν����	K��7�6��M�2��}v఻`�����y�H����s��������Ah�n��aN�<��6��L�ZR$�HY��\�Ľ�\��lMH���x�4ڗD���_I���3����&����oO� 3�u61����