��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�#&��#�<����蒋q��x2��+���Y=�$�FxV�q݁9e�^v���U����~�����:�GG�BIF�,�r�a�BW����7�Z��z�A7Է#_L���E��a7 I�hn��.�!m
J��[���~���.�c����Yձ-w������N�C`3*CN�֍���+�K�f~�aם�eir� �jz�?��	��@&2�\��Q}<*�#� ��XG3~�`5D}�"NL�ú��-��ī���:}f��Zs�L�<>R�s;��:=9&�O�b(��M0Q]�Ө$��{�}�7�����^Sq�$U���C@���>TpG��-<�����*���	W6�������ŀ���3��I�9� b�3T�(�j��Z{k�J�<P���7���>��ۤ�<@��F0�^r(R�p(5�Pj��%�����E��[�6�;�p�\�
Q�-�6����M���C4ӳ���3rƈ>Y��E
ps�O�soA�=��4�����cʤ�j�����:��	��S7�������B6R�
��]*�Sp����	��v��@ݭ�VԱ��$K�p��G�Yc �XFr{���΀����M�Z�7P�y�ؼi�5,�6\m<��5�FD".�h�c082��\�I)�����$�V��"�t�k%�R�Or�P��.�5��ma4�c�
�H3p�ĥ�v G{�����L��`�d�u�.b�$�V1E%&�&�ݎ��<����q>O�yW��Ƒ�B3��+m5�.����p�(��m�Iw_�1��um��1�ɵ�4s��Q3���O*B�k�\�T�3��.2؞#3���u�� ��]�E��dz`	���Vt#3�ǭ�#n�C�*�8
�t�J��T-�y�	�B��J�/;��*���#��/=�d��]��6�_�d/�#��%�H����S�7m^'���9�����
��<��[W5��(F��sy�����)�/�8<'�^�3�^@��g�Y�q[���)�ݏ�h���}H�.J����iR����g<�g!��D_�8�D��h�l�/������NZ��4�ز��	vZ$�'�YD`���df�s�y�m����֧��s �,��݆v�M�_�YDlq�&�"7�yn��]i�6��ݸ��꒎@��S��6�����C�لʀ�l�ґ��_�x"��娸�/+��V��8���u��np?h �/�J"�x{�ʞ��{����=}��a�1�q_*�#��B�\X�S缹�<���P�J��>}e������� kRD��*%�O�%�m���ˆn�i�4�!��43ܿt"�/���Y;d0$��#��/�
5.�G��}D}C?ʊ�����]*�M4k��l��I�q�A�����i��!��p��S*�
�%�ڕR���6�+����H-��?P)O�=���2�sk��钡�]i#}�Զ�Oµ�u��k�Y1��m{���t������r��d萒fq�[=]?s��+��i=ĕ��ǹW�!��Q�k4�ឃ���7]}gP�0ӹEڧ��+# e#3���o��2�10SQɤ�lE���9AL��bG�)�8_AX�\$�G���`�E�9J�|��B��,I�M4��g����p�-����q1�;�G���a�e��x�{�Ѵ3I7�Y*j�1�W%f�����6��7��uJ۶w�+��1�="Nt�9!&�4��yZ#�R�c�	��qi�.����j�cÚ����^�tS�j<SD�{]��:�\j����q�w��ud��	܅����aA��/�:��T���������yc(M�<Ȋ�e�e�%Q:&����G��Ma̰�+���K^d�,�SKPU��1oQ����Z&����!�.W�h��_y��>z��?>����e�z`(���S��� ��+Mp�e�����)YA��ټ���jP����5W˒��C�&����F�7�Ae�3��!
-��A���:!k�p�
�?�u���sXQ~�}��&}�����9�D�e�\�"�z��m[0`���2?���i��pb���n�C�dtڠʘ��h�R�����>5ZQѭ���pR= �7;�w�dc�C��d���[��r���Z�:woþ�k�5U3:���Ua�xr-#�0��u��L��2@DRj��y�c4����e�=A������PC�vE'�'���,��C���	�{ؕ��8ӗ��f���%�$������aXlQ�BB�2[a�U�Q�������Z���Z���h����$��w,�"�x31�-1�mdȊ��%p�z]�6h�'��c���<��n5U�P�fY�0u��DN9��miNE��'�Aa"�����y��im�V'����F�8�YP����r�W��RmIw��х�"�R �����L�v{[p��(���@�����䧊�������V _bS��*���vH�6I�ۿ2U����G~*�����$WG^g3�
^_�UtZ5S�)�4i��������R�I\GV�BD`�Ǩ���3K���9y��o$��b��� <�4���d�zhѺ]����)����͸����ѫF�6!�HS{�<�&�ܑ�(�T�!.e`K��I��6;!(�L�'��F��]v��ܴ՚Qx
@)H����ӎ&Iӌ�y�.H��!g����ӿ�I��6��KQ�+�,v9Ν��&]���]���,}�R3�c#%�tۀ1T�#��y�
p�\��U��.տ��=��4~��6�ِn���T����;��)������8m��mOX�.�U�Yt��G�k�"8n�&�Ƞ�
��B~ ?�kH�g���W�{R�ӓ��8� E`���{뇂-�r���=x�؊X�ԑb׃�3�)�����8]/�V4i�6CPq�=� ��h�W1�
-��7t���-Ze:|�oߨ-~�����h��y�$�8%9�����]�zMBv�{�<�)X2 ������K������ϰ۽Y?)�[��]�~(�k}���. �wL-L{���GU��ȠԜ�E^�T��	�7k�d��l����Y�w>y�ߒ�0���|e��7V�f籾���F�Ⓢ������<���;�
Ak��g���H�������05�����!x��w:��a$��䳉�tY�36J���h-yU 0x�=�:��<S>�: ^��9���P��߂ |.A��T�^�E׾Ւ3�l8���p�|6��Y ���9�V�5a�ٜ
[s)6�ݐ�,�R,�O�T����/=�C�p#B���z�W�Wĥ�CΞ32Y�wp6\�Ѩhts��=f�9hI�c��ӑo!�J{%�C�28� <�q�{h�O�t\"Ws��]��%6pتpM\��W,��d���A͵**��O�	��3S��	��d���}}�^��~4�R�U��%G3?��=����l���e�RD���Nw�aA���X�V�B���ӆA�� z�vfr���o�'�+��{���g�#W���\zz��-�˹w���O6j����*�e��`�dT��XQ"��3�Äo��\�.Z?�^CЄa�$[���Ї˅�f�C�q��es�my����3B,D���LH�����|�౬�@8�p��}(?*W�N~�#a6gf[����c����"��PYZ��5e൭K�uu���Yf����Z��Nw����]?tJ ] I{���WӾ�	I(��m�*�<�w�:N0�c!p:7F��r��\����fS���&�BR؜�%�K�a-�~9'��.SU��
�Z���鑈^�Ni��f�Z��G�ť-���׵H�M{��Y��͟����J�w��ςF���`���YY=��;g�Ʋ���re�/-ܫ�f00��-E���0D��9�/�����Z�w���_Ecܭ���xa�ҔK�G�m�&䓽��"�n-�C��zFY[(����Ma�_POH�b�{�p��r9
����Օ����k�=w(����.�=��&��� J�`�VP�#���_A�S��An���ӗ��@�]�U���U�<lN-���f�A�����ب<^��eI�\Di� ��JIWҠ�E�Bp��,��{��@�b��w�c�J��e�vUD*��Ѽ9��]��b�Fa����9Ҵ�P��I��?�wc�M���1�қ�;�G.�o$�G$��Q!�P��Y��i	9%�\��c�ڬ�*�u�����gr����plH8����D����8�=LO����9�*zc�ʠ������*�:�"��w��,������Z�ZIĀ�_&�����_d�"7�d"Q�݂f�f(W�]�V�'�g���6uG��hh�#�L��d�ݻ���rBHϪ�_OS���l�m���#?��)z%ɱ�M�A�{
��$�a�g<�7�y��#��mC{Lx�A�t��h2�Ӥ��SYۋ�K��W��=u��̻Ϣs>��b4xt�v�
p5?2��*k(��%�a#�^i(�<./�0�<�r��s/�*��֋���o!�B	T�Q&�S$�	�_���V�#Ы��?�1�N ���{wd��E�{�*?���ɯ�E	N������G�Q>P��=T"�@���W*�z�g�E�����KW�ޭ�*6C��a5�"c��`��������;����`,P�Fb �z���t�'�j��?#��~�G�`�3{�������	]�m�&eP�RCnX�*�1S$N�"�ڑ[�LŹ�no���~Ab4wOﰮ��q�f��"�:.�6�D�!�ّ�Fv4� ���a,o�Z���Nn�-q�h����P�Cx���'��ٸ�n�5�0�X>1uϵZ̝F�ð�ms���� gT	�3��F��r7����E�Z��w�B���}��I�39?�?�Ur��9d���j�0xD�|�?�s"��u�����EU@�q� (��/k1T#?�DBVB�`!�)v�B|z����H쾉Cd{�7��^�5R.��&G'i�����x��?��A��#Mm�<{#~�"�˄Te��?4�drD-w��_�MLs�0�3�D��)n3�^U���[J��O{K�-��mqX�Ӂ��2�!�"�+Yx�@+KF�Cݯ�Y����W�x=�0?�!����2�oLה�^�W��)���W��=1��0���Ժre���ÔAbuKƎ�bP�a��a������x=�0��;2h���"K��2L� �ۆ����Զ.��ʜ?QW����k\��2��e"?N��;��c��z���Ǵ?�9�:F[�X������S��;�%*��c������rQ��W�yn���}�����ҩ`t�ge���Ȯ{b}H�m�"�����9+����
/�I���H0I(?{������0�������~�"�d�����՘�%�=hө�#{�:�]����o����7����Rڠ��+�����yb�DR ���D���2�y�ZJ�����Y>�O�*J��W7���������8{ŷ���Ce9�Q�%�^ff���V]���������J����%��������5�o_x���H����a�
�w�_����!�����2JL)]�CL!=Y���mm.m�G�<�:�ЦR����}_*c�1?ͤ�F�4��F�?�udJ*W���Z����dX0U3��t�!�(�Z5�!�㤈lkFI�q?���t8V'�<�&ub�@c�~�ʾ@������Hc�'�"��X�x���y!����E��Q��7d��6I�L�2�s�YA�䒍�Q�b$�Y�CB)��]�Pz�B�MM���P�28w$$�E�۴���G���W*TlH <�氜���	l��鮏��Z-[�!yΤ���j*�q�^�&��M�����.�684J���Á$��l�ɵc�
^�Yt�-45�/K˶0y{�����YP�I��}YH�R���!oho�+�_?+�AK}��?4���a)jH<M��-��lm�'&%aY:~)��3�K Ǭ�?&7 ��GW9�9��߈��̄�w�Z8w�f�<J�Vu�X�7��"���K��)B���Y���gW5�\ǆ��JpP�^��`^[.��˞��V�#k���s!\�6�I$�`���c���Y�qh�흗��J�e�������r��=!4}߮$|qF������#d�i
��{���h^�H&-�H�z-Vp��
�@Y����bV�+#��w��){A�>Ύ!�-F����ۍ)~�-T�׮��\~Ą�.�_��QP���x5S���3�9����+̽�=�����"_Fdj��g5��
6�݃�b��m��0��#�����
(�w-i{W�i�C��B�Ӄ=6z{����2U닍�r֦ۢ%�d���,��>��D�7S
-��+�n�ֽm���%Wk^�B���8���_�x=y��ʱ�1U������OJ0�"���� c��Z�x::@��=A�*c-�\'����_���(�#�;I&;.ZQ�O7��1��S!�S�Oe�/"���V��cV>WP�~ze�K����)�F��ć��n�7�tN��L�>��J�D��q�XX5��y��#��(��i�jvWu)���϶/��#HT��+�����L�m<Χ�)<�߬���m��^�dm�!eN�0�T��7�mὢ���*�n�ΘT|:�	R��ֳ1��hҁ�2gR�C�$��l�@���˭����s?�a��i�n��;�J�x>@��ŕ��┖� >�:2@ vsNH9&ӳж	�5,`٢;Bx�b��A竱���S]�~P뚋fC�"H�ud0�'�a��[\>%/e�7|�Qgj+b�)yeBY��!����rT
�ImSq\�[3��M����h�"8lR��gg@�<>#b^f�D�#ɾb;����{�oV��ՈBĤ�tͷ�h��F����8��}�|��R ���j��Ů�T���ڄ����Q��a��M١�^�1�ȱ�XحpJ� v1�!���#'2(���������i���*�o����)=�m
�.����<\��G����k6P
?�u�H/�~�oEW��_��:X9i�s�G�\���@CҖ���a�z��	I��z�V'�ttW^�9��t�+n.������IPqN���5��#�lz��v�Q���m-���*�蓘�@n����rA��n�����͇ �%[?�m̊�ѹ�) M��n�k�f�t������}���C�F;�Ӧu�#�y� pԅ+FaN�\���>UF��z�vz���9u�j���t��'NP/FR��0��b��������G��fO��x��QW��?,��pV_�$�B`�粍�2֜a�wQ���j����vE�&/�9������{ü:a4t����Π񽫗�a�^E���&�`n�7>7^TT�K-QYnߩ�4"OG(�kk� |�M��ƀ�B�$��1\�~��~	+�]�F=	V�kX�7��N�v������˓C8���a�.!Z�t����ݚ�O��DfC[ѦF��m>|���?�C��HU}wR��G��^����``84H�vQ�hA �:B��}�(�=�*bC�E����8W��~d����x��ZXa���2K��>�g���kT�?��|A�G>�6����?�G\�e�N�pF������G�{7�g�.@��B��͋��o4B_'hթѨ�ͱ=;�݊,$�Ι�	;e�R�i"a*�fi�)�MSp}���1-fJ�bU���9m��"ﯡ�ŝ�ZMy�MB�)�#��4���ʀ�qMbsM��z ���{g� (�=�P&�:�Hr���� �a�E�fG��� N+���f��1�>�%*y��(�L�G��ަ��*/����S؈t������~p�k���Fk���H�p���۟��Ljк�95�]t��CN�/����P�c�[7��Z���UX�\���7#��O�P�&�������<����^"�o��F*rNբ�6�qS^6�s�P��ڼѽ^�$�)P��t1��}�Gc�����,������ˤ�tq2�\r��ȍ��c�9��+)	b#]��Q6�G!G�ʧ�l4{hf!,~tU����9��� yJ��@��>��q
DKL$��ExJ��A?�WD�E߶��ޅ��9%uޭ��+�=��͛V��m��u�Tm9F�IY� ����_��F���k��d�������c2�}���u3���q�^p�۟隇�ŀ2%�X���!K�D|?as8�$�������W�H�@�_��V�$K����9�o�?�5������L�[�����g�Y�^�~:K�L�G��k�'���\��+>������KA��)*�g���K�0��F'���*��saE���DѨ��a�7a(�bQ/H�wp5T��Lg�H�Zz�9������7�pd�|�N)�N{%h�y�6�,�j-2����#Tٙݞ��Vp��k�6��e�xt�'��C$E#�����o2AAe�� p�#'�As�r�>=�d;�Z{����{ '�a/�),e$(�;�� ��N�����-��evL�I�;Z�4���)4��}���d�@�J̋6g̑�����U��)�005���a��^�(^����ku���H2����w�`oA"���`w͒����J��d���1B8/H��H���ǃ OKrʛ�h�~��:�q\t�u�"y���8��N�C�����D�{���ͮ�B[�u����]��v�`���7J���a=�֔��r���	���c����S��ZFg�P����*����Z�|*Χ�屌=��Z���JuÁ��^Q��/�{��x�����W�p��.�'/�g2�x�Y���c�nI'�7pްd^��;������ �(a������l�@4k�		e�0��.�8�ڿkȊADͣ�%W�Aړ�/��Pb�@�)�@��5v��s%��sϲ���-�?���'�K����,���.(qvWgu@�J�O��nd��	��� 8pp�7����Y��`\�)��7��q"Wrt7>_�UuՉ��e�����l���R�a}���u'��� �V*�P�q|��-P�������T���٭p:����dc��� ��Myqd(lX��|�M�B�P��*%h۳�����9b%�n��i2�j^_O�֌)�^:�Hd������Z�笺)X������*eq���zߥ�c�6"(<��>�G�0s:�Rԩ��/�RX��+�xs�S���F�YyNz��-I3�-���P[]�ʪk*b��.����̦����s���:e{.rB Ntb'��si��(�y��@�u5�S���:
S2y��C�P<Wj�Zi����xA�ga���W/�/�ٷ����dY���u� ��H��8 +�N�-ekŊ^��2/q$��������G�6BJ��_�)��-�r���V��Y���E$��	�n�M�4�W�@���3y1ږ���M'���H�_�?�͎
Y�}��	�.e��2�`� ���J�r���F�0���,�l~o �I���d����l���\�����K��>vK���NeR�ϭ8��cpq� �8C}�m��V�{�Lw\7���Jin/@�Mrj`F �h��&+u��QZ�x�)�P1��6����Y
F�hY��3*K\٢ҙ㤶��x�"��rU8]����yVo;MHbZ�[��׏\$��4��)`��y��O��1��Yh|y�y��t���W���&{28���W�iȽr9ۨ�\M#b�G�?%@zLԪp$X����������,75� b�(�H=,�W�uVh6f�q���̜�BS�@�����Km����2�8l)���s\,�?1z����IWt-2�7	� �3���*��Dba��L��S�q���ˉ΄U�w2Љt�SkmЗI�U/�.$�iL��ZR�6�s�Dc�����A�����{"}i߳��"�p��ѣ%�I��=m�#^�wx�
���r�;�AC$<�H
|�z3W&AC�Ӻ��{A��h�š��|����s]U�+���=!��jOH��(o����S�h�,�e��֣�	T:ݺ*���{��my�v,��������Ѥ����!�΂������A�-!��55��F������Vn?���M8�X8d��F݊a��Y��u]�{fve�}���qĉ��81��UK5���|gx��'w�1���:탊!jiJ���Vdԇսz��M�,��a�y%gF�n�����w�s����4	,Ā.Dډ�?�
��R�kJun^��-����s��MtwZ
P��i������8�IY �rΘ�p�B1� �P,��Sw��j;A辶`j�7U��9ۿ���\n�>�j���W�2�ksQU�O��[��:i��t��R��eB
s�zq�ψ�P�QKV� ��-b�0�8c畚`c5Ӕ����3������C�IGn�j�������=�w1�i�*�����x�cTL?���_q�[�EÄ�	�ʢ��&E�O �<>�i@������cUt
���qL��3�#}{#쥥&`ތ�tn���g3񒴔�K�N-�u?��;�wu�����:�f��?!�Ϭ�5߸���n
R��۬�}�3�&�Şn���dó��ݶ;OJd2[���!�`m����T�gkʬ��"w%Vo�Qcp����� ��S�&�/�t�@�$ә�CHlF��^t��=^rS�M�&���
��O.H����>�v9��ԇ����O�"--'�Q�������	���RG������X�TWꃐ����A8��y����s�����w��K�PC�J�����F��c��!�XE`��ie�Ф絎�����zb|�V�5�����_QGg��R�xې����r^%�wy-�o�O��ШW�B�&:��ρ����ɃD����<h��a��y'�ޚ:�6Q��ZI_��0���[� �⻮Y:o�d0�?<�D��q���/$�������6����E�[p]�����XQ�QKֵ�[�����Ru*>ua��Ff+"
��;C��p�p����E�+͡s|�X�s@N���q_����s�i�d��.��y�%{��Z���P{��yd�=�:{����G��+�N����� �Jrd%��r`V�1����p�Ԅ��m��*��4�x��NcΚ�����[O���#�߶5��ؽ��N�AzW�L$��(5fm�oX��lU��WR��!]z*3�j�k��S�(F��0��h�����{���N,#4��ސ��ze�������t�_���&���\�'���N�r_/�R��5��T�B>i�峉D�˶����P�{��sR�H ��8���5Z��伎��zc��ˊ?�)!%w��ӳl�=#��lݒ5T@#���fE.�mD@z�I�BF��'U��S��4�Do\��g1�{V���/�(p#,5+ 2cۃ��x3x�3�^�?����n:�`OΣU�űU���s���������<�qg�������*�'�#��l��61#��Y+�����5��Ot}�A���F~z= m���i�����mRI��UL��^pK��7A�:��Br��뽛lcO�*,v�L����S���w��Jh+J5�G�<K��&Y����0�Jƫ��m6���C�K/�/]�H��R)�������8����e����D��$�T�1l\ߋ~]'U�Q�.C�
��B��U	OrV1�짱�]�<��H�e縁'�W�:<Wd��^�=m0���_�yn�ơ�r�p�Ѣ�ݓ�SxƲU�|�t��Un�g�1�I`����պ�͏C�G_Z*����j%���:n�1��'�q���/\=�R��	pr=����n���=S�y:ZaN�%/�"!P!��Mq�K�"�P9��n����I.�#����a�	��7�ͮ��������Z��ЍؚEܵ��E ��=a F����Jn�b���s�E��7原�'	gJQ9͑w��;pP�,����^[��ѿ�u=T���|Hw��.9^2*}�P0k�[{{�-���ʣ�bfؓ��f2�L�p���̬5y������20<-jHc�J�=� Ir;��H�<�)��wzQ	�P���8CO�#CA���c0����0�e�FDټ Chs��F�_p�=�3^�ʟ\��I�@����_�:◖I�*g�� R�xϙ��?���g-[����%����;�I��Y�pE�}�\_���Eq�*���mz�,z�S�e�ē��k�f�?�Z�v>P<�.�	�3���y�땆��
K��th�FS�:)��[���d2b�
�����������
Y�^*��f�yc�cs�h؜d%h���5���h�L�RiO�E�g�V�c5�Ǻ&��:���&O�5�E�����nJ�'�.�fV�=Nc�S�z�_ =���h�}�f��M�)"�c����t�or�dd]�%:Ѯ�F�h��tN�eew������r�-�UǑ���/���ĥ�Ih7l���tl�~$�eƫ�x ���5�@�-���7�ͣC��S�T���u��])�.�FcIO��k��m
ZD?y[nَ��I��%6�ܑͻ!�|
��j"����S� W��vUT!��)�N:U�*$Ӽf��{0#�.�JA�toO:M�ȕ�YRo�,��-�׻U*/.0����t��Ѹfʬ�	"�X��b"HX�-ZهV��a(G����9��9�����X�	}.���_���A&cf\g'-X��3w�61�bC����(P��IcjB�9>����0�C�@p�Q�w����'���Cѐ��T��L7�w��8��j�V���1�c��� v�n�t�I�`F�Cg�c��"���#����>~�ڻP$��=m'a��f�ʓ��)ZGX��bވp8U����(���&�p6�q.:*�k���A$~�ގ�uZ��j7�����?d��~��0�
���$`���	CvG#8M:�׋ഡ�S�s|ಁ�ƀ|/�a79q!���Ra���K�p�c�h���X���?`<8t��J ���K>V��î�9����]Fz�X(�z������<���	�z}�
-
���W��	���[\��{�X �QD(��o�2VkuL��)D��.f'�P�jm�|���1�SS?��q�aB��蓹��H��c|����W4� L���/���^�I�^���K��̼,5a*+#7������q�P8(�N�q���a-�����h9����R�Xfs��cv��>��c�����8�41z�K2h�h�!�R�""3ʕ�QŔ>t��ԙ-�i�#+��W��хKo�Њ�4�hA���j���Nj���E��+Z���{���cZ "��4���i�W�{����mY�q5�5�ʄ�2) !��x�]8{��j�,W^#���yl�d�ZWX.�|�R��ԓ��;c*6����J(f�pQ������z9Q��!]�j�lm�C�%�#�0��z�0�]��NMp�T^5�����e͙��0����m�|�6قSc�r������fLN�d𐃣�^���9F���"C�}�oS��֬��q]-*�I��}�asM���aT�"�<����ŻA�l��I��:����ȃ�6�1rOx�f��	�_v�pmNdZ2�{8�(���%��PK����wsUk_�=��L���3��Zºic�Y�P�&������	�������i%�5����ځ[��L�`�)Z���
�:䚍�;(9%��v#�xfVJbG����|��U}L�1����:��� E>��1{/Q�����Q-�Z�����ޚJQ��.������݋��=�?���y<P���M�l��5L&��X�)C{!݃��t��)�xo�G������(����O?�QE)%H&:�3�iS2��� �R��=u6���&�����@<��6)M5ۓ5�׳���5�V��o���T�-� ��r!�� �G?Ѭ�� ����?�i�ؗ������V%Y�b���}.GM�Œc����m��&q�i7��W��A�-�:��:RQy����hC�"K��ڱ�q�zQ�#��|!���w�̀a�g6���]-�1�Uu�ǚ�~E�9��`VQ���P��N83��٣�����B����B���^NN�0��'zag���d�=(#"Bt��H��;گߦ��P�`l��
(�������tl3>��k��7W �Z2���vYka[�/
m�\���b�IhXNњ#�O���k\\V5�V�Y�4$EB��2�J[t)��M�0/�%��E1�H�4 ���:�ot�?�Δ���
�-.K��̰�[���!8gbYK�j`&��+C6�L^��X���B[�_��o5�W�&��G����X��r7��հl<Y�3M3�*2���f0�şA������ӹ��?��e[�2�F���-�Ђ�r��B%�!��S�O-����7�{2eN>(�Lg��x����Q�6�/94��i*4��AU�1^uW������?�Ha�C�)Q%7y��'F�-]Lg�� 388�L�ǃvN�2����8��\ٟs\ԩbK�'�'ޡq���*�2��Y�+�zr�9��:�����-��Ǎ%X�B��7���^��J���י42�fzg:tg,�hE({R����,�%��35�F��-������������i7
����Ҥ� X*%�|4y�M���$s0H'�Ŭ$�4���މ�_|��.e���I�?�k(����P�-Ƒ�0��;0�/`C"Ё�(�: �^�����񧒡��v�]���5qGbP� xPfJ-bD�O���1��������)Q���"���A�A���몊)�@4�q��N�`D�^z~gĮ�2a_`�ج#���_?����r���q=v�Ykl����8���C�)�g����W<��Z�,	X�:��`1IM�uWm���D|�8u�s	����9����<vF�d(f�`6���T�Iw}�W�z֪i�@�E�� ���'�R�>c��B�����4���to�4;�|ʎ��� >��\&_��J��$W\ޞZN���������TD��!���L�`V�5��q� V�w<w�xe'zm{��^Ð��3t��[`|d��.߯��*�� 4�Lv81��|hۻ��� E 6��w��i���E���v��ۖb�m�U�qym`E��s�KQ�,G��D�Ê�_V$�@Y�ߥ8��}H�R�6[�k,�Tr��ßN�;..:��XA�d�n�ǮWoO������J/��<{SB�ģOo��m;;�h�H�S�ZW��ء�X��"�9}Z�x����9XrʧU�S���춞�e����/�F�`,܁G��LH$a}ā�WV���_w$������=Iz��H"}�h�{8��j��J�ȕ�{��� ����/9o<В�):g�I���ӹA�HT (��jR\��Lx�	F5htTۦ��_5�뿾��y�9E����t`5l<jٗ^h:��Ɖ5˛_�Z��-����c���o�$�7�W�	KD���Hv�Nc���\Vʿ8�[��1�0��E&a,?��D�/� �Z�_���Nr�k����5:e�ͩ�Q�B!@y�����$����?l�uA_�qH�"��#���2�=�nћ�c��N���D(���xt��$���WW�/���;yb�O_�AN7��0�H��r�C=k%���/���,�%���Z� �Π�ɿ��g[JTH�<��ߦD0Z�2�����)�d�Ԓ�,���d4��Xߔ\�`x�ݐE:g���vī(QI|�S*c�Lf�(����4Gt7�_���<R�(�Vq6r*��b����,ǞH8�7���Jc=L'Cy�!��ܑ��c�����F�l&�ظ�4���Aj���ᗱS����`竀�åy����q�����&Ոާ�0�L�e*,p}f�|g���N���U"�Hb�Zڪ����U��U��a��Mdi � ������(�ky�� ���m��Y���^��;�#aR߱$�����Z0�����X�5p���Q��:(��>Lve� �7v�97��R�6d�#Q�Z�
_ʨ}t�D�~Y�EN_���(�y�Ř�k��l�����%_��Zjj��n:�)R7��Uф����?�q�?L��9�c�'>��NQs�&�s5-���,=}!�zT
~n��g���W�=�=�@q:�;���~G_̆�P;&H��P���	� O�G�ݭ�}�j��<حEoo��Q	��{�냠+�w0°�œ��\�	-3��3ĕY�6���AZ�
��99I�(�-鑆��5����qu����u�6PBb?H�O5#�����;T5�=�l?�eQ�M�����hH�@W�D[~��O�oB_KaN�@�>����n�%!r��]>�FϪe>�f���w��Х�4F8<Y#��[�����y�v�	�?g=u0L�J�Z�"8#cr�90o�7��{Jo�Am�7j�P?=��M+���Ԁf슜�X����>�Ŀ̓���~Ѡh�,���z[N�KP�R�7)S�`E$v��ġN�2c^�ЗY�]�`疒K���bpLm��>2S�M2�^9]�&�KJ���p$�頵nս�~g�����0'!�v���9N}
��д�,?�=l���L4�5\��8���V_��e�.Ѭ�i���uj"�7�̔c��:qD)$�Y�V�w�8�+bI��Ը��Ѣ%�v�[�C|
R�Ls3 dI�
@݅A6��,�a�B� b����0;[�qj���y5A1�V�+�Z.�{2�2�u���!n ��Q�c�G6,��M�#3&�]��j�f���o��2m%�X<�rK���_���Q�����%x?�WPlu&
X�ʲO\�՜�ۼf$<��a�7٘�!�Jt���3gB�׹�.3HͿ��d��X�Ǎ��p�q��t������Jo-��$}�|��̿g���"�ycc��a9�ᒊ�曤������`�mt�8�7�̻N���-6�@�n��e����yd{y{�9�*��AĠԩ�lV�᪭boU]5�<� 6:Q睊h+��M �t��N�uS������7P��s.����;(�5lkW�������*C�7�u�b�� ������t1�P��z҈s�������L������(o4T���X�v�;%�Δ��kZ��!/q�8�fQ��b�Ӭ���bB�]�c���ʄ?,Y�&��R������YI6i�%�� �bn/�2��`s���iKh���t����h���X��&�y�n8�`Õ�I�-d����_$Sxkb؀Np��Ϛ<=&4�����칽��w$9�����`Ti�ɐ�)U�Kd���)8Yp�ߏ{������npmD\*�Zeۺ��M�*?��7�4�a����f���Y��$�Q��\j)1�0��Ȅ27���W)���Yd(v�p���{S�č��l��j܋�/��\��g��R!g` {��}㔸�R☰�(��iX���kj	�G�TϬG,��5�:=ݑ59�N{�q���(c�et��)��1�L��Cx	Ns�U�ڸ�e��ct4�>e�s*-��rt1�$�	s��`��؍�����7ĆR5|�gd(���i
!�Nc����>qWyț��B75F���{<d"���,h~xv:�	�����Ǩ�ղ�c5�-9������\��N-�_p�Lo���,���
��O��q�[�TM�V�
jK��[��-�4&C�}Y���Ґb�1&3��m�[C��}S`��"t�R�:��3I�(?�.A�E]V׵�M�igD�6�hƌs0��m����bXP��u��`��.�%&یu��8*�,�8���GV2QB�?��[^����=���`pA�Q�N|=��I�)r�U� �Bݱ��˵'r����y��{���|_��b��zt�4�W<�zc���S��P��ђ��j�Uj��)ǚ���b;�a<�w�ǣ����c/��K�C��ױ�"��6�����9YK�����\1�֔��߭Y@́؁�gNg�������r��2�j|0C�g�h�b����1[��!^�ַ��ͣ����%'�+ɑ�*�S��-��ۦU56�?z��hG;����mw�i0�sە]FN����	L!=	�',��t+��z{�x�r'9��:[:mO�~e�B̰�FDh��n?��<�]̘mᦔKkl:Z����ס�$9.��2�_vK�d�BC�L@�HvF��ٹ"iގ�R
�O�:+�*��r�����<��Q����?����8�6ߥO��'�2b�s%�]o3Fc���pq�:H�J�|FH?�-!�"x��zC��KF��&��p!�oK\i����(�	����I5$l %)���nN�T���p~�GZԢ3AҲ��i/�܃R��[���|����H���@P1K�WڈN��f��`���Q'Qb�J�	ߵ����1�o�-?m!��� |fdAf�<&p�ƍ��m��\����Ya��N#�\@�I`Ě��+W��ߨ�yFbԊ����_�v��ۥX]"���8s0��~_�i�ȼ`�\�@�bX�+Y�����v-�!]�% ���-�2N)��),�f\W2{2p�\������Y��k��}�2KRHgpL����="��b���I<�"2���Sy��.�E���^U#�F�|���'7��-�N��4�)Я�י^Qc�e'97��r�4I���ZmW�������B����A��GQ?@�/�(��� �R�Q�����Y+�'�c�A�P�P�GCB��ʧ�j�D��<�Q�����잸Z����1�q�h����w����2zO<���"�����ɇ�!��`�Eq����R��Q�R�џ7`A��_�\I<��TDl��D�;�f� �H(�+z�_����^��a��uw���Q�����V&�X���9�5��.:�Qtt�a�ߨBbq!I��͐�Y��:1k��N�7��"+��`)h_�
(,���Mu��-Y2f��x�ׂ۝�+���E?z�h��@�ȶ�^N���`�c��sWl�^��q��M���ݞ}S+0����qaq�R�&��؀�7�"��5�����j�]d�}���7N��=�l愝����&v �X���[<���qF�{���Β��` N�R�P��fTS
����x� ��<á|	� D�q(�)5��^0��s̏\N�  �v����D\�`=�}�^�f�mՂN_��P��B���̭�9B�'s��/�$X ��<y�16(�,��L��D����Z�l��X�庑4Օ�P �+�H�H�QM�H�K��jn��sJ�H�Z� ��z]+:˰��uu쇢J��H��E�@dR�BCB���o�䥼_p��?�R��~j�y~G�爞�k�?���F����@��/\:RM���,U��EP��Q��5PZ���c�.@���L}�X�����i� �TC��sX��~���f1/R�8����#}vӶ��m~9I�_z�q�4��컴q�K���z�T�8���s�o�A1�X��mJo�[!5����'bom�c�����}!l�C
m�k�����2g���l�!�����_���HM]	�x�6��(���;���7��o�R�@d�A�	?��� ?��w\YX�74��>8�l^�<t���$��'�,u7j�٣qM��cR�����#U�Οg[<�\|F�c�1���m�`ԑ2Ҥ�4��*���� ��ٸkZM���g�G=�:��ԅמy�WH�t��.�t��5[t$�j��2������ܪ��88�$"f��xE[�+�Y�����P0������ރ�s+�ы�G��I:v�w������Fx㟅
��n5^Ie��W����������n�&ؒ�t52E�'��ͤ����B2�$gfR�'���K˴Q�M�	=�R��[�6O��A��KFN�Tے����E�́�o���iW�s�)���i2�p���DK(�hvD;҇Բ����ID�2��gt4���cޝEž�9�N�-6����H�̲Ώ�Xt�Tn:Bz-��` �\�b��?�"��^�~��2�2ȷ�t����Ӊ΍"j"P]7���N��5��}]4�Tv��D�h-u���Z�̕�c�jk�[�-���A��kz�jm��ѡ6�o���[e�ᧆE�rU Cv��/�*r$���2���� �%��h�L�bb���3�n����!������Y�+���X5��[����D������c�*0	��f��O6�	�ł�o�/x\�?�4�B`�K���i9���:Q��>p��E�}G�#L���Θ����반�ڒ|P��5t�û�N�V͏G�:6X������������9�>'you���\�JbP��quc{�d�_D�	Yy��^>�f�BB6O��8���_W���&(�%M�Dj�R�\E������iR�r�_�d	��E�Z{1nZP5�1��[�[�8�GVt��p:t���䈵ʒ��X��)Eqzt�:�[��p'h���*���=�3x��O}[��cMVڊS��� �G < ����tr��rs�v�p��>��$��r��)ZŇ�s�cT�z٫e���˾���d�� �BA�-#��b�]��1Zt���ⱄ'x��P�HL�XzSLS�M��E�9����p�٬�J�&�*����7�!<��,�	=䳌j��vG�)���P��[�a�AS��W�"��0��2�� ؂�6׹���F,�=�ؓA��;�o��)Fl�5��H&ڞ�+�V5�,�laO�Փ�Ù^i�wk�o�J�q71��7�~������b��6V�m�MJ�L���a�F���X\������r�p��D���aUs`���G���&#�y��ʚ���!�
���6ߵ"���ţPG�.BOmGCI����y�}/B�;˂�^��hq��NZ���.��p��Ϩ�*$��|'�;ɻ�#��ݎ�h[ Z��ԙ9���& ����'��5�;���Oċ@��6=�7��������Wl9��ɦ���}�/:���$[�N�!��52�+m�#�ҧD��q*9��>�KX������.�瘁f�ņ�Mǫ�n�!2���"0hw�J�}H �o�F� �r� }#�����v��1��RU���Q�di��A�@�K!�F��L��UT 	)�I�M��p��I��S6#���b�\����闄���I��*%���KG�Epq^���v�y9�d��[�����u��#B�4��B�^%����d ���Z�k�26�JSX��݇W�Þ�e���u��1�,���2�Ρ�9�N�ɕY�ͅGE��g�_Z�n��B1������nyxP8n��I[�,�vк�(-�[�5%/��w7@s�+�2@�iX�c��E���1[D��^�o��r;�\����t�=�n8��.��N��Ԅ�ɻ��EgU�]����R��8]��HM��28����uғ�F�W�a͘)���-��j��~�cug{f�Zz��V"���Š�(,c��ݨ��?��P�bM���Y/�@8���J�O�(�p�����8={��"�~FWKXxA�w 7���z�T�ʋ x1YӇ�R%N��N����;p�Z�L�J�{K푸���/�2J�!FV<[*���!�;�C]���JaWi��E�L�-�Hf��RAM( �����\$�j��Q?�؋�@l�҈��Β�2��� (��~*��M��ϕ� �?�2�{��4�Qx+^��V�y��%t<,�5o<<�#{|��)�@R�w���H��񑮻�սEt�Q��֏қ�{�&{�������l�:;����b:!0L�b���,��e�O�����	_ࡰ������c���@}��������lS��X1@Q�W~����](�	���0���E�;"��֊��Z���?<(ȳ��V�"�DP���T �rq��|(R��.h��%g�Xҙ�T��9�:RɧҚ��w`�������L��?}��PFgw�O���`��<�\vg�P�p�]]TF�w{����=�ι=p��b�)=yu��@HJ�׋_9�Y�*�!>�U�߱�3o��j�����s�`�ۧk�W���$����[��g, �����o�Q�{z�v��Ĉ��,�b�"�!eo��#��{��WS� Ԗ3�h����b>ʖ�@
�u��)ʺۤ��3JL=o@�������)=$vG�t�9��C��\�$9�p�q�OX� Q��l7�(n��-���!Β����3��T�3�!ЗN��#�5��δ*Ndj݅�b�DP��U[��	����PmE�!��Q�Kӥ�������H��&���� �ι��$}�E��1��i���� G�����ts��32>��e�_vo"K͘�V�Jt��	M�m!��7a
��BZ���׮S'l��F��}b�M�K��q��|%���|><V1���+UgoY�U�.<B؜�'_�T�H�����`sz��T��
��&"�b�{�s�����P�=(��"��6�����_����6��?&6�۵HO��:3��Z�V�#���'n�����XI���o�*��|E)bs��d�w�S�b����i�{��=�5���Ԑ�~�A{�3��Y[�������͖uyQ���	��_Ӛ��'���am;��A���X��ׇ��3�Nt7��.�Ҹvƹ�k�-	m�qtОQ/@d*T%+�h"�D��q�غ�o�RZ�e4 �|��x�*� �ϖ74q��6���o�z������c�2�/�'��$����0 �7����)�8%��H�$��gQ���r�QE�&h�����R�*t�n��!��h�1���J�_D � C|q���s=��Q,�w���댢Iħ°X�U���X���:e�(�k��eL%Kohxh�o"x^��d��vT?e@�������=����u�s��I?��H�1@���	�i&�^�р:4W��} :1bd�@�A���v��f�R���hAdg!0����1�YL9�;b)l^|a.i�e����^�p���Knq��ǎ-,2�( ��r�қVu��#��W��^�����T:G� LI2���V����/���!R���	��
-�K!����$.�Z���z�o�Dz�%)��&;�|.�/t��'���Ϥ~SZ#��^"��`!إ(������b���(�;e��У1��8�$���j9k$+ I����-�&\M�JA�\�I��zj�U���hdc�t�b��ܧ��FG����^���2�JF�Ck��2���y{	�:��D�OEt���X9��\�u���yk��Aj�0k$R�i���O$��P�C���4���b���.�$:� �&�Y��S�~O'��(���T`�$/���,0�-	�u>EE�^�&�[�2kI��~>*�i@��v�]&i���i�,qF|*�5���N����Y%���u�٩Vt��0�T�a���8y-���˚�vRIŒ�{����N	0Mf"Ђ�MR�FL���Kt5�(��}EW�jǕH��̏��Y��-�j>�s�k�A�	�� ��6PJ#Qq���D�Y/ڥ�*�`�a����]������0И�!�ɟ�+�D�KP��8�%�u
i��Y��Y��AY��AZ;tH��הh�#1���S�T~�8�9<�t���zJO K:;�/�Jx<F��rP�1K/t��Vx��[�s:2�ڞ�u�������
�¶J�N�Rk\��u 5�i��4��HU����0`�j�?�����dT�@� a����������0��NW7��er<���5�o}0�|�#�X���0��@BQ��5L�A�����u�y���O�8��ε�qbF}�/C���F�۝�p� 8�#*1�4MX�)��z[CU�rahڽ!��Tb����& j�85�P�vd�$�T&�e&k$�*Uɯ���;��l�Ѳ��������m�y
�[���,|�K�yGGa� <#�k���ȸ�	�^|����nX���,*��h|Dy8���8.�"����9�8�%A[w~!P��b±�v����O@�L�֯d���6,�8&/X�g�t���Y��ħ�c���{=1tm-�pO��	X��o��fxL(X��(&�{<���G!�,`���;��w���@K�@��ȵ!�ޅՐ��<�q��η���^%C����
�W�Y�}����l_��>w��Lt��T8�`*��`����,�e�.�d)��������Ǉ{q{f�� 	]!��-�wE[Z|�NY1v�t�~��AI�L&���M�#j�	-�q3Wx@�#�F2���mO�;=#0�ڹ���ǯkS��3��oX�zy�A��
6eZ���;�ޙJ_�@7,ԓ�iC�v���f�۞P(>���	��d��Nv�A������0��
>|n�^й��Yg�b(kS�U��1��W:n�ҹ�SԌ����R���.�=k��B��C�(;Q?V��.��ؙ$�*�y�R�?6^$5mz��寘�m�����/,K�Q�hI3}��"�hAd٠����g4�����,���G�L7���g)7�*�(;�/|�l'���}���I4C�q�5e�	I���J�r�h%��Ps��Oo���KD�k�=3�᭓��\S������Vw�&�v𕗦���^X�`DY~o�:���,����\�-M��~�a�����R�_�:hf�QAZ8?�L1K_-Nb�&B���Ө���~�ڟݘh�]
@�^eI|(��$�K��z�����hq�F��
�uf�sI�,�(y�wrۍ!�e�,���B��=3�h]#�u(�:s�f�E���H���Z���Z�w��\xN| ��K�����j�t6�;lT��m�4��!���7z_��S���,D�ђx���m���Ms�	s	ٮ�v����I�Q�5AͶ������+dW�m�DWkk.s����� �P�#E���5����Xd�/XqR�۴��%g�W�Ԏf�τ|��'d�b�i/����װ�-M;m�vӯ�l���#��n��sj�&�g4wW���f :�s��r����s9��O�� �dʕ��
�j�@���%���=�<��nţ� .N}����p��&�H:��,%X��hNG�AM?:�����M�,��v�;���z�NJ<SP��̧���n�?�Y�`�i��� +��M��%mr�*�Ҭ�����,u�5H'`μ�W����ߝ�����~���ӕx�y[R��Ր�xy��XJ����tɠ���%��U���RbU�;3^�w,E�7��Xn��'?�R���H�ʉ6az%\(�Y�hE�\���0a����h�q��ɜ�h�&��:��s��R� ���b4�O=����gxv��|p�Y��y��/��߄��G�U����9�Q#���N-hTW�{cq�ê�R��J���? ����Q��+��Q@������8bh��U���*� �q���ўQq��l�H��ٛ��>[���� � �:�xrJb�p�«E�(
�<0Z�W2T��GQ�h�+����/DB8�4N�H��6����{5����Џd+��m�����oؚ\���|����#؇´����T=�E���uq)Ϩ�Ѽ��&�&U�|�2�CS�=n�: '>cK�����r��7��Vf;Jw�d����t�H&��!�h����w�4�֐Y�ZԶ��y��i���	x���ݩz�������WA���V#Η-��)����	��I1��MJ��{|��03	�q