��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ���Úx:��_F51��H�s@�ek�>վ�N�h�%���up+@{�`�+D3C��?>;Lm�hco �$̭h��
�ڔ���X��t�h<��S�{��5nǇ�o�p���]\6-�-4�����>S��x�Y�2�z���{m1b��#A�:����d���	�%���ό��P�m���+2���*������?=�&���hJ�|��
�p�:��޾�*���b�1x&ʒ׭��@-!��f�r�>gx۽��y����]r�o�Q?�Nx�bF[-;@ �NL=+�B>�.	�"߇�߸
)(�h�wk��k�w��K���kD ίl�[ys�@�@�ʍSp�/np&�~��Y�!&������D:Zh�.�s���z�0�CD�s�h�:�x�2�1&7�ZCt�n�
ǞAL�<'�]� �g'�5�N��<"|!ij޻r-�n���N�@���Q@��@_�aלv��2�|x���_x"�k,E蛩�lk��P�>O^/<q�D���oA/ǩ��a^����Ժ�T��x��vy��
݁�e��D��3�LB�'\�XW$����h`8t��-��:#��-�R,}�2v���M6�;�I���Ŗ�!k�Q�o�!Y�<�jmE�[i0es(����K�i�6��=��7.�P�'WZ`��g%C�b{�������U`��%IZ��F��_D�_�zB]j("��t���� ����ʯ�tS��/S-@��~B���Z�B(�!�IP��5姪�Κ�Rw �Fn7��8��.O[!!��:%D4 K��2��J�	����!�(��7F^�E7�;��KB���6��e���L �]�;��+���M�!��s/d�jSv_��Of�ش3�;җ�{`����P���^�A*<x�m!owyG�4d���gjm�}�}��0u��L��N����V,5������y��Y�n���Ӏ�H.qC�����ǵ3'�bϩn<���P'�w|(G�(O<@��'��� �oQ�4�p���W����*��·E�_bX���F{�-�+��z	���O/��l�@Y;����aE���"�EN�y*
�8�aX�i�( .>�1�8��D@�ξ(��%k��IQݴŰf=BME	�R�+��E�xJ�%Ե@U.O	ᕮ��٣u�!;zL�G���^L~]Af��j%F8�6f�6h�A���Nv�e��+��o_ڐyK|�����t��]_i�u�^Y����o�LE���~��vBr�KĊ�r.=��t����I��J�����P�ֹw�϶����R��w�ek����6$�H���@���J���{{�6.
�3ӟ��)9���j9�10D��~�^+6����R��C��k#��-�,�z�mc�9v$bq��1f�I����;�y���}���q�jXҪ�4pUU��4������V[�4!B��C�y�;��C�r�W��uM�}�
Fu|�β_7������t;9�\��s����������:^��^���\ձ�i�k�e�%f�ng�Yr�G�Tw�����x�;i� 7j�`X-1(<=�D�0b���9�V�/������yj��?�aMt��ْ���0ĝvؼƎP��J��-<xݺϜ�n���E����xQy�G�v�0�N��-�ko�J�@�]���`�����{���ճZ�s��1�'�F\���||T?g��f8�
�w�cl�8��85P��	|-$�����-
fPT��Cs�rHz�Ȭ��ܝ�����lS۩&�U>���(�-V��/ZO����v�+wU��]K���-0o�|�;���:��b�\v�h4~C��߇#u<�˂�1�u�(��]�n/(�bW���,�{
�cup`SM=����$�s0���|������\��Rg�e�^\���q������	0�h@�w�g�S���BҺ?��~��V��]8�Ah�YD��"(�ن ��wgRG��y�i���"|i+t>o�N�'g9�}��~ ��CS��l��z���z��L���sS(��p��Z��FR�G���?�[�
5��Ӂ��&���)��w�g��Z�'v`f�#�Q���l�!�{�6i���^�9"}�'�I�\ڱ��L��D¶���X3���Cu��`$i��8�2�;��]C����+nb��rb�l�� ܪ���ۄL����E1���1O��-@���)Y~�o�5؀NsC*���f�)s\I�F2E!2e�tE��Њ���Н]b͡�����t"8���>����d_���*�����)"��ˈ��ޚʮ-�U(~R�-���2���?������DS�Ք�LF_��2��>֐\�푣T�SA�)�����&̈H�$ m�[_��#yM�;�
�?�;'fG�v�qh����D?����>&�l%w���ѴP�	ak3p��9>��2��N�S��\#{p��q����-�d���A�u%�}���:�B	�F�����yFG`������+,8L�νԷ�V��c�eᒛt����)�U�	�_����#ժ��@��nN��Hˮ˚v���A=̵~@�w���� �C��#(i�U�c�X��7�	���-X�\�X3?+m��-�~�g�FxB1s.���g��l�A妧~e�����/�c[{,��eջ�䄙��F�c��p�9_����%F(�	�%fk��ή0޷+;��60��3�HG��N�O<؅�����o]�5�D��S��Z�2�9U(��r�< 
4�I���ؐӭg��g�q�L�Ѡ6utW��@�M���`�ee�G4�V^}Iְ�BM���az��	���-}�Z�la˹����-�8c����ټ�ߖu�jczYIr�T�~�g���R0u���|���7�S	%#�\�T�H����a�b��ƍ����aZ��8S�����?_4�]��/���AiZ�J2�r�ތnjǱW�A�j3��Ee�>�\�y�k��
)r�)��J��>��EX��n$Y}>ަPH�7*��M|�A�8����k���7H����V=u�=�J��dai�^%L�P�X�zs�|���_&;�k��!�z�Aa}�)�%)Qi}C u�6�O<���;��B��򯨲���}���-u�?�§������	��"�N�����c�26�7dQ��M!�}צ�	,��� @}l�ԃ=����0VjJ\�엕a�E��Җ�shn1�jB�Lg��i?B���&!�KY������� ����Ћ'�
�͢��D�P�������ͺh��xYm��iq��	o�N��R�f'-`�`��x% ;Ax6���׆���0;�,I�����jա�d]�8��w�ކA�[ІTq3���*֚dZ ^x��ӭRC��=�� �xY0�=h����":rK��c��w��@�����V�ѹ��wL�$!�ek-�y���#�l~?�]R�d����ԲDbn��x�j�.@4��G!�<��@�P�Y]�*/f�C����ek��qr{bչ��%4��ڮ��񢇚�*=O7�I߈!&'vzz��-OD�B�Fb�D����YI��h*�SV�S��� A��c��+�N�)��Lט�9o��Y�3�����$�g���C�no�d�PbK�'�`��;�Z�1��xi�\��xl@e4b�׻�X��|��S���,	e����q����4���Ċ*-�5%�v�wX���B���ax���D�U����Bm�"�+�IFѦ�Z�v�u"n��o�=8U;H#����)�����Vݾ�9��ȿ�)���ϨI�r.��n+k0��~p/�E^@��G�c��E��R�۬�[O8���>��y�i{h�`;\��=zC����QQ��K�h@�Q��e_1��E����W�2s�O&u�Ż��/��~Ϸ�����+D�jv��\ ���ԫ�y���h�Pƶ��w�qz۱�f���[�R��(�
��>t�i�hqs��G��FhBy�����rd���KA.�R���kL;�$ߝ	��������<5�u<d��ϫ��D�:v5��b4�tT3n�� ������X�x$�c?bd����ptg�&�'T� {�f�O�J�C��E�h��6+_!�4���v*mTu۩�;;d�x�)ڹKE����d��߉��� �D@��Щ�*�4q��X��ѐ�W<��z��Q] o%8�O��e��{\(y�0�l�� �ܣ�TF$�˃�fR'����y^"֌�fq��m�x2D;�9�cs�w!���q��-����gˠQ��k} 8ayNŘ�q�o=O�̜�*�p{j{������r�m����)�WP��-�@V �ZgZ��<g}��p�?rV�b�f��i��]/+�4#�%Ƅ�Y�f!��_��:O������#_�켉B��6������^G��g���n.����қ��U��\�m� Qv5��J�C%q���n��<,����8���Q��[h�t
�+��'*mj�鴶nw�����HN�	,�Oo�f�����&`d��	�-���x���!L�J��/,���ƍt� F�`ݽD{�դ�V�}ƀ"�Ygo�K�=�'poH�S��[@e�6Nq�[͕y�y��������>��N �����\����6zu��vAKd�2Z��Z�*��1�
�6�78VYt�w��D�HwW+h4GO§�=�2��� R����%�P!񵘋�?�6��%����;�7})zҸ��E���+ NP*}�!�`��GB�(�����߹`C/���ȼ(��� m%')O(�J�@�e4:_..Oܿ� ^�J����)���AB��k�Yô4F�69-y��(	��R��w��xw<��wj�AF@�L�J4[�X�9���sWK��&�^����+��(Т�Irv�c3��59K�J>|a�w�����~����,x.F��Z� ���4$���j�~ʸ4�ƈ�V;���{�}�"���q�����޼�O�X��f�|�sH�le���)�uz%/:��P���y�x�I[�8��GH�,��{��NEА~��>�JK>z�\o��P�4EL�^يf�����j�8��%1㟽���t����q��G������*nL�xk��^Z��#=���R��� %rp��cl����:�Y�z:B��wi���`/���A��L�r=B��?��:o�8�iw�8̅����������A�3/\]4��sd#��q����0	����E��i=���VR�렇�⹆�o��(��؋��j��R������y�i�4���_a/����`�1g_PFIë���}$)��H|YaO�� |\d,��k�J�L�QJO#�W�<b��
4���J�Q;.�6�uߕ�}�gm������e��6\��S¢
tsP �|�?��م25�~�N��d��� LfX����k"�4��@���,��/T�Eֆ
��30c�f�vu�Ux;��Scr�o3ErZ�ktl��
��l��a}#���dGL�+��l�b��G��>��4��*�^���q�!% ,|�QW!�ް�)�e:�|�뵇൞C�b� oz]7�M�mYHJ����,L��Nݸ�?������r�f!F.�a9�����1X��/��p��"�M�^
�9�n/~�	��qy�2�2SOO�y��wׇ���o`j��Y$�_g�%֙ms��;m��κnw�~6<gao�����5v>�Q��6�°�K�e{t(��{ u ͫ��Va68a 㔌,$Nl�������97���ЌH5�<��ъ�x�_s��\Aa�B��͕�8��e��=/_' |"s� x]�+X�$Q&��R�9gl�0��?[�9��RQ��Sab��O�'����8�r�U#�V9���`��˵F;A(��hSkP�B��el���^��߼CP��O�&3z�?��f�ҾHc.5��S&�/����t�����f��߬��/���:ei�����u+�Oep ��>\��M���P}yL����"���ϊ�9�f�[X4�ݒ�(Og���(Ue|�x�*���*���@]��dy�?�U�Wp��kd��DiR[uN"��M����:��o��X��xh,��\ k?^��YZ���4-����b���:��7P'����K��+͊(�.Z�ǯ`B9~��7$�6EH_�.;��2m����S��x�����%"��,GBgE�MJ�ʾ&�u�$|����c}+��|P�:������գ��f2!�*2�1��[<����	J�
��i�i�N��r�d�]vĭ����%��Q����۴�@��X!�`h�=��i���&�cӖC��8��%�y[e*2_�{fn ���4�����B'Porف5ڰ|<8�Alt��&x3�/R����K�E���?��~,c*ٌ��x���_�?z���K�&��C��G�O��՚0�U-�+Y��tǒ�˦O��|ɫLb����qfV �~�]����bp���ǅt�u�����-2����k� ����8|������M?K~F> �s�v��/��`��l������gu��!��(ڤZ�lĚ�H4`��5�7����dX_1�2���S�ϖ=�����^^��.��X.~�&M/���F�B�c�<EHVLkG>W?�B�PW�D1
K��_�G>b�"w�|��5}T�I�!��k$��hf/*�AuU����O�5	�k��L7�ө.��%�oߴ�F(I�9�Y�z�(�7s�S����o��cówyg�?�Y^J���'�-GWB����Xz~kzJ
���B�J��� �2�"�,�����,I��W�5r�����av�-��q���#�"#�:OmY)�l%e�[���<��\p'-�ߛ�Χo�6~�b��ޱ}���^��6$~]z��3ԱX��mVkbM����r�*�|P�ō$��ۙ���"銐=k�}�X������I�=E�N�y���\,j�{���Y�$���ٟ��کJ#�4���|^2�����BF�\9*s��yP�R�8���NV���0���J�%�:��w�'�P)��j�p8�{�|\�;����ƌQNnkz�p\��}9��xM��>��:����U���}I@'͢�����3B�5��j-�.�� 'ʪ��6<��F�[Xh�u/���r �c���Hzx���V[౵Lg��/M1�q���m}���V��������o�=rz��6�t,�6�Ԕ�u�b�vʺ^�l8��2��u D��М����툋G
��f1���_v���y/V�C��S�:����V}d�83��vpD(�?�i�{H�[U�y�~�)�=,ؙ	���s+$\9HL`��8��70 jye�I�Y^j�����N� p��ƚ�K�س��N��%���B�jp�����H�~��ǡ����Oc�bV=���D-�4�r�иӧfD��W1=f�#+�7M�W�{�[�w��a����M��r	��> g�Ϩ��o�`b3���YCc"0��CA�Ǣ:)�1�b��YyKf�0*㫂�V�mc#'[�SȺ���@&N;�`!F(K���ZS���nd���93X�}1&S���R���s��o{*":<g��!�lG��3���=	tK*N;��Y�׮-�K%B�����vu�+��0G0�Wi*eR�mzBT���e��]��7:�/m�Q<?-;��hIՍz�	Ə�������뢟%�0����n����2�Xj<j�N����\����7��mA}�9#>��UP8{&i+��3#	*Wlw�K�)L��ظ$�����N68�.�.^��5�ab��e�O�s�1�����_�֛�x;W�%O/���ښ�����1������@��޽��V���J�D��IꝹ��G���U�~ �Dj)<l��>Ɋ�aU���)<���s��H���e9��&/�b��5�>}/�6�o;�&CNH�vs\Eݩ��K�y�R%�g#�QGb�<�a/#u5�=�贮�{4�Ɠ���J�����H�,�e�'����	f.�;��l�e4�^��d�<	�'��N�k��]t!�$�f@=e���º3�6	�P'�:`f�Z����L�����D�C���ƾ[�`�^&� ]�ɜi��=��D�����s�J������b7�e�_4�g�*����ݫjj\ZG�� @!/��)y�r����"��<�k2���+��&���x��jmg�@̙�,��p�ߤ��F���9!��D��cFfi��T
i�]4��" ����l	���]�$��j�S指ð�CS6��yX9�FL��FW�&�ʶŲ�A�
`N�i������)fJk�<5���,��8��z�Hk��BG��r��#��3�hC@��半�˔><;��[L\T�q�MA<&9Հ�\��#�&'�������'bd�R�o�b��7��&�W��O�i��lc��x�7��n��P֭��eΛ�mf�<<�K����]��*�'��4o��ʒ����Q\�%�Jњ����f���!��őn�¼i�t��h-�Ld;�\�Qh���9�`w�J���*�$�/�b�F-0�u6f���1�Z�Bѯ��Å3a�Ĳ�,��c�P%��I�mz��{y�P�=�(':��j):��2z H��8v�aԬ��C@��Mrݒ.j�]*:Y�)w�>|�d����H�#t.q#ۼ�M��4h�4E��(0��z�H�)� �D#��f6����W�҆�&E&�����������&`d(��#�J�6�U�~P�gВ��R��A&ܑO%��;���W[S�Z�Jc��"�;g�X�iD�޲�W�C���:����	��p+�D=�k�����w�*���ye���k�� |���{�"�����oz$�t=�N4��{m����ۥ.�=��ϫ, ^���!kￄln�QC���!hlI�e�w��ζ� AK�ݼ���N��qҷ���E�KG6��Jk5�Ω���q�	�*�A=8���1�4���ڰnw@��u<�"�e](�Z���tv_�~)K����j(�h��J���ধOt;�h(!ʨ��X?�\��5�-�?u/�SА��Z�f���.��:킭f 3��P���������S�}����7LY��Cr�g�Sq��B����o?;��U;z�$��_C�!�ς��5Rŉ���NhX�6!F�6x:��,&�:�U2��ވ'B�R<%K�����`q���YK��z�~�w�J��D�j����}J�_�;�6��<&��5:P�{D�d�(Xn�搗�}�`e�KKV�S���x����4SNj��WUY|��_'}�E�Q�y��m�'KJ��l��6�h&���P���gU�W21L�3)���l>|ije�|Rjˮ.z�����(���5����Ƕ�7w���ax�_�����g�+S��r��:�@Bv�E3�"T�&`l�5��z����B*���Ǣ�f蹻�χ��%|v��^i$�7Y�S�dS"t��0��I ��P�ϙE�z��D�b�'m��ڬ��g�t�2y�]\�aX|��ck�f<ėJ�I���uid��m�&J�����|[�S�i��	"�/��FR׎񾲂 �͇J[qf������wJȝjrr����=7�	"H����=�a��_�L6T�-P܈� ��^�%+�o\��?�~�33aQ������~t&����y�]{���Z�@�h}��˩镅b۠�	YĠJaK�����ˏx��jWL�����VWo	���T=��@	[�2|�P�����t��2Xw��X�\�X��Pʩ����e_�2��Nf5o��[d[�#d3���6��+>#�����}�E{/$�&ɉ�\)N�F0ZƂ��V�+�Z Z����+��(����/�E�*���3�Ct���I3�4�o�꿖4ܴ�p����]U��|Ӕ��v2rD=WT!��MJ�vow;�Ef�L�]��p!÷^�܍�e�_��A��q���X�%Mp`���Gc�2���9E��*C* ���jw�A��Ԍ��>�'�|"f(=����������p�SOشm�KH���|��^�i/�1`�� A���Dt�TVrz�#�P�2H� ���r�=F5Z>��M�$5.-��R���8����`�ɣc@������:;ٝz��8
`R��U:�@�v�ܗ'�P8<��iv~[���})�kr]1E��f�>uIL�ш5�h��"�;.�c_�)�XB��P�j����<����%=QMk�8O �z�t�����_k�`�ܺQ�H4��ը܁#���w�b6�y��.�J���w#^���J����2������4�����u��`���L�쨻xWH� ���3�T�|[t��-rr��2��U�7ڲNv�<�\ZlY� � ��U��tXu��V�1�U�c�︄?�*�D�u�bFJp���4/�{+�ivp'ز��|�e�$�D�;�w�O��%��`x�Q��?��^�/�B����PQ��|�ij�ళ+�Ϟ�=@�Ez�]t}��}]Lv��J��Zru
+n9�2&��������d,i���s�=l�/�*�T�.�,g��2��h�������u���к!�{jC*״��$�lBzΔ�{�Gr�����a�9��>:j�,%^)�q�䂹��������f^@6F�?4-�̷�IV��������j�Y�+R��$fTڦ����ݳ�����cp?%��2�	�Ӭ�a
a��w��rD�3闞Q'����?!��V�.��F
�"�#����=YSYv��ǎ;�'��������NQ�$ ���#�D�8m�"4oō�Vw���5���~~*n�z�����Q�+>��4+ś�]Q{(2��Ӥ-��B�U,h&{ąeO@}u��X�A�s�鋑���X8��p��k�o�b��P@YF2wQ�3�����y]�2��?�?�$�0��?�4�^���F�mY8ے�2�q)%�	�<f�nw�Joaa�o�~������c������A���$>&� P�M�:��іF�kZ$��$�ۆ�J�RS��&O,4�M@�>�D��gK�� �W�9�Qꊤ�9X�l����-�|�]糈���:��]�H�����Y���'�C\YLhh��5�Ffx��&Zh�Y���k��-�<��lז���v0p�X�L��$c҉�G��r Z�P�L��[�,֒ɩ<k�eZ������F�N�:�}~<��;R�����	���- ��=��u9�w
 �>�5�-\�2�x�*F�;J�0UPEu:����q|]H�2��z}ψ��h��KMS������h�͛�~x-&�'�!��'&6N��x�a,L\!���t�.�Fۏ�x<O��]T�6nB�8�a�~U-��!�SL������ʒv�<a>��l~0�;���p���������#y�Ě�rQg�����hU�T����� 1@��AQ5�Վ*F��}*xڿ����˭�Έ���:Sx;��|ʖ��I?Pk�����.mܗ��JԴ��!����@N��n�,2���w�����o�
Z�T9;BCs���a�0a�7��u��{��j~ ���H��`-@��J�f�:� C�i1��g��?��X�͏p��Gy�n*�6�E���(�GV��Y�����r:��:��Ga�Y˅7?1`7U�<��tĢZ�}C|��&�*�,ѩq܉$~1�S��@���cÆom�߬�B/�Zu7�E!��飤�S8�	4?a���[�݀�}�R&������hu��3�� 3^�R�����Us9
6�N!��V�ՊB���_H5�M��.1�2ݮ�8�C�D��2����co���y��:V�2�ߥRu��1�,���%7�0D���u���M�Y$��Ǳ׽���J� 9�7x�*0HF&�5	L��A�|Tk�ư�u�)�[���9E�I�����+4@A��Q_�F�(��2>.�����i�z��1�/%�t�vQe�E��D|��ZVQr�J:.ξVJ&=����x�؜�.jTxzMb'�]��g���_������-�
^�� ��!�I�G��y�}jL�2t�lˢ"5t/qXE�}k�1Yi�e����B�6��i��=��i�A~NvD��O����i$���sᄁ��H�z�2�?ٷz?v��~��
�޷b�"��\Ga����Z+�4�9��$͒o���Bt��4�rs�!���XI��珩�7�ܞ}0MU�,���@�JϏ�·���|@R�+ùK���VH y�Z{_���|cY��&Q��M���%$3祎C�ȁ�苓�񖌇n\���dCخ �I �&	�(�\�b�ץ�Y�.�d)�~�v�\�:N�	6r$��\��:���Z��>1F,^�`FT��T��f�U�tR	�$� ���Ǘ��$fY&�;�`��L%�\Ǩ;�������Y�4Eճn��3�&<�OV�A��Ml���; ~���幰ࣕw�Kd��wv�����t����)�R���a=��gc6��!s���)�b\�4���/0b����rD�}�1Ҝ`Ͳ:Hac��O5F�F����E��l�R�XP���aQ*�w�j��m=����$���C��L9�:�^�[6���1�.�?��ac��W)s�p�pd��WT�n߰0�}�+���2t��Kޚ莎�I�Z갓���Z�$��K��P��x�~��d���0r|���D��y$�l�B3x���
{F�4|J�*�
�oО�q\'s�\�^��W�s�3 r���nU�� ē�0R�#&���1;�OH|��'�������d�� S�U�d�H�!N(MPT����&�ޠ7>�z��+>DlT衤g!9���e+i��M�Eiz��n(�ݨ�弽�����_2~��>_���ۭL�l779�Ĩ��s�/�W(�}u����cn+��z���Iw�����;�Bӽ�� �J]���r[�o���lf)l���1�JԳL�_T��V�����W�{��b�2�a�xQ"�,�Z�0�4��E3VRTX�RC!I�c����W�\M*�7�xW�-�1Ȧ>1�1��� ������K�c����'���󲼚�Y�[��R�V|7�E9��f���eG�c��	��:Y�Bypl�ߑ�Xhn�)���R���������;f��/t/������<͇M]{�����L�G�s��OE�j�}�>��C+�^�"X�a �KH�p�L�c� �ƍM�쯅pk�D(��U�S$��gp��G.����So��O8������v�w��@.�=��nBJ�Hm:-vz���ظE{||��qu�:x*���ᩢ�w�'9�WtoܙvL��l	W��0�y�~�I1*9�pGK�=���T�b��ýv;���*Opqx%śE��� ^��PN��'�X�J��vJҟ��}2�Ʃ뙯������������ނ������dJ���X�0}�,�}-�^(h.��Û�	HQwѻ�O�#-���Z���e�c��d(I(\�Ӎ���݌��v<Ƃ3;�f�mV���:["��1&]�|q�o)��ܿT��2z�����81;&�S2�J��4���ej�nesQ�� '\�� T��юm�x�ݽeq=<$������H7�����[
M�_��n�tW�%�4�J���,�(�K�9\6)�ms�#S���
?�X�a��u5�!~�\�����^W��-ie9*Y��uJ�v;�̹k�Z�^b�����?���T��r�ko�}���c��1�������^����s�(76�P�&C�N�0|���Hs�� ��({�,�9v��7�q�\�����Ŵ0P_5�+5��2�a
%fL�s϶X���&e�w`��9{��>u���h��ݥ�z�i�7�hӔd�?��]e��B����Y�8D���u�V$�����F�M@�.�Qa_K;��;���n�yd��E0�� m�Ő�.a�)����Ly3pz��oڞk,�N=�(���2˂d�n��kJ�c�2�>�*ܺd�5~78.�����:��J�X����^T�i���Z�T�(��Yj@�QZ�8x�'�"�.�%��B�5�s8��(�u{_?�Òaw�-1@(��ôF�MM#*����Ք�>����F <�~�Q�ؠ��0����љ���&=O3����ꆟ���X����ѝq~T���Za�&��ҧ�d��6[�x�.u�� ��P��ג��5���V�]���D�|�?J�h�yН
��P�B���P�{�A.�mԃ�<�W��p��s!ݯ�t�uт]��l�P��u
�����1��[��xY�]#-��p��͡�W`#zsa��.bG�8�����EH�hL7l=���ET��[�g��?�"&'�g��$[��{ܕ�s�4R�Ҫ���J]��Ҏ��8E�@�(?a���?�QV �^[E��}�cTOk:Z~��u�-_�I#�r���8h�A׌���r��k��Ӌ�;/Y��?4��U�Ŝ��m��hR}g�D"_	����{<�ǩx!G�d�9�h`�!
����r�\�L
����q�Qa$ڡ�
��F��	�C.�!�*	�4�m�)�.��m�X�73�mĹ���`@aKZΑ�����z���x�a+������A��Q����al=a���Fn�H��pVg)㭝�D�j�^)�_��_/U����(�a�}F8�#4�Kp��r�>����/f�;����}k)f[�x4���!����XU�s��l���b���X�
��5UN��Z�N�k���bu6���^3����S0Fh��YѮ@T]���ԋ��I�f{��(� � .�|L l��<�8�H_�O}T���C _�7�3B��cLcTgs� �m
.��!������w�F����-ж���r�2���k��H���-��c�dy4�������޸�o�3�%ޓ!�y�f�;UMf�ns�L��I��=Ϟb���A^�>�ۀm8.C�R	Q4w�T�4���x�@r�A���xG�y��>J�C�/���=b������m�o�-}$��l�A���r"-(G9	�qi�вq���T��?Z4#�w\������=��������zq���puK����MO��V��7GJ,d�#'o�!��e�"��^.�������� �_G�)���6|6��n�
���3��@v�4�fT���\��!@2ő�W���K���E�}�V#�86��͟lꌘlt�AXb&T��4`XP��}:^Q0���\��P/^�/E�j��?ni��<ڶ�8^�����Y�>�C�S#���u�����;,+a��0R�c�~Oc�)'�	X��~J?��UԺ��Jd���W�C��U<�v��y�c'�!�l�����|6��8���\9>A�JW~{�H2�6�tm&��9�����͗��҂�zE_7�؈b	i66�׌��w�!~ �kl����BSIצk�wtkh���#�!�,B�
�t�
��?��>��=1$%#OCuG����m�p1�d����Z@;�n`E�>u��@��gT��ܯ����S�щL����dDL�o1*����+_ͧ|"K��jJ�3����w��)��v��'��W��xX��O�۩������u��XsBX��5���װ:hb��0�ao�t�$
�,�1�2�i�ȳ@�Sy���g�Ԏ�jBA)�
8��j�[._���2f2I����3�+]F����oVE��r�Ywu
y���`=\���IP&�	��Hb�敔�i89O� �����ǣ%�� �Y����'YWR�#4�}�dѠ�+c!?i��ܴ �C�����������q�؀��P��<�Ř���k�Ri�G�	3@��$�ZWa���*�<K�d7唚b�Y�i�\B*X:��/����U9}��G��CC��븛��fa6b�߸�'(�ڤOD�ڗ�QgؐS����g���G���3�z�r1�R���/�k.Z��,vp�X=W�wIʎ�Zr��"`q���%�oq�l(�)�8���J\O�����Ң�#�q&^��LO8�q��
���n�m�89a⥱3�4�z�u�L2M?G9�sZ8�Ƨ`"�g���D���"\{I*�B�Ḻp4�A���2���?�q�qwRz+���c��9���j�!;0��# �孞�,R���� X}��U�j�+Hɛd���5;�%Qu�c��&�<��EҪ�����=�J9�b �?�8|��=֠�	�/����qf��&r�t�:W\K��͎P�J6��\7�(��%N���e�| J�/8/yb�?��T��^p��6Gz��
'�3 +��d���D��5wI��J���|��I��4+E��N]��u��.R|��A��5ȶ��l	>Ɵ��}��X�f�7g9]ƶZ�/��SOIC��h������iM�F/+�(��@+/��KP�34�E��3��΋��+�퇞�{�1BE�&����4�	�Ĥ��̪k��ܯ����j>f��p9��̽h�%��0t@/�D�8�Iܡ��4m� ��U�d��j�T\�6?�����ɧAxa�s9�����HI��*"�ʷ�o;KB5�*�́�?�g	x&�o�,0����xdGC�	�ӤC�����m>��Ear�7�~�rf��U�w���q~)���s�"��%�Tڙ�!B�ݞ��˄*��LE�Ӽ"��6gB��Ô���h}i�Dj��R�����0D�{/���h"dgG�W�	
�ǆ���3cu���F\��h L4��=!~���/p�h������������ȹ�=�o}�V777+�_I�Erq��r���@p������'�7�m���8|`L�7mzqK�%��B��ZMS�`�6��:R���[��;C�壻0��A}\e��v�Rg9K\�at���;���7qWw,{S:��/��2'��3!R�-�id6�pM?-����U�q*a�/�)�o��{��~_�oM)�1-~)�  ��hQ[EW�����3c\X�ً.�/��j��80��#i�c�C�@��Է�M&Yܿ�Zd"i7*A�C���D��[R��z�_���W� ����b�i�Z�:���� �I������A(%��_:�U}!kp�T���f\ܣ�֍�iҊU!�0���w"
�@�M�wvz�ƽ�È,p����{]zﻗ���)�d�B���W;s���/�n�r	 {c�f,K��I��j���y�,��5��0)��PY�Ԇ�	x����	}V���BT�単���L��~�7�æR�QBZ~��Hhb�-tꇩ�G�!e����y�nm�8�.��V#t���E� �&o�M��)~3	>��%�M����C���JH�����M���J� Y��Ob�1�wvI�gX=J����D^�iX�L֘�/�;�P3�)%z&�0��TH��Cr����S讫~�F'}/#�i����U52��1+]��yU��'���G� �lakP�Շ�/�����3b�$�"�@t�!��lќ������ny�E�|���$[�D�p�<lJ��h�x�=Z�:Kz)?��a[;r���sщE�P��oX-M,�W�ۘT���������*�k	�,��R��܍7W��^oA��]w�u����`���Sͪ����Ff�E*�<$�D��h�j�y�?D<@a�)'�^#�i�RHq�!���aR�;��"�u`s�#²�1�y^�FS,tO�+��
�fX0U��Un�2�8�F=Hk��KiVݍۓ�I[/�d��q�����@zpW��%_I�5;�2���<�j/��Z���+�F2p ������;p�:K��~�����~��M��1�"���I��4'8�y'�h�I�)��z��ٞ��y���ϙ�j�a�0����E�&N]�R�F��L�MvJ&^�4S(L�T�D�*/��G���N���vG�����O���Uv�M*!;!L+�G�9R�P�}<���
�AC#�����S!�JCbR1o�Hv���iW�0¤��^4���i�uDq�ZV��W4�I� �� Ż�-����?<���t�T��Qb�G�:ڑafءd�A�x��Q����-XLX�-���ۄ6{�������0_���)'Hs ����F-Ѵ����E��4����AXRbѣ��ka���a�h��kф�8���2wB�}!�C��\�x؏/1����^���%�w�EW�/�r���hDu-��* ���G
^��V���1A�]Z��v�wOo�R{������<�@n�m�3vJ��H�U�w�|,F3)ޜ�"�p!�"���M��J�|�%ʼ�(̜A`Sw0��b>�眂���/55�)��%�iNN�t��\��Xc�6O�{��l,Te ����v"0`4y���ފZ������~Z'L)�k5[�(�n%��?0�kѵ9Z瓳�[?0R�YC�k����Sp�}�{K��K��?K��-9[s�
�\�GN#"�M>������L��w�{����4j#�swA����/g��i�Ґ���b�M�3���
�U�/�^5��*5~A(��|��0�����	�$�̹:��8x�:_&$��ɏˏ
�R�m���k�
K
�h2�ݕ���zk�h&dŧp�β�āV���!��8���+	:��A n���.�����\L/�y�%~�rո�b�g����R��UWq&�BMOv_��+iEMD��
�ssр[$8* �r�a/�}�(�9��>�1��O>�z/���5��i�9��%|}�� )��l�,+�j�Dv�J���Yel����b$C$���*ա�ߓV9֞����pO��;^-dh�7&8��U��Ƹ
����'sj�즦]2w[t~��{������4��q�CY��V��mH{?n�7�%]E�X�48f�T�'H� /(����2��3����y%�D��B?��UpѧD-����ן-\���rW40�:���_�A�r=FV���a�Ә�h��;l-;U��\7j[[�?���\��b�ʬ���n�&�7-|"\4V���K����H�B��=Ƭ�V����R� 4�\�V�DA\��P��i�n�P��տ�v�(1/�����y*%����t��C�h�s|��֩N<(g�"�IX����zyI�;�c�|$FO���5ww������sZ>E@\j�f��<�"w���2������8M׍$$��\��e+�%��%.ڣv��rE��LG��ɱ��(`p&[��o+R<�xT^�w����yVL�������!ye �wF��ʄ=3m�I����,<ϩ���`K�����#	ia�*����o�3[��繀>q2��*���U�*ce�){._F�J�*h�OB���V3����c(o$����!�R�P��˫����s&�%���xw�j�͹dP�L�:�r����)����?4���!�X�?��yJ'3����+�o��л��,��~l& WJ"��S��	��㔁���d��H�r�}F.�Uy�C��.Zm�B3�h	V����!6�9_Gg^Ȟ��7�ǯ	�-r�ļk�y�w���2�_LM��&������F4#�؎ �����bA��S�Q�Ơ�Q�$c����z�+#����n��Z&͍0��+��Q>�����h�ma�ͲJh9�&�RJ�z�~O6h�E���{�0�j�x�nb_J��εd��'�[_�
� �kT2.U)ۉ��v�_Ԗ��j�p�q�"&9��G�n�r�H���$he�s;��F�L�@l5?��Kc+@��F�M;�LVP��O�闣M��/2D��
~
�4Y oI(ɽh�I�wn`��s�1b�r�q��n���l��A�� �(l�챌 ��
��iўE��*�ޢ��w�D��]ts�a8,V�fz�P�B�ՙ�z�QQ��-�V�޼�*ʀ���@ T���U�Yq��v��B)���A�˖��Z*��d kZ6v�UА��+����X��"��t2#r����5s������'�vĳj>5?l��;UdNX�#������w|�Ȥ:s��*Eض���]J�*F�����?=i˞���	m��憬�x�/
�a��O��//:�h����ͱҫ~ �� ��Re �p{��H9��r�{ol���5/�i1�'�h�rX���b�(��U�p� P���ΒS�ڭ���K���"�-�����}��aN�mQ(Jb`*�-%7�-n>zs�:�ɉY�or;��O_+,T�n�%��@Î�}���J�c��#1�!3~u֖���-�+��[pc�l%������p�Pѿ�w�� F���V^����A[v�d\��8ԇ��/�c)���fs]�����8�.i��֦��٫�y@�/-���|��	[�V�	���O�P�{{�C�>k�!d�ڍ	0�#�hG�f�2}���9	|�ctW�Y]��2��кDI�g����:�e�&$���}��ߨ��>i�>��y~B����2�}�+�iG���[���8�P�"�}oW���3���M
йL�����Wip(�����lNm9����;��ȫ��t(��2wۊ�7�J��F+@̳�J`9��M-+����r�Lr�*H&H�^#�]�V:��L��`��&+M����6���o�W��=�D�D&�<��[7u~�'�ųIʥ#\���&�Al�Wr���"�?��� �2�����~��n{��7W?aX'l:�&x�6��Pnq�sG�g�D��L�_Pi�	��� &i�B$(؂_O��v��V_�ԩ²�:O��T��>�q+�c��}n=��B�T2hZS6e�*G��pp܏�@�8��gˏ�.M��0w�eӶ��E�)�y���-�#V�5M���p��~yh�}�X\���X�҂�/n�w]�Kh��Bl�&��j�)�E6��ps9�G*P|��b�y�pҏ�"�l���آb��|��㊃4ʤDq��g�[��~Z\��-r��D������@
����b��tg3]L:C��b���`j���<@�l[Km�#��`���t/���Z�z�k1��kV���2*[��!��C˗0�4���@H1f\�#�&gG���V�("�E�~$K���!�7C�v����̽�=����FfI�~A�)`a�[�)�,��T	�~ޖbi�V��u��p�$���:P�l0����{�qٴg?���(}bW ?_���r�r�e���PG|���U����@X��w^���޸Z�O(csE����(}�	jq6h�aR�����Psv>"Od��5�����0t�꠽�f�v�3�[E+K�79هSD��}w�2�M�8��ș�y�;�^|�
���r|��fB�q{����0=�d�-�}FAr`1-�]v�X��i�+�-z�����F�X����_W�*|fN>Zq8��d��[�d�l��I�+�
��dŲ�_6��Xġ �J{;ƪ�"�N4��: hM��v(���<��_\G5��\�j7t�Jw�s��f��s�FVH|��ݞM������RP�C	K ��JjN
lg�ۇ�_��q}4b��I��]�]55!iJ�D�)M�P-IY�x�<����s�S�2�#Wg1[����o�14���י��ey�Y̧E��W��yߓ�㱰,{,�D��U���;z�	�e��GD~�wΠۻ�Q�[�[!�Y���ݿ��t�qP�a��_WE
������g\������3��l��S�k��w�āN��H�1��wO3e�x��iA:�����r�r�u�Q�pS��W'a��5Y�GP��[���
B<�
�"_��ቇ�J�j�ˉV��
����Z3�ON0b�쇶4E��`E�챉)r�`�wD0���h<[�K���1&Wc@��!`��1y8�c�WZ*�%^�J}��;k �Ƚ����:���W�}*A
��8�gn��UX��	8<��U�D��Id���I��
T��I��(��,�E<!)��HU�=���f�A�~6���x�R	�s�M�0����@}�A���CT&�m��O� F<�/6G.O��X��R�Yv3!�k�) ����\6G�z�bnjՙ*�(�f�Q~�P��&���wׯT�<('w�G�i	�a��.�������G;h�7u�$M�v�-<q%��eLz:pm�"�(���ڍ�jVH?��
�^2�Z}�9�ā�j0`���B.��A|�����YL�,(]���,��8)#A����ϙ�g�.��p�i�:�J�A\ �/D�e�7�� �)�xO�T>Ǽ���A���[nx$��N��m�j��\��);y��@��r.0����8[�� TVj|�;4e�"���a���U��1~y�_ �����j ���,n��=S�R��S��'˒����:A�G��@�~Y���t��i7փ�L3i�ZOj�>=�$�!��bu�1)oU�mҾ
8r���@\ӽF�`s�f��&��p�Lfj�<^�5w�PaN�~��b�`L�pz`�n���Hkr���ؽ��ɶvR��	ߴҞ�.�D�Q~�ĸ�s{�c�N�!�&o��� ��y؝�~YeS�����3A4��)�� ����lh���J��S�� �N&�(Q�*�D_�`.0ss|�]���hx���P�E�5PC��td��BL��5���d��D��I��>��YX���N��� A	@�@�BW�<�`&�����Ү뉧+��!co;{t�<]���Ӛ���7r݁�xa�#�5䶐B�� �,�R�s!�O�u�szӊ;�囯�n�9Z�����&PU�E�v/��G����k�ۜ�+$!I�Bi���E_g�-�����Bh��?��2�ʮ-_B�@�u�����{��{{'��`d7#��^�÷!��G�ΦF���.e�%�����P���gnB\��
{��}���� �:(��V�%�����qtcq��pՃM�;jW������.�:}�:��P��u ����!Mm��J�hєs�u�k���_��KNEunܑ�e!_�)+�ִ�|�IDPSR`���c�B)%�c��7÷~i{+���̿8O���W��K��v�O ��6������U(?{����2�}�eӨL���D�9�E�Eňb�`!�er�?���ߧX�)H�O0xrgJטU�m�$��Oܜ>���*�Wg��ƿ��S|��oO�N�W�M�C��NW��c����=��?�)��^b��gƙAC��,�;Sa���^ٓ'���:��l9�\C�W�f'�3-sU�Sڂ�ǳ�v��w��w���B����ϫ���ݜ�)���IJb�ȇ1R�!VKN�n�q>n��8�]��t��>���b��ѵ����� �c�`���:� �-���kܗ~�-p��ҽ��*e��X8P9�y��� ��kݾa��1A��6Y* �\�]+S�V�mӿ:k�e��v��7�۬hP!-��]>�]F�����}�l�,��Db9�1��ܰR7�[�;n2���$�,NƷ6���&�^/[�܆
�y�=qv\t�����|�����V�.,㦦2���%&���[:��GV�OۇEb!Zei��JΔ�E�?�T_�p�_���=��w1��c����d��r2؆�:���b�K��i]4�'&Q�c��H��c'Q�a��XsJ��v���
��ڈ���*��Y%S��J��I%��ʘX��x�&M*a�&�ݮ4�[_h.g���|w=��=���L��u�J'Ʌ�>=�s�?��ȫ��!��0�üòaH�ajT�Ȇ"g8[uO�uW7 %�l�^݇���CQ��f�y��)c�`#wx��-�ޝ���#�>(��r�&MEl-E�<�j緗�KN�Ox��B0����]��>�dr��z�q�}Mǹ���� �خ!j��E2r�X|�^��q;^�c��	/ΰ9�S�XO�	4��O�<�Ԛ��b2-/N쐎�[sd�� Y�M`��HY]dh�9����3\E�H�ő����zެ#��V�8�_�]�������ٮ��q���+����c�9
Ax��4�]�8� �&��Φ`���YXF(@�b�W�l����������A�̩��H�����#����W�lʝ�_>5<�&��R���:/�AAro*2y����n��=W^�aZ�~k�|N��r.g\jM���)�=h������X��h�^&-�8/�-Q�%����]���)Q$�����eC��������Bb������q��.A!��~��uN���"�~xA��A�m�����3��R&7�ޏ26�Rٔ�L�[&]�8.�"1�/�'s��|�x�4���y�D��Ez9~Z�$]��1�ˎ2:�o�N�G�r�nJa���8�kC�������!3��0QmL�
8T�=��K�DN���+�M�hJ��^�l�	�U�����W�	|^��q)����c �� J�jCD�F�~�"���p`gv�D�@ޕ�o�;rv1��֮�l�)���"G��		k�����ѳ��xd�N�a!%TN[&Z��fƿ��k/o0��bA[y�'��-�aQGN'g���U�@1�����
�����HW�kd&c����ܾ�����dj{1�h��2��:Zv�TK��N�Wj �yݝz�D���[4iz�4ۆ����[G�%�L}�L��+�6�����t�3��"��c�1Cho�2{�=�"�����Y�	M$��U50J�!d���_0�x����@G�x�_���� o��:T���.k�z1��W�=�k�$Z�,nO����cJGXm�B� ;�f�����R�7��C܀NkL0A ���&�u��D8ǒI�]�<aT �*VڨW\���֑�G��Z��wN��^<2�c�l9<eټ�-�k�0VHl��9�pJn�q��3K|�C5����G��ÏN�$�jM��d2��J^�]D�;��\7r����U���( �)�	���]��*ɩK}����s�b��6�������M�9!��4��3=9*p�Q��\�(���uA��*%� �ܦ��&�҈� @06��yK����U{6�O�e��{�2�V�Ç-Z�X�@�����$⭜�r��o�c�x������2�e=0��E��+++�[�=^�BqU�"�����jD�=�����P%G�%@����uw�K��OO1�xP/��O�Q�I���Df��|�hO��h[#�t��@jB�26���܌�LZ�����ɮA���SV�s=��DGk�/���oQ�Tb�()S��K*F�#��JK�:�Ҝ@Z&Նd�z���]�OcX?2g!
<��Wؕm��Bԓ/�!SW���AE��n�ʜ�����)��0u�MLC��za�B�y&I��/N�9�,�W�����A��a`S�Z���ng�o.v�5�.k�0ϐ�B�j�6T]9X��P�����~3oe(:��y����L�xG�r)UgU��]ν��Kh~��R� �\�Ǘ����:��]�	�s,5"k���W���y��0-7�3H�3�ʩ�����c�=F�'J��m����zӉ�����̀�cy�8q,����|~�G�dVk���p� J)w�K	��W�;C4�)DA�#a�2oY���>-��2
�����b2�%&����0<b���M�8��E�}("��&][L�_���B����2{rm@��f
���bl%�]�a^�SE���`d�����p�rFQ�ul'�/�~j+��i�E��8͞���â����tG�A�9����@�Gt_���$�?�bO r�3��	�'��!�]�?8g���&���T�VEJ�<Ί,p��B��[<�ݠ���*e�9��n��|������;�_K�V�ԖD̞S���+Ya�rEO�!_
����BJ�U֬���B[F���S!Gi�A�?��	-����(بmm�z��nwv�H�᮴���|�b���N"M��w���b�$��ȣ�b-1s�(���x�RȘZ�c<D�zP���&#�x�h#qlB�z/"Bn7#D"t���47�̈S]C$��K�2�D�����3F������c���Y�b�.
�-����`���L��`�͢a����x���(��d���]Pښ��C�A�+@�i-��_���v0�I��1���2���f۹�E�d�� k��`�^�^�~[��Kװ��@� G���KR��*E�h{I�����fR�|��.1�}��ٽ1�5=jM��o3��z���n�-���m�7hln�F����G>�A1���#���0���*���-?7d(����n5%%����gS��Ԟ��$=���Ί�):v	P�|��A�T0RsD?Sz�����cc7��3��ͻj}�g����nHgl�GNsa�g%�����[��1`L���:�;נ����@V�-;��������a0�SJ�L��͒zƽǒ$/��r��+�S_Up�0.���j�Fs��I�t�.7qk�����Xo�B�'J���ƈ�'h�mze�S�m���'���6�� �,�-��%c��s bS= #����9�NԄ:�p�ɐ���]	�A��G�bC�r�]��$��D�����uaq��_�|�N�TDe"��8���xEo���u�P�w��
{�q8Pa��~�VJ�R.�Jb�x3+�BAmA��a\Cߍ����+���΃�u��撌q�㧻�
���z5���~�N>��pA��$~�+� ���"��8��>Ǫ�3���� ���[9N�!��NE���Q�nSU�6�`pM�b�ۤ.r#�gtIC>���8��]ߔ��>`}��S��v3�䧛Iז)�DAr��:}/�EP��qzA�5&8O5�f��-���Eh�9��Hc;*��-6���|X;UpIs���hQ�/�ii�vI��PiK�^��O�=�j6k4Jl�#��O�=X���u
��#ղ�"�y�fj�x<�Z2�Ն;�q(r9�˫L�}Oa#<y W=�Ҙ`+&�2�d8�@����5���%J���ۉ��+��ڍ��u߰`�L���IK���*r��@t`�pW�g\C�����R��
~:F �9�*�� h�Ì�ӕ|����}��MR�}� *�D��b�<]�N�	�ST��q �.�$*���'��1�ne"�$e���v�4�J"�|��P���b:�7^�t�1���%u��/�D�n�;_"4�A�� Bv4_��|*�H����\=��:$��9�ڄ�$[T�����K�(u�q�)�=s�T�:<|,�P����ֳ��L����/�/��[ۂ=�7H,���ӱ87ةz��i��2�N���Xڂ�Wt���!�m��`i���ɛ�E:�H_x�wm|�+c��}O��xKFZ���k���b��4�m��jM����r�
���\J��e�K�lH����d�k�Q���ئ����BC��f�?�a�[4S��2���pwz*��]���5Y�����Gn��D���	�����$<Z;�b�N)r�h����Ԅ�u��u��ה��iɯ���ŇԽέ����Iu�m��L��f�n�g�d���Zڃ2��*S�(�Y|��a$������$�}������������]�,��mC'�}a�$lQ�M����2�&.����j~ѷ�,j!B/F���)�8n��I�ܦ��t�
�N@ /������;4$�
�m���cs&�1�M4�>��6Bv}�����(�Y�-N�jk���Y�[�Mə��^Ĩ�RڿB�<o���8z�4�L���������A;v�O�-�������vys�޷t��?0��Bc�&���gHSQG5ʴ�=�uI�,1;�*�U�+c ��ݶM��,2���M"c�PL�,��c�O���ct�4}��nj�Og��WZ�hd���ǿ$���߈J4��0Qyd=&r��r aЭ�G9K�N��-��/�1�*��yn�P�~mV�����ׄ᤮7"+p5K��t51^���D�0���<� ��/S����'�F���<m�GZ��hi"�U�b�Hd��D��1ӝ�L�>l�:�]{��S�!�06��~�(�:1MŊ߃� �y���o��,˦��P(&Њ�Tʡ1:iV.�t�-N���KnG]�<@;�.��d�(��^�,��&20�Z��D�����.�je���T=�b''����T#YV�r�){w�(m4.O�r��`Gz:��rj�B����]���5��v�z�#K,VI���v.t�|4��AVx�y�Ox�����g&��o��g`Q�s@r7��h������ųX����v�	��]6A	�pl�՘T�۱Ər���{F�x*�>7��0_DlP	ZH|���jF@�%��(���� �u�%��3b����5-����fFh�³�VaB2����|%/��}7f�k�i���?R-���Jpݱ\df@ػ�,�%ĸ~�E8�RQ��a%C��XpDK�F����Xܫ��� �y����/�2*���ok�ϡ�+PL�0�[���$Mޙ�!�S���H���k����i[8$���
Ȝ� �����qc*pg��-[[�B� ��/��8la7����&1�T�T��3�%���RL1P۹{@��Tm���w����:1%%[���R	�.��'�h�~Z�o��=>Mxu�+�͚�>�hN���Z71�p�_�$��W�ie��{HÚ���2����5u^�����0k]� �I��r����JY���ɲ��l­A�e�8���Ѐ����O0�Bq;�|�BOş��d
�F��� �Z�u;�	�����(�şjh�
�Y�&�������Ӡ��A��	���++�����e�%�J�Qo���9g9V�{Q���2>9�h
.%�lf�E��=NC�����	Zv,����r-��s�*�ᖿ�:����b�* D�S���;����a}�Mw{늁��	�5�Q���6:2ϥ���,�I�,�IK�~��<�H���i���P}��7l�����˿#A"v�QY�"Mm�)0����Bv��a'KRH<��$�PE�y+[�ڵ��a_,��r����.�U6��M��&��~�����0��	�^m�GB�6�uH��b�F��;'	����)�Z�P��12�UY�3������Z�"�G$a��u�^��a�s���:~4��S�>�o�F���<�v��4w�_5�v�]���e��3�*oH��n�2�!j�kc�3Ғ�_��`?G���Xd�fV��7U�a����M�� c� �����Wx�]��WA/��|漝�e��5�ZE��8�PeJ��;��H&���G���񎸳��#�-ZvÉ꫷�������Fdh�3"D�6O�އ��rډ��E��dz�w�2�%v���%��5h�~߼��QQ���\���4�'�R�}��;�_�4{yØ���!0��?[��$
P܍���l������R`K���k���ތ`�Ev݌E�[޼j5dZnl;9ypL8I6M�]��v��e��j�#�[#Ky{I4	t��ݒ jկ�����$��RH�
���#t�/�q4�hn�s8�]8����c2b[]��2.�����M�R� ��\QU/6I�q�7^[�9�e+�TV��ja�����	�˹?�g���Jw���E��S���g��(�T��`�eͮ�F�,K.��=ҭ����/7C�p�֌`��γ�WA�k�7���`�r#�<Zo';+l�/L!����J���C�4XA�Y_�@��P>�Uw�v�j��̹����beA%�I��1pƔ�:��@1��*���Y��p��z<�Xx=��+��pg���A�h�
�	�Kzʰw�r�@�Lv�"��� ����!i֊���ZZ	�#�
���T�Z{��I�p�����45��]W���es����ۈj��04�'m�O��bti]X��zM-c�bre��N�G���`~�0��py��j�t�� 5D����1��h�.���qr�٢Z���sLD#������Dt�~�7C�&+�v�%L��λqf��j�8�ƺ�zS��ٰ3z�yk��=��|�>�W觖��`mcD��YQ�I�;����t�{�������v+��-U[�2��&�EQ�/v4��Z܈;U�Y���wʬ�Qn�F��x��/;��p-�wS:)�G�u���1'�3'�����7f��-��͞����3VN��=	ۮ~UE�]��*�_(��y�n2 :��{'��a��[�77+���,�)@x��WVU����!M" �<�^�_i3Z�-m�O�9]gGI�+ϹO��$���ɮ-�8U�29�4/��ѝJ�<b�dv�!T�c�i���]�U5	A7����9\������mV�b�l$�G�����`O�W���9ɨ��wӶbK��C��X���UX8���!�Yvv�zz�O�T�|�?]
}N�A��O=��oJ��AQOL�{{�P�J����ݣY�ӵ6��?���NOYؓK��Ns�T<����`�΍��M�w<8a1�S�af�^�J��+4l���1	�uDwh�>�q�T�,�n�۞V��#�"��N��@�Y���u�+��R"�b�$j����K{^�=�"$�I��(-��/�V�αhBIIc����Pً��~�إ%��G� 	�@��-& 4ק�2���V�T�	�����lٷ?��ϝd>-�T��à ���͸_�I��^F�*��+�����KPS��zh�����Ֆh�&W.���+���L6�w1���-\�>Z��~l@��LB�8�z���
��\��s����k��S�g���H��mu��`��,X����)o身"	]�Z2�@�q�9M��2�1�����8l��(e�쳉�@��{���ʶ��L��	b����`��j[]h�a+WB�	:s�u�GR��+�/&�m��F���R����-՟1%��hZ��Z=���x�U�/�$�����y�Z�����a���ɝ �Ƈ��5�,���i�;�d<����d��2�B���:@S:�B6sӄ��3|�m%�??ҁ
4�|�=�M@�I�T�8+i���\����!:��z���E=��p�A������s�Q�L��̞��YI���n��5�o�%�tf�����7��0�)�_�Z�ѻ���^ly}/���(�Q_�g�X�Pi�Y!G%I�p�UR;l�~��~�G[k�C�QA��(A ��)UR�Y��oF�	�m�x�LKK[��tФ4+.��@��Ǘ8����"E�%T�f3��(��6%�9�����p�[WA@�>��&Y����5��KBB8p
�i�����h]�V�&m��Fx�b���H�t\��+��ݡ�̢50��˓�����KE� Zqk~�Y�T�Ӏ����4��rS�S����2�~����A������$�BX���LSy�:���Ę���ܚ�;߶�l6�k��#�c��B�zu�17�r卦I����	�b�8dgb�:'��px�Z��ҏ���^`�I�m���ʫs|÷6��T[���(I��b�4/B�D�:\��Q�6z��;����(�����%�����6��@U�� 
������$aV��`���jF����fO��U׌ª�a^_8��^/���O���ŚAx���3-}82Ҳ"�� )�sjuzR0M�Ʉ[���:��МJ�6�[������%JjC@<�y��i���\����$NҪ��Ni�� {n)��Z���0
�s�	�	w�E��p�eN�Hn4d{����z*�����ND���l�W��XR�vĕ�� p�򾣳V�-���b�`����?���E�1}�C���57�X�8����ɀ��xx��8Т�e�Zui=�T��gH'? ���vӳO�KR������� 2 �$��(I�XdH���%��U5�:m�L����9i��G��,�%�?V�(%��_t��a��V	a/s/7�F ��ပi��r@��dS�(A��'� ��W���0�X���ŗ��"�[㢅�*�a�(%�� D�������պxd4�G��4&p+��6��1�)S��*폛Cʔq���IJ8�'��hd�kP�,ƶ�/�k����!�@Y�EƑ��Yo���~?օFo��[��1Ib67��ܠ���sy�i{jl9����y+�}�@m��[O����*+؋A���;����l�fsB}6��D�%o
&�*R�P�d��c�ũB	sn~��X=0[��eX�R�W<�֏^:q�*a��*u�U�r@�����eW���ىd�2M�.b`����J���|��&_�q��\���m�{�T����}Gf�;b���Z�F������+�	{�������z?�=��K��^�k���qDsi�q+�<�*<������l�>�Ɔ��ߐI�4=���m��H2����f�~�H����� �2�62	�zm6N#�+��ş«�"�*,����b��אT���p(��íb0:�-8WD�yk�ܙ$�ġ՘�s1l���w�����(4�Cݘ���y�i����˖�S��[QG?��z�E!vLsن���70g�- Ʋ�~�T,�tl�3���,�3	�Z����+ԚMaX�aJ�,ǉ���C
�=D���=Q#��۠�4��Ə�r����%��	w��%e9���[Se�I��=�r���jq>�W�1T� ���b�N��+C�:���a$�}��z�9��n�p�/���q�'���ɱ�5���Z"�/�979���晄��y�I�1r��8��. Y��'`���0���HX�|�̑�<���6�c{\�m���ϯ�5���A����`�p��k��P7m;D �2m�-�ees�T�+�/gF��īs8ɏ���_Pa��͆z�w��yik��R'��tZ�/3��i���@#:��S����S���Ȝ�v��Q�Z�-�=��9���М�b��"1���b�J�ݥ�-�$K�v�sw׻�3%�'	P��\�?�ģ�g�@���@��y+m"��܇1���Bdf9-,'@
��"��oWw���E*�"�!�������h/֧���v2��9��#��7(�1�?<e�nDc�8=Ъ�������1e�Wi��L񌷟��y���7�mÜ��A%C~�b�U�U7�q�{\��d��;��<�vZ���Q8>sz� �{lMzm��)��'7%��d>|(u�_{)̟���,T��$�p�/�e5��7@�ǟ���a��{���e~��)�3�ՌF�4��)��UL6ogv�u�����Bs��>��U��s�{�2ɝ��"��(K���4Zd��!f(ElRL��`��!_�q-���*3no��_���\�A�:��Y%�]�B�������џ��WlL�A�S.CM�X�5��M	�4~d_<脝-Q�����X䉑���M�p��������)�Z
�#WV2Y�۾�~do�.���6�&zHY3��r-L�)�40
4����D!��wfwVN�m���S-%?�p$�v��62�PY��t��ф'��e����\S=[�
}"'�sXd\0ST�L~I��!]w28?�Y�Xf�n,��2q8(�Bn���S�@�7�I����$����L�o�W�$�z�)�dr7��N��4>c���J���m׍"n��.s�BSJ�/5˭G2;݋�_���*3|,�fL��IϏ�f�$|���|o��.�K�Te���"�o����- �	
��D]�W����D�(5�~ƛ@π������b5���.�h��8}�8b(�;����V�z�4zr����%x��
�����p��~cA�p�����1m���ؘ��<��Z���w|��,7Vdi&w6�w�=��V�d�S�)�su�#g�ܐ|!��W���A�$����W^lF��"��t���;�Кq6U��M<J
6��7{ʥ"��7{��c��p�:�l40�Yϋ罕�t�N����ҝe�4���Z�I�ue��9�ѕ��e���Ί�l�4w��ۧ���ڍU����Qa���ݢԉ�P鞽��+�lt�b������K�t`̠����\�K,���J�栒}0K5���Z�"���4�
x�n���N�8�h����*ڶL7����䓆'�"����e�"�9ޜ��|�%UZ��HS}���,I���\{^����t�B�c���ܣ��
\?�I�,�%���.����S}��!���L�d��/PM��]ׇ��g���u��Y�J*��gG�)ig�k�Ż�Xb<�Z���$��e�CV��@܉Ê���xY��F_�z����Ж_�ae+[�}�B�Уp����B43_�Q��%�&���7&Wr���לY�j�
����(���L��pRw�S�g�1�ܬ\�w~,�9���M^����1��se~�||��W�Izn����-�Ǫm���j'�<�pM$�5��2�sq��Տ� R�x�����˻����Y�4%�>�:*��̄���X�]t���ه�)�#�y��(�����[8�!�hn��|�?�Nm:!�=�,p�`+���V�t�t��u��S�����c�]�I��R8�S~�m=W[K��g�����)��TϦ�廁hb>q���6��K^�1�y�Jkތ�4p�[�I���X���|Gb4�ժ'���`�ݰz�2�*K�w����铏4���8���:ǬZ(�Y���������v�[�x�+ji?��aGfBN���$"G�nA�ou��IME=���l���������_�1�Ə�<1�!K"�y�'Co�V4�e��G�fZ�b5'�_ ���,]������Rs��_:����:D*hP�[ۡ�<$��]�y�<G�sQ�L�wOR��lq��{tF�Be|g�h�����)9����D���d���]!�v�ƺ�iF�7rR��9r�Q��?a�'Q��s�0�Q^į
Ԇ�0{���ݲ޳	���u��>v\TW�6�H��;E荊�׬�g6�:���#�aM�ڊ^�g�p���2*mv��+�
E��_a�~̟�Y�潒m�̿��S�rU�)h��Wګ�<{�K�2T��ʍ�`}�R���0��@�� ¼�$�\X}����"��̨g�^h�Bl���V!s�xeD���h �e��]F;d��G%VӍ�+��E�>J^�" � }�
�w#2�N�yF�<��#�z?�]E�X!��>��!6;�����LJ6:����ͮ��4ov;�֦�/�Ʉm���)���� ��DnMZ�ɺ*����y:�]�$�x��N�����R�����m�D�&����!�A�g=q�B)5����Ƥ�.mfz���g ��z��ݢmG�$L���W[@޼�g��5�f
q��Ƞv\ED'0���0V@�b�-(vL������%."���d���zq)�6���+sZzg�(�e��v/�T/v�� ۝��dٯ���	ɐ��'� 	jw�	K�=/*���-+�����K���oj���G@5���)�3? ���8 �`�llo�
�s%��_���,���4���e����W�<�Nah�\�����Y�D��J�� �,���(��U_��j�V���	~�����֗�����[i>�7����Tn� |M��V]��@,P��X
�t
Q�_Ã�|� �%b�j��&;o�T�'.ٷ���p(�t_�W���:�t��o;�!9*I��
�P�ZJo�EX�Fc�mۓ�!ؚS<}�N��oh�\����(��rTXM�"��ʺ1+�4�TM/c運�M���^K��}^Or�����U�(�*��7r�`���{�F�����%��>;H!`޽{T2������$��Q{t�0�wJ��{��2{��&O������v-N2d�ުhf��S��^�V�z�W4�l<��W��#������	���>f�9n���O,H��iw�h���4��W��{ �#���4:�ۯ��;�;�z���׵	�#{�̕�*]@teoq�\=_jm|$���׀��������ƧVj�^!
���̹�
�-޳�@E�q��<F��kcj�Xk�,tC�x�S+�x�p;
�2��VK��7��4f��Lu{$��ln� ήH�TW���V�4���A��+@�i�q��+q�d�:�d���Ñ�$@�]�0���/����Y�d�>�=k�&֤�
ڶ��'J]�2]cv;׏$��������$Cke�5@��>�U�4�����ʙi<������u�zx<�e��m�E����aB㜲�b&_�I�al�Qz!��]S3��}�c���9������կe�*����"�6(uG�]�Bf�^G���$�Ab����C������$�@=�_P;�]���!a%�X��w)���N�?ɂxF�{F������%Q����r*�|��z��XSq�oN�/n$����~r��(t��XPU�oУ�9Il��yڢ�Rj�2�4SwN������f7|�ت�ds�tL,Vl�ҹ�D+�������gGL�ߏxԉq
B������'9zw�l|!3و-�E�D�k�Q+*2Xl5pϕrJ��Z�f��&������UsK�R`�Dr��ì��D�H�3Wa�?~�Vţ�%/u�*5�V��qF����)Ͳ78v�%!#��ɂz��M����g�@Y)��b3���Ȋ�,���p:^2��9��dKӑy,�B�<'����\C���˘�I����G�j�;d
��H�}���S�`�-q�u�o�a�I`5$���� ������ �AH:W�M\�I8d& ,���_�>��!���} �5(�������)�5��F�[N��)�F���76ބ�,��H�8�y���ߒ��d4̸e��oJ3��e�$�����	e8"WJ�]����S�3��l�[��>g~�K��N���V�Lfos��¦ϟ����Sn'C�$1ϵ��Օ2H�Ͱx.'({]��ecv����x3>q��"#�>���=\�)ݒ$+���KW^5UT��/����W�u��4����6���yn	S_����ݬd�w6j��K���(/�f<���-�v 0���5�ar��-+ނ�-�2Q�u���Аf���-��Ŷ.�� �(_)�}�����!��R��>!������F�6� ���Ͼ��/yE>y�bĉa�d 	�9��)�#�Xj��a!��=��?�y�[����O���������@�:��UJx����Y�â��qR�"�|���x������w��@Nu����?�/�S`J���V<^����H��t��`���`P�_;�H�Ȕ����a�:��� ���EiwEV�F����@�x)8gh�Q���f�~;�"N~�C���uY�g!^����{���Yv�Y�cH���E{D}�8��
>�/M��B�l�4�L<%
�|x\���[�����u� ����'ʨ���R���`'ޚ����Ӈ�� ���|p�����9��׹�m���O�[ !T���@��0�RG��w9a��S���|5��o~�P��R�Mo�"<��F�ɡ>1:$(��DbE�-`�<�2��Ԃ����<�$�°�>��G�����I�jἯ ^{59Z�H<X�T����r:�	T�� �N�)! �x��3{�a^V]�v�_�iB7��\���̿dX��@�n�H`0�/��4:��� tK6Wt��J��$��'%�5���yd��� ](��f����E_���T�s6�mf6�Mv8���;pklE��4���w+ud����v`��q]�U�J�Q<rO0��A9���ԹD�@��)�`����M�ov��C	Ej�����4���EI�Â��v��wn@E$�� G�@:�42B�Z�R�R��1k�r���)�+�,P���'�5���A� *O�7�L?I
��x\"� |�*�ײ�8�x�^�Ŗ�`
��`IB�L�h�Kl��c;��0g���]e��ĪKx��1)������
1m�VX)����4�zv��z;^ ^n�#��!Ao�T�P�[���ώ�%XΪ�����6�������������@PS5{��	��uu!4�#4��PoF�+mw��n���y�0��BZAd�����@Q#�
u�",����l�w^+��no�ao����/ͅy��\:
&?)`�I68vl/��ZЧMHr��4�Z ���Z}Ajծ����_ws�`�V`��x��?1sz_���=.sx獵���g@ü�Z}��-H��Ě���9 ̃]P�A����t��G���h�J��N��J�6~�(��k&D��{[�Z��(Pv-�K_���eC*�7�����?�[�ݽş+�iS���JBWI/��і�n#*���4�o��o��T!N���0��A�U����������7��,�#�V-�R��O^E���R`!X������c^��	5鐞� �/�Sڐ�����q��p�}W���pa����"ө��/�c�D���GnP���un"cۊa�d/�º�y�O['�q|�3�׺f�ܖ��;�̦�Z��i���k���6�Q^X��(���Y5.�A�D������j.�_���S�}X��$g�~�u
�>�����Ӝ�U�I\&�\-lǀ�y��D��l~�� (,-���wy)�rN�$!��ˑ0KǸ����81Yxk�H[��N5yD�J���X	�~pYђ"[��}�ؒ1[� Ŷy�5g,���Gm[N(ic4������\]�+j#��0w��� �_)݋8�({��q٨�����m�����`�����[���I�-
�������R��;�K�]z\���T�����AVdP�uV��(hQ_�G�qaҮy֣�_�=b��F��ĸ����|�$L��&!M�-k6G����F3��*���ďz��U05L��y�K��m��Ҍx��L����5��ͣ�^��M�	Ma������s���h�qM�H��lpl�a4��O� ��bo���y�$X ��ݲ�[�+221q�3D�,���M#*���$�~�����+ ������� Ya�:GwḌm��΄M��)���*���-٪�k���l��[[��2$c����^�\�r&S;5E#0�cL8�pA]�bZ]S���Xq� ��b�������g��B��/e�$I2.��a�<Ѿ*�Ǎw��|;��2�[
Sr1.ǧ�ష�'�Zت֧�n�O	 ״�#�BG�3sm`"��?���0�o����9B]a�G�B�\l�wEr���>'ƍO���7�wJUNU	��h�֢)SQ
��If�џ�����ᗛM�A�6I֑GX(W,|K�a����jG�'�6��֋%�`��j-nz��!�>�3I��g�P�RS����h|$E����X"��{g#8#?��%�ԑM� �Ⱥ�{�F%�} דG�{���d5�tX*��259�;���^V�qp��v�i���=�-P��R֮�t����s�F���o?�M�4��x�u,�SEڛ �tw�D�$P���4��$p�/�H������Af���`Z���fkn�iaHY�vW�(+���*�o�׶%����Xr��_Y�!y�����Ү�Y6�"?t U>�mYv"Z�<��xA+co�a�+��� L� !�L�L�f�0ku�	��0�jj��Qǎ��J�̤����$�Z��Y2I�L>h���j�W.����2�UӴ�����}u$�Q0�B$��ǽ���'�ֲ?��Q��@��D�y����M;VQ*>c��۾w���T)�*�b�k�D%��vQ�p.�%ۖW3�J�us��17��������|L=.5mm �`���~$� ���w�S��X�F��U��L� ���ͨ�^,�Q���ſT�̔���V�L�hs�n�a��<f6a��`��y	�Կoǌ�Ƒ�sb��g;n�t�~�&��Od�ϒ.̵7��Z_�zkӟ#��<�R��>��И�߷�L�kPC\��٠�-�Co��#w�
�!��	�> oNҲc�/�����l�-s�\#oՇw��h2�W�L��$}ġ;��}�Ҍ��wc��b8�dRk5�+��u��/|n�,VzZ��ynx�^%��0_�|��i��mf��"��$�+ɘ&o͆Cq�{�ƺ��U!�JyXs�{�f`W�1�X��x�Z?�KΫ
P`�����k�M��S�%�Ҧ<�m���,�s��ƙM����#3�.U��[��w�?�	RpQwR���7�5��{���W����m���B�ہ�?E�8i\�"��o�n�3j�� X�z)B⻠u�h�vP4h1T���i\b�F����}�i+�:��k�1�z ���g�n.׶0�D�>O	�"��C��&��bÙ�/7a��6PNU��9��hԖ�qBu('�N��h�*�
�W���S�2��H�n̮�1�5yPP�P��/	%�����n�&lk��N�Z�����p�POM�7��E��z}s�g�.�X��&�� =���\�.Au���� =�)="&l���O��%}i�.���a��Y�#X������c�Ā���^2��z����rb�!Ot�'�S�#�X��hzs;�I/��;GZ�ť\��'y�}���\�a#������e����;�M�BXT誢Y}��%>�����]r���ޯ��`�������<��<vh���0d���¿��T#J�E��G���ı(�8���+F�ME�H��k��=�R�h�f|��dxҶ�~`g����O�/Ln�Y􆎕ft7V�A(��[�K���y�Ŧ]��s��b�s6)t�By��ZP�:i�B��{�%�q�����j&�(j��/"դ1�zZ��x������$�&@mo�1Sܟ$�;����,�s���(>�^�a0�$�߭R4e��=k�ڱ��"x6�+H0��.�dyd�+g\+�_�¸täR�ȷ�e&n>I�vD�48�:P�/E�:Dw�:l ⷡ���C���`A� c9�0S���v|�\2 W@ BL��j��2z�4Ȟп	�,�T	�Z��QU`}��ҥ����D�]��)��?A����-
�9�;�1B)�&��,�����C�#�>�K����xD|6��
V�Ӳ�(JdN���D41�-̒L��%j[��	1��������-���0�"Mc�%<�N4'|�."ۖ,��H�c�l�a�)�+{��"��l3ކ/=ӷh	0�1V�=��cX��M�|ʣ8��ZЙq���8�1�7�>���zn��	���Q����h�f/goI0u�t�x�N%5Z1�|��PE�6A�o���V��0�c#&Lz\��3((֍K9N�&�����9s<��J��Y\�3��7��O�
ܞj!����.,5��5O�b V
,�����$~}�"��7�gƴ���iϓ]��;w�͑�%$!�c}[��x������Z+Ve�h�כH��b~�n|���~����zx���9	�8x�Pq��hy�x�n��Q驘�"(|�Ω@�������y�j������~~�m:��s�{P~r�-�|���l&��9譇�#�ɸ5pѠ�;�o����=˄d=C�X��?�S|�팺����Iq˅�*����Bn�r��C��-�i����(�*��- �=n0�������+��he+|��H/1A�����Z��V>�1��Z���I�vOե�h�1@��|��X���[#��Ķ�s{1��`���'�*��
2v�����%�]� �n���z�w�x4ڪ�:3��y�
�-^2�D�m��!���䀉��nw4=Q�u��lF4���R���C2�W�uկx��{e-�-=�N��t�Pb�B��G�z����޿:@��@U�P�V��Y��x5���!��w)%��}I�]��ԁuY۲���|���q���t˹JN���~�f-����@<>�S����S�y�3��&X����ʶ1%�&�����)E�*`j�`f�;��}��fq����=HvjO���5��wS�E��û��f`C�^�g2���QHEX��Y��q�_����Pc\����դ��U��T
2���:j�8s�W�&y�@2�<h���lcU��qG��ٿ�&|UBkԨ�!3��>=D��c��0���s��F-�~���!�%p��'r�(C!���ϯ���퉭����d<b���R��l�'��>�yi�L�l���7���;��&و_��=df�����(��8��~�K�`�ޝ!.s��?����s��k6L/3�G�Ed���>A���oT!N5�N�������/�Z:� p�:�V�i��}9%E�=�d�>��y*z����߁��//�$��E^S�4�\,���O�����o�/����5�o�,��<�!t�=e����J����m
�e�B>i]�*hD�jJ�"�J�~X�d%@aǞg�$��]��!NE�RSL3�1�B�t;����#��Ŀ�P��1��$�R
��4��u�����`>k/��N�`��zr����c����ect�fq��u轭�T6��L��a����)��0�F�''��**��p��7�����M�}�7�鿈2U�ăN�h�J���)�dE}�:�Q����ϒբ0�b��:"�P5�1���W�6p=��DA�0P�E�p@�jn���>���
��U��B���)��Qⷴ%��N��Mx��X��7���.	�nx*%��/����o5����>�V�U��Z0��|��U��U�y���5��9������w�qd|�)bB�]e�e��}beL8�j��!|��+IXo �5�$�MP���L� bZ͒�q`.�i�?}���-ӺRuK�w�9�c��
��	��{J��C�ŕnVr��U�S����}���k
e���0�R�k��J���k�M�r����݊�Z�!wt�Vر^��Krx�V��}�!���Rz+��މ�DPS���Y#���f=��
n`�.�������⒈��I&'��t�q�cu�%�|U;�ah�V~��7�}� �R�.��0@C�L�*y���}�6�۪���.n�^<+��x�"�F(�Aֿ�D`(��NG7(�y�,��2la���5���[Z~�
eo͢�ݢ��7���~����
����>�ۧɦ����!��ş�]�����b����QuF�*��ą3�Qu����􃿛ړj&̵L�D��ս�~�f��Zy}��EN�F�"4Xz�ot������.tA=�\Ж�����O��In,w��&��^:�G�c�vJ
Y��]6�H��]��"�٪��	����if�&�_K����B�5ϼjQY��&���fl:=�_!/)]��r%Z-|�XD5+���4�\D��f�Ϻ�>y�HT��W��i������pt9������>�.u���z9�[h�p�h�Q�4��ٛ��脾%(AdP�b�0����A�pBf�����[AV��Q�s�� rV����5oG<�{6��5���2�B����3J9B�2��z��M]�5�"�c��<*;mfA�
T��e���n|�)Jd�Ks�K.���&�M~���b�� �
����!�wm�����Ց���Rt�q}��bWE(4�h[|/�	��
Ys�
�ͭ/9�ǋ��/S<!�������%*� [�:h!
�FP˸<��OP�8����D��?K����v&���[WӯD;���I��F�N�K`_����C��(�Ȳ�h�aD�G ��[��P�����<'Gˈ2@칒�[�+�Q��6�|�i��cA�򖁴_�-Q���Ff8��� �̦��3Ѷ���4}�tP&D���g��@ˮK�+�p�v�v��]�OB�c���%J84���F�����Ḡ/���:����K���8�"��n��z'f�SN���;t�U�\_V0��j���U*��2�I��m�mR��ȵ�~I{� 
����]���{ ��ڱ*�㚳�+�,mu�ͰK��bm,�mR��7!�|}N�@�:�*��s�rxz$�Ɩ;+j Sr�ߩ�;5���r�zF�Q-T���X�J�m|��o�����:�Mi}���슈u!$
&�9v����6Z�"�`�uG��̰�QQ��IPd�gGIa�L��tc(����"����� ���˒�Ɖ׼Bw�|R^T�]=:�HW�������v�u��
�U_�:g��WS�Nj7~��ʤ<Ǜ�U*��q���^�_K����B�y���ʄ���n�9��Dܥ���3ݐ��l��i�q'�"sҭ�|0��ɴ=؇�F��>�S6�I��
U���"Ր�d����������ċy��Žsd��W?�f�K ��~�%|�\p��~@&�A��FV�[/&Uf��d��	�\ZJ�߬x�iK�멺=�ucQ�1�`�XB2{E0�9%N��e����s˔����ݒ�3ŉ�h��Sm�5��${iCu�3;ߣ��5�P��
k�lu�(� ���z�k��[��#DŚ�Z�o�T�E��0(�T���4���rh�A�DR�*�z�o��%��T�V��������<g�H�����{	9!�;�L8R��^<���P�ש}��u��r�ūQ��b�k(ƪ���y���� H�κ	i3 ��,z�%� z�߸�h㟏O$�5�����WP� 7��Ah�]��9������w�ג�x���@��<�&�1���Q2,���}�΀�`���O<�c�`�S�L �8�C�K�bF@���T4�Սr��E3Wv����_�c�s�Hs����Ry��#�B��� �.����M dJ,Ao��������*Ïi�Ɖ5x*!����ǣ�_T�k:����Ar ���t�LJ�K!l5�<�꼞,R2��bM�*��U2�@sS�3����u���Vn*ղkPz�'=���X��c���<)'��l�6�z{�-!�����<_hAʲ� ?~3�}{},�!'u��iUxX�<��W������O�������E�H��Ng�{�l�܊��(�� �llV�q�tb�E���@���-�w�"i(��+M_o�K��j��1��gFZ��M�L,c�F:�V%����%Js�b$$��K����<ן��g��?���w�Ʊ*  E�ԣ��k�f��I;F�S�Ë����/��j��-�]m:�f ��K=v{�Q��"���i<�x��̩|6�D5(��OT!�Q��2�L��SB$q/#�J is�kR�򩤘���M�Q*ƸX���e���M��`�LY�_�����p���T)��k�y!X*�N��~������ݗ�4B�lCb��^�Aa�s�+�R�ߥ�X;(C�-O��7e��6rBL�HD���Ӭ��c�H���Ͼ+%���hj�gN.,�??�BU&�=�����Է���+^�����ԍy����������P_�V����"Tw�K�>�P���u�
*2��Ճ���A�/���t$f?�g���_����q4b�_��Z\�	�D�ۻ2��̀�,�2��l~B�L�7n![LArP��:�V����~Z�EQ�Is�]c��1fAһ��Aja���*���{�9�/u&�B���f���=��>�ӮUx�B�N�`wX�8l�vR�lV>N���k�v�U^n 1�Ξ��H9а�uٓFn���������%<�A���D,d�ɏjH���$s�T��Xb8hŨ9���=�,X��p7�'֕n�k���d��8f�l�㬍�4�y����1�ޗ��I �^ӄX�qJ��1��^H5kw��ⷙ�4���X ���Oٳ�37G���'��nqW��Z��V�@�ћ��Hë�ޓ��HEF,�is�E<�0�J��`"��&�v�~�`]̰��E�3��Fݑ��O���q�6܊�/dI-���é��k�����R}(C��ag��,?r�����h����m�VEQe��2�{[�O��|��Q��o�J�#��� ��)�	G�#�e�U�>���b���CZ���'a��\���z��c'��m�yg�n{%-!���SY��Dx�j>|�m�H�|�}��նLT�v|Ng+f�6X������&�Cm�Mo@�%�}|엷Y��&q��a�Y�>;$b�4�Γ(�ʗxN���B�[�f���'sZ�_��VOA�G�2��]���+]��Z�WY~k�AW�[�,��2,%~��D��n���f
Κ�v���;�o��*(>]�R��Aq��:�C*��$�DۗU�.����+n `Kh�iܮe*����c�������H�̇�g.�wls����a��ube\ ����R��4��a�XVΨ��Z2��mh����:s��W�Q��5��XM��C]m��_|q�?p������6�f�0#�Ҽ�eT���X��@�()Rϝ�?!���^��*J���ޭ�R-�谺�&ӳW��#xS��v�E���p����eB%ғ�,��\T��;k�} �V|��\��/P�k��˶F�_k�֟�ۇ��M:o���~�t�D��.<�:[����h�LNķ7����I����r�d,�ϰᆯC��KP���C����,���}����7��t/k����i>ej˭4)��ࣕ���d�5��t��l�DX���J�~f����-f�NG�ir
 ���'8�۠+�#��z�M���_���!D]�����k;�v�xH�*�Ϩ�I�92,Y��6�'�ǎJf?������e��%����sU�C���ķ-+֖L�E�q�����TyL���U:+�Zxɺ)����Me�DnȻ��v�tkl-�*����3��Y0 �!rRs�?�!9t��K�sR ���1u`,���W۪�X���A�+����>կ��"��A����RBU
C�B��=ϺdcMx"��"��{88DH�D(��i��;޹��-�&�?J���I?����8��9H�<�>��!n��ac�L����}uZ��
# s��p��	)�M�#+!K�*�p4���k	�䊮�T�3�F��|����������.x�TNd7�{�*Ry�>��Z��K�����&�� e�@i1�V+ܘ)���+"tU�1�trB��r��t�^D��������L&�n�Q_r�^T��,�o��Q���b�>8Aȗ�����:�Y��bV�r{��b3��(p�����p�+�v��G�~��/��W�'�q���.ا�A�N��N��;7=�7�CC�2����T;N�t6��X�� Gi�!��YVAа !#b:�}L��¹|`�O9='�ؘ�� RF�2�J=Rw��3����	�&�����D�1d���D��)��;��`̘�o>�	Qn���\�L�`Hm'�x�3��U��
��/��3o��.�E�O�����c�b����Q�	{�V��#o���Sl�ŕ��{�q#���$�\�46s���>��7I���g�T;-�CLS��I�O����b=�B?� h�,%z"������%B���c��[��=�8����� #�E'y)Q;�K�# �MJ���g&���gB���p�e�Ў2�T&p��>R�̘ /rԌyj���z��|'8���2b�mZa{���K�*�'��j�ߘ̑����� U/6Y�f�F՜�U��@R;<�t�{q��ov�o=���w��q)�k/�b��DDQ�ѣ���v���b�^�a�j�C��gDG�_�i��
���*S�Ȥ���??GyX��k.����`�+�(W�Y���$}����\,ҏM^O���a��G�c�MH4Pt�q��\Jd���c��P�0��ܬ�<<EM��˥����F�z�,��k�
��F}0��ܪ�(�Ǘ��\��⦎.���
�E�c�8\��z)�xڿ���kެ��ka'�`�;�����T�,��Wy�2 ���h����{5ɹ�oP��������'`M�`{i{�D�R����H�0��v���X�x�>Q*��~�4��d^��*�N���f3�N�d���W#�1�ylK-���4��l3��t�%���&����ccLb
[�	K#\m|d��@��A�/x�\3�^[�P}��s����tWw��)��U��ǳ˯P�@��ΦP��;E)8&s���\$��E�k�Q�P����0�_))a%�ԡ��b�ytJ�oLo��gI������}�0˘��~�.����d��Wm(&��l髤[.����"2K��v��p���uޝ�fj9m]X����6k���B":�
�[[a��Ũ'�j����8EU	r}hj���A���$��?}�ӕ-�'�>��՚D�]b�O5��2��.S�����j�[z�g��`�V6 Z.�t!�V!�$�eZ��)N#��p�^ )�� ��P'm�@/�e~��6K�Ĵ���mV����cҏ��Ʒ�Rs����f��(�P��w-���>�0�fem:�� sa�%�/�6�]n�	�'3�g�UQڳ*�-�3��IWk�i��ˠ��rh�򙬅�䊌�Բ�/�,@,�Cc���I��U�{�A�c?m�ح��ʎ�;�ԅ]"�=s���k�R��WZ���@%�0fO��!9o�e�]�اG_N��[W��k0��
��|�Ȳ�-�i�@G�C
����%�,DP~��<Y?�TPz�j�IVn��ܥw�bo˶���@����M�~r�n��̈�&j7Pb!�.�
�tk���
<�M��^���M��!�/�r 1a�ȝ�p{�1M/3��|� 6cƥ%5쇨
!I��#�V�*��V�*>�/���b��~i�X������p�Z��*�R�Z(��]��0FvX�,��ϭl��>+3�}���xyqc����B繒~N�?�IW#ń��;�dB�e���Ҏ�м���f�&%9o&H��J/f�%�)웰�LC4���B��r%[�|F��F�)���`�]���B�Os|n��_�2�)��a��?��i��F�hI��o&�+e���z�%���"�k�<�@�H�Ox�������[O��H���4�46R��_�i�������{�D���3۞��Kc��z���F#ͼf}�yR#�6�������f������v��rB�̋������E��f2z�����f�w�¢�K��C4PSf�_�X�P�Rm�*���G@�PT���>�*��
�Ox1�Ӟ�64�%f��� ,<�d�:ʩ���b���c�+�	��]�*�g�������W8����&�'��B�V ��x�~�Q/���ݲD�l���!�~���o��	�}��h^�l/a�k�~�Nwq`��S-V��a�<�������|�����f�#�Ԟ=u8�t����89�K���
����r������gp�Z��lݎ��:��̙d��\����a��]��+�7���Mg2_/����F��e ��?b1��q"6����7��w庘LFJ	��5G��#�SY�2&���
�)�w�6�c؎���x5��yh��7��V׆��Qc�uu�j9��ap�+�d��QL��Hbo�	�*ִ��m��MՖ����_���2I*K��N���CJ�	]�Ka��Ȇ	��b�=����A�<*�H�of+q׹�ObE�g��!���{��?�5�)�I��l[���\Ԭg7~q�Y5��'ntK�&�P��]��8��W�x7-��R�!\�� ���V'�@��ю�"���B&~�(@�L��KA�2�r/?(�8"#��>E��5MLZ~�0嗺SY��|[ɰ��0���a�Ub���G���7U]|���*<G�{����![�����uk�.�.�%UcW�繱+I#��������[Q���9��0��)�_���̚��yi��gV85�[h��hL����$���T��t����61�ҙ/Z�,�l�ǉ�(F9��(ChS'H���5/:Ps�@0=c%(y�IgC�8��u��B���V*����ƒ�z��y�uº���+�"�M�1w�fH"U�A&}��Ս��G{�3[��Ц���ǭ�&S�D�� a{X��dV!�pJI�UK2�d��X�nؠb��^-��~O�Ι��g�t,�L����ޕ�z-�p�Yp���X��~��Zr�K�;��t@��QӞ�҆��Ds�C�� U��@���t2�5j�}i{5��˾�F�ݰ�?G1nE7f?F�$�p�����L��[ZN�+ ��#¨\���pta�d��h6����e��9�.M_&f�SP�?9g�w�r��̈́7��u�1���L���"�'u�O'�j��K�C��r3D<��z��z%���-{��&�:XU���3�w�p8�����G�3�6	��w�
w���3��Z�/ϝ@��t <�7SI��	@SK1��@�?�[�HU>o�c���M�_�p����׻w�U���)�\.#�Z+����4���ʋMy<a<V|��� ��
�9l�_��O�@�/���~�z�P%���[�����:��L'&�0���i4Hk�u����B�X;��)Vn�5բ ���;Y/�^yS�K�A�s�_���v�PR�'x���d�(��4�B���i�GͰ+AS*F�g­#c�|muL`��و�i^��.����S�g����]��s���F?Z4��J%�����	����k���"�Y�O�mj|�OP7���"�W�kuc#����0�~�����~0�xf��Ԝ�1�.���4�D	o�����
Pl���I����$)��}�F��ML�����B;��I��dT6�a�g��'�y�	��'}�p>��j�@�l�����ʗp�1��_"�d�1���12ɼ��(�"�.F/���\*�W��CӑW�H�Y��A�a­r��>:6^!^�D��e:� ���}y���/n(�B��oҪ�s5�Jn+Hv9`x�Jp �w�T�W�0T�[1��"�������y6:fa�S�[J�ao�tJ��G얁s����Q�$los�o��m<��U��g���w@�~s
x^�8+�����"�x+�]z}G�
O�g�z �:�����i�*��)�SM�ͺg��]f��bع�4�}1HM\�f+� �������-�BcG,e-E ��1L��-ϐFxI���۬\���!a�#�'>����SU��R�~&S��S��ߧ+�t�C%�_+���e+�������o��WN>��xM:���a4j�<�D�	z �)3PZ����f*/-j�2�b��QL\t ��dd�m��sFk�i�˾П7ۜ�&��i����ʛQh��{��6LU�����XI`���\CZ	4b���*��d��HJpC��ĮD�?G���8Ω﮶��������j�b&�}$�ͯ��9��z�0�
�q��,�%�[�V��1�B�gЍ�O�8Hc��Ey��Wc��Si7���^O���v�(��1~ä�.?iM���^���� 5ր\��<	�ȫ�߅�	Tb�˸G&�l�7ح����"�W�Vy͛��Na�Վ�%��`�(����`2�����5�RL̵�f�2D(�N@�%���s)���"�V�	�}`!<U6��-@���{s~�0�KK�:�������zy�����*�Z:� �}�Q��`tIa��ε �&��UG��i������z�I�5B�Eh�`�I��'3������
���0��}:%�o��P5��u_ӧH�|�/MH�����(P�	��S�M�@X��4�Sf�#r��� LbG�ܒ�/}E����ә��|��nL�8��Tu�Gy��3I!-�s 㲂��G�d�����J���F��y���Zf�]�I���ؙ���;���*�i@������G�'���C�2���Q�D�ʶ�'T�p���с�;08w�9���歕�m]����ݝ��{����q�:�K��$�nF^�9?#��TfP|�A�Ϣ�KR�y�`*��ʓ���|^����O��6��19����[_�gF�]�
�������^�el	?��l8R���eK��B�>XF)�Ub98�	�k����S�)s�%�8��')�����+���[�=� %"L;�}��$�4�CQ�،\��J���#��O�A�+j�w���<�ற�vV��O(ߌ�闉=�����ՅSwl�@K��o�y@����?�.~ۺ�Y�^���̼2�AZ������=�-'KR(�*��ah����E���3�Ҏ,�ҲW%��I�a"7��3k�]��Ea�
�Q�����g�;��&By��#f�.��5��~,i�=�u�_Q� !zL�$�th{�|P����1X-t�:�gU��y46��w��G�W2�V���c#Y�lC�
�y6o�xXh���o���<���}��`Bм癫��E�+�#*o#=m�{���>Z����C��Wm��~'O#f���� �s�W����M���<Ԟ͛�4i
�6�v[<l�+�\�.���9��c��������$t�	ށ��7�q�C��+O�2��.��R]����X.�S��[�a�0���sޟ�K��O�&���L5Gs��7?�Y���6���<"�C�/qj��k��� "����9��v����o>���5A�R]�%�2�Ν �������������̦USSxB�.R�
BA�{y���P��=�^�hϱ8�\6�#��z\���(���������0v"S���_e�����J �k�T���p�s��rΑ9��E����,:�U{7���mA��R�h#����l�O�8��T���d2���>�Pr����N�
+�T�12�]�V\U���2R�d���tAa�d���[j�q��<�vGPuC�<���E�9��9����HZ�I�b�J�m�W��ϭ�mE��,��V�����D&�ȶ�!��Fa%����t��t��w���(�=��ͺ8@ F�]7�w�g�i&�j���s�T���5C��fŌ�G���9.#�E�%1�A�-�]�i/�T.o({rM1�?e���ĺ-u��OT�%���1�Fi����"{@QZ��<ƃ�0 � Q-<T�$�����Jk�0�仮�Vg!�<�X-������:tnzt�<��6�3�Z�u��p|9�+$��������l�MS����4,��S�ā���4�����`�$rg�i=bA5�7�\N�-�[R"����W'"�y ��kJI��s�����!�@�H�K�k��510 ��%P݅���V�f�Y��K�m|�W���/h`P�I ڦ�f�.�`]Y<?b�<��?��^?��L��e����3'_5��hd�\��ԩ��X�T�:��֍U&��Υ���s�4�����'3IA�[��F��Q6�M'>D>$߮�n����=��^������^[Ɗl������c�AW��u[��u)ʅpϾ[�ך9뒜��n�/��������=k�a�/���i}�B���u9�����1���i���^s�|��`��y�U\� i ��UE/J��
]<�;���Kh�� `����֏&}�F���ʾ|�:�]D4/g(�TD<k�~&���P���K&��s��� ��'@=6����V����yc{��`���n���Kt����_oFڨ� ��[A�8{�0��x�+�'k��ʉ�ZKRB�2�&�Q=�0�������=�o�d�����N�����?�&LtQI�G��ƴV��	ڈ;��s�-�=-���	����1l�5�[���jέ��m�� ����y�:�X�;)��]49�C�Oz�ҏ�[�Q��FI ��$��~��j��G�`�UQ�Mv���M.���.u���{���(�o����-���[���87``�j�i��r��}���H+�����Kh�B���`ž�9�g{�gs�C�*�d֗x��
F1��RD����Np�ɇ�mf��0���	əAQ�m��om����p}������ń&�bɧ|�@*���C&������Gb8BUT��̵��Փi0]�d�V�Jܩ�h��e�H)lO!���#���%"Hȗ�^������U�J�y�]�8��a�ѮhQ�C���E(C8��-��Z��R������Vם�k�����.Q��u�}ÀOd^UE��N����d���CA��"�m�f�@��u#�����d��&3bF_�]}������(r�H����گ���N�s�f�g4UM*S=��M�TS��Q���.�`<�!�ܼUi�s��6���W�Z1v�<$�R]�� �'>:��Ff��2����:�V[���� �@��c�*��Dl�-*X�|�5��R��?-b��/��@EROF�ۦ�k�΋�[����=��s5B9L(\�K�KU;����Ϙ�����"C22T#6�U~9T���'��"܂㤍�4zϧ\9@ntl- #)��T�j�2ݐ�n��PV���f�ʋU5�y�g���$�w7�ICK@n0�_ܿ"}���������W�=A���S�_7�'^��-&��G� ��	��"	��{�7�����������~f�1�?{@�Q0~W$��Cz�k�efHV�4�P�H	߶]z*��0����nM&'3��X#XI�p�wda�ճ%1P���o"�cN�c�W
���G�

{�>{�S�0�(���|V�y�$Oq�U������L����Y~:.l�w�MMր�
��,�Ӱ�����ޝ1�n6{2�$��Kף�e cR���8��j�ȍ�����UF��D�	�q�YM�At��w\w��z�Z�4�/���!P��_�¹Ő%�gչ�h%�~��!Y&�����$3���0{P󫂼�m�j��)�t�i��T~����M$�}?�T��ӡ���и&>�\[��V��غ֟�(g�ǍU�ik��KI
[�v�	�guK�8�n���Z6'�$DK	X�e3I�x�ݒ1���V*�9�Y�wT�*���!EĿ*���<a?$6Cn�-T�rۂ������=n��R-��D�Oh`;�=K,�[?����w�w!����>.h�����ٚ�;#hr�:�c�/Uj߃1&�ӷ��B���l��@�XО�i%�/�േ�j��x��b@	k����(��o<�8�Q@�MR������H�����C��6���}%OhA��3z���MUz��o���Cs��¦��1X��.C��Ye �"�~J�b�^ =�V�$�%`m����@�/hS���$χ��R݌T�.��ƍ��N�u�C���}i?���-��^�M_h�f��r�,�����bϰ�,�2�J�G>�O�C&­a�� rU39�<|���lp�(r�y����+�DQY��)YR���e/�yG̽��Qub��<�:J�!�M,<�\@ـN�-Ћ1K��_�-�j�^�W*m��^�ͳ�"�/'|Mwn�GtuA�Y�Nt���T���G�lh�b8Ӱ�7ҹMQ1ķ���un7tW]���=d�ng`*�:]ʼ�d�H/a���{���P�+�#��``V��蛈	W{�@��.�������d�:�m$��\d��eT��<�?֖����A:��$h���3�!"��NG��zo"Ԫ��`��tU�&ヺ����L�%�����`�|�&�8e�	����A���\����q���f����~'	ꖂ�+�H�  �/�Q��rd(&	!r�s�k�k������`�AFn����xH�L� ��j@kIT��rr�.����DG�K"��La��0�~jb��D��~��'��8Ҥona���b�Ǹ�T7�r��}�<C��7��Ј-��7=�pY�ً�b����՛ ݚ�Rg�~����V�VyrW�+�G�ȌME���td�R�����K}X����i�������ݩ�T��'���� ȳ.l�[P*��󿢭C]l�<�8Q�PQ��;��m��S!����y����l��������r������:���2�du��@O�s�q�n�`Л��[�
��d,_ma�����_o������-�#
1#����5������Wæ"x�n
��Jr��c]Ta��!K�}����$�w�����׸�0O���a�U{*��Ѹ��7�H��P�QG�Z��&b�:��AD-��!��4�(	�����T&jA~�!�V��ǌ��g��.6�m���T5�v���=vzt�\�p����yH�SUّ��U�_O����͛޾��+��$��J�Cl�s?�����[
����B��T�Dq����\p�8;@7��\�Թjp�||j� ��7�iS��X`���-�o���V'I�g
�]�8&�7�����<�;�6ÃJ�`��MKU������#�Mi$){Ҟ��D.z�i�L�L`W�kE��)��{e��I�v.r��o���+��a�m�����ck5�ف�Ϫӕ}��D��H�x�h;l�W�j,u�\�Nq%L���<2u�*k�ѕ�zیYWW&9�_t���aHm-�N7c ��P-�wݮj�g��������`�����Qc�C��ͺl��x+փ*�X���yR镻�!G��hH˪��~ l��T}�>�Mf̠ ����<T��V�aD����]�5����W���x�h<�W5��Z���5{�\LQ;\.DW�	��6|[.��K��l@�	��X��е���:��l�5�f� �j�D���t.~I"J?�á3i�x��E��]<���a�6���p�	���6G��?Q�m�Z=gJ���
��!4$���X-�Ačl����rM��¢(;a�&�	b�u��/(rT�7��kb�o�V
;�R�x�=���ךE�E�=����ɐ|��lh�3��ґ�.���Ls骁�gl�����;� �w������ne9b��2k��-ۋ�<��C*�;8Gk5�����Ik��m�PX��ԩ��o��D�WjQS��
�$�3]����MIq\U�iv���DGS��TT����� ���	%�$V`���)�%7/�0�* �g>@����|R��fM� 5c���1�1t����9����><B�w)~�����nwR1t�A����畤���=V4~�"��2P�Mfޓ�H�'T]+a�_&I
��9�����Xh�縮Q��G���@t$n�Y��"c��ˣq!+�e��}�*��Ε��	i�3Lfź�x TS��	���O�GR;+M����yo`��=v����ļ@#ͨq�F�9R@"A�+��պ]ڛ�J�0�}떅U�tм� �� ��9�����d*�,��H���t������::>�$CF��#9����F!zq��S���?2%"� ֛~݌��H�K��X��BlC���������˦P��> ��,N�/�G���r歬��(�T�݁�z�"w�po\`n�8݉HUK8�+*�]k��zx��3yË�������<��W_��~��ۼ��Hv���W�ǌn_f&�8�O�+w~!뜸�/⍓�n�1�+���#<�q �j��%��U�9�/�H���J05��k�Ryț-0�]�D���� �Q���;��6٪�E�s���¾y2��Oޛ!�q�?��;�q�F�!�f�9���\Sx�3ޤ2�r�}�3+k�e�W��w	N��E%�����f�̂;c�6;	�NG�׊�ڪ���(瘤j;��_��A&w(9S��zK�)�[�/��n�y������R�U���<�`�c2�^Y�����5ߨw��]�	���	���%��5�{��P2�=���!�k"C+6곷���Un�'�~#�9�7OL9dZ����+�Т;�����WòB����^��n���	;�e�E����VS�����X�3JM��k6��p��(Jx��� �uL�^�3,��&�Vp7�3hͅI�R�|�{J(�Mn���92d�(8M��(��Y�A鼭�pr�g�e�O���2��T\��ܪh	��~Q�D�&cG�W�=oq�	���Il��\�Ov��@+�c���*��S��/���B�,�5shga,���7߮S;Y�����P�b��fT�ieC�b��'����A5HYU�?:�$�����rWfZC)�fY k�V�4]c�K�L	6d���w9dc6@��o�����L(߃M�wPe�7���撀X��ġ����L�˒�E??��Le>�`�ꄅ�ϲ����B�T�2C�v�M��@�G?U������������o�t��ⲱ��<��Ku�Ŝ~q��$�E�e��RL�d���T���Y�\l�	8�0eں�#�WT�nr-I>|d9��\RJ{U�M�Cė�_L��ￇMo�:�.��� I���4��z�w�.R��ͯ��Xf-���4� ��C�2^!��O��!�|�?�gMj�Y���$Hm���H8H�E��)D?8��D/�EE��)�P�@�:}���o����'T��{���3D���	|�qqG�3\Z�1�S}PfM�S3-�x�����^��Ě�O ���8��iGE�i�^g�_�F����'��*�^�8`��+T-{���(nˡ��g	�@�������k��'%����{�NlC8�������Y�����x`r8|q��DF�a�E���@��Dq~��5l�0�I��X�9<H"����h��CB��ؚ�/T8����"s�K�»��_^�.��K-����&q:!�@�i��5P�<���M����.�g|}ș]�<��VD������Jܸ�l���d:
�>;.l�W+/Ȃ��D��W]�U��QH�u�� enJ��(S�L?�@�գ�>����H>���8��BZ�J�;�ץ��-R�;�m]��T��d�hm�n.$N&��z�<�Y1�'��vԀ�VN�c����x�yWi��ѻ#�?��6��!��$���/�Ű2ԫ��Y� �*G,�d�r۶D�` �T7���b��{�\�s���i��͓�J���)!�o>��Z5�C�-���c�n�����,�[Ö��E}w_�TY�<3$[x�Wl��J�� 7AG�щ�1.���*��8�j������MyBP֛R5ܞ��nĖ�;�9:�,A��-i_��O���=�(+���'ZR�{1/s��e�b�N���У��.�Ŗbgڋ0�Ioz����{i��%L��3%^����A: i!I��ެD�5�OPCo�c=��[J���^�u
�xa�T��oY&�����B =��2��:�������WxO���7��n�e.{�*��*_�:�)�#g�� l)��lw�'[5"�\E��,,�
.g�=>�O��j�߉��	{\زQ���;�}��֓b�EU�.! Up�6�2�m��/��rk7"�~/u�o�J�;�e��<���%����àlzU�3�W"-E_��/����5A�/���$cҁ��ּ��*�e%��9�$~Y`k��A:C��(3�8U����\GkWU�ԇo���������@O�(��~��]��v�j��\��L�RY��V�^�{;��o�'aj�)]�e�c4�Ed�����ǲ�ݮkz�z��2��E��N?t�M(�{����3֓ҝ�� Ϩ�3H�8x�Ȕ�F�Q5N������,kS�i��U��u�u]��G�`����*�tk��\��2hL͔��@&�y��8�0y��QK�x��Mq��W�!���T,��ebv���֞�x���n���E��먱T���v�*�ђcg�S�u�d�X��ȩ�AKKc��x鍕��
�y�H�,�m����e0�����zR��<��:�u{n:ۓ����s�P����1�~�F�s��Dg�:d��֡�cK�Ob�Z��m_x���UA�j/U5�\8K��-����#��;�UoƦ>����6��v~�_n��OU��<����3%Z���,��.�6�f���K|��{� �p�-�c� ����w���x�M��p[�a?���Rv·�R��rj��v�'p�LK�*U:Ι���}��v���1���T�f&��[�O�mT�-ր�<2��s%2��|�y9*0����(~�0��!{�d����Ce�E�$��ңv�6z�A&�Q��I)�;QT��D,?>������� q�g+�Ѳcvr�-��j��V���)�e���T�;��KN�7˱7�L��;�{��h[F�`�Ud>e8�uJׁ��EF����=�-�߷�[�0G��}�cpa��y0m7#��(�{�e��[|��AN�w�zH�ڕ��0+�2\s�,��*�� �!,'oE53!Z0�f��d����č:���m��N ��U��<B�5UqU�N�~l; �r� ��r�BLQ��*]1Բxѭ��"��x7ywAz=姻B�H�T:r;���n[�8�#��LIJډ�g��gx.a��~�!Xؑ�8T�����U�I�D��$���,��:����;N��MZQo~�R�]�<���UJ��il�5��[�U"���n%�m��e`�������B�LMk��H�� ��pI�����!G�$���Ƽӭ�%D�փ%����?�`X	���xp�͉�J���IY��5Ăv�QC`�Y��f��	�Q�\pd%aE�6,z�������+��#[U䏅<�+O���v�����Y�joHX��D�5�xZ�_�Ô	�l�v��k��@(��8;ۙ��z�J�[�cnJ�)Gܸ)�
�Ln.RZIP��2��	�.A"`������!u��YP�#X�l�O+kXv_mr��{����M���aW&x�Z�D�X�d�l�����ߩ#L�τiPڼ+}h�~�X��f��mC<����Z�
�Uhɑ�Z�������!�\��u:�W���V����.�G�Q�)�-��4�/O�Q�Ӎ��d){���zxս��h�_l��6E�Ob}�4¢!�=	���x��ʎ�B�0l��rcSR��R�	�_z���^h��g����\1at*y�!ar�$�� Jp��t�*S������b��Lf�����/�k��d99b�)l2B�r�P-q���
�v5�� ;1?�j*��I����<%�?7��C`�g����9"��E �:��p�u.�Y�"��!�~�$XA]]ކ�i��,W�Ć�Kޒ���+l7%x1��m���t��<��n&�å���\]�I����y2���%�g���*�M�<62C��P��x�]�b�s
cF���cD������3'*�k�ƴ24iJ_�D:�F69�v=�ɮq�+�	1,?.����x��8��A��@Y�z"ͱ�_7}0v�Mzh����A;�J������OpG����HȐ��W,��������r��i��ޡ1w��0ī֨�@8�O��f�\6�o��9�
�yŜi`=�HD����v1oo4E��2!.?�`p�2\�>6	��9�J&�ۙ�Y��+�Ƒr��b�h؛#��v�d��Od�2e�j���r�Q���>aS ��)r��/�of�� ����KP�I�S�=� )8�xh(�`di�K�~Z{_��^V?�qԜ�:k���+�x�mX�Y.ı��H����F ����6ڋ�"�[���3y��q��U��v��uӽ9��$���=/��V���C�r���p���&M7�"ۦ�d������WQ�Fg��?���O�1q����F[햄�^�����r�|G2�M����N�g�
��0�p8���c1�Z7T�HY��if�w�_�P��k^4��B �"�lV���g���ħn�d��"�(�+�RUF���e���Dfổ��?hTL��<��?���b=*�,>��a���4P1��8.��ZW�����"�n��>4�y��Nl	"�k��賡>ٲC9����πm*-��)Y�鲇U{`�Z(�vs�ƭ*���c�~��r�[�Ts�܍��7���f�De����x�`��U��@�in���G�� |���%L?f�4](��{�ӥ��z����g\]��������1��"��n��v��:V�$%Y1ߓ	H�7��8�|�dF뗖��ANI��rNv�ݳ�4J�|��߲��@t��a`y�|�߮?��@t�5�s��2�l]É�8�-�I�Ze>�Z�\aN�m�$#������-i�%э�d�ϛu����'7�B��[z�uT�0�Pk��bXp��L'-���lS�k)!m����H����٤򉀙��W�<rʘ~[]�m]6��0�����E� � �z=2�� "�\����!g�YjE޼\3V��K?O���hs�1;���[,!����:F/P�_j�����ڟ�(bD�t�}��?\������Z4�c��[��E� ��G�6�Ng����N�n�+E5cg*�F�T�bTQ2s4���l�� �VY���y��m��p�s�{}�1�tg��h7�oZ/3Hj<�f��]�6Q�$���\��j)�� ��PX���/�G?��^(�� ������	ڒ����@�;�O~)�#�(8L�v[��ȩl;���"�b�n�ԏR������g�c�����RD�'3[�ESA��!b�����yD����\Ʈ���_��\�)*q|&���Ⱥyo�f³�V�qƳ��t�7�W����CbU>��5l�+�� �$��"�س��#7�?N��D}c�)׺�ID�#pu#\>ܩLؽjMI���#��������
qŁF�2�j��9ⰰ[a�����t^G�k��bg�8$�';�I�yd"V�dl�3t�е��b�q��I�����>�m�E~��_/�	%���H��}qc�����I���Fa	'��$�+�,c��Ò�woaԭGn�\(@0������"6�Op�/*���Y��S���`����\���e*��JTmx����~��-N���(!l���|�Yߚ�"�^�t����V����g�Ҿ/�V��RsQ^���İc�R�jW���Vd�S�.0��#)�[�"\S
"��p��I�$���O2K�}~
��t�h�z��j ���s/�����.}�z�y�Ua��Cm��=��3g��]��uC$	�-|���~ߺۦ�T!S;��J��K-�g�`��`V���G'���j�q,4G�WI;�p�a���v#2��Tq/ҧu�� �.�k�IZ.5U&�k�q��E�q}��`(�n��'��UY�z3	vjr���Vu^|2�����&�ߨ"�}P�w����}=%�]2\H��B�n�Ňӕ%��4$�fXS��{�rCà����X��y/8][��t���=k���؇|�ӛ�ay�f���gp�##Wu��v��?|�BZ���Oc�������a(ʫ�x�&�^�:�ek-1<Ů���/���nz+���cYֶք��FH���$+��w���J������>숺�OL��_4����q�]���?�ӗ��K���S�#������sVС���?����>;��>H���J\�!~��ś�7ׁ�p�-� �1S��I+��;o�\^ �TJc��h��
By�ώ;gO������S�Ҷ@N��&��`vC�����"���6J���jT��M��+Ngc�vS�`S�0�&�t�V�Y�Js�3>���u��Y��[����=�X����KRP�q�` �ȅ���s�ȓ$�>v� ����3Z\@��;�;�E{O�5���8�͖r6��B4J��݄�����V.S$�dd$�^Yf\B���l1�> ����{��"8j}����n�\t�����{l�]��.(G�A�w��j0W�b���Q������D�?��h�fc�8z��$Eb��1#	�К	��-�1���k�5�*ms��u�����P�rW��eGV��6�[��+{��Dm��t��F�ٹ|$?<b��NxX2��@��~(������L�x�Mv�O���D;�ia�����Vxz��UP�=}Ҩg~*��7a�=�{���ڋ��4Ouޢ�y1ɞ�A*��s��jf�D�#�l�@�t�E�KP�l�b���]&W���ъ�t��q�V�X:�.Ƀ�@�2ƝB)rMz8)� ��)T�L|Q:�R����:ͿV��^&MlB'כ�D,�Q=�yG��k�R릳؇W[P�Gq��ӆAp<�/1J�M���k�Z@�c[*q�R)��RȊ'��̡`�2�QdT�Nk�R�#dh1#>�K�?���������;iQlҖ�$�p�-xO��e�$!�&��)t����qTxA}? ̮����|
NҾ��l�B5YW�y�`�z���gY,����I��G3d��jGX��\H�k��c�o��o�������a�Qz;�%4���ބ�Z &�&G����<{�2_�P�4�c���Y�X�N)�㜹��݆f�x�EBz��vncl�<5=�9�%£�jq�NL�t�ؠ���f�� E���Y?gf������g+v(�q���VL�5���5)�x��u��E�l���Q5��7�����4�-���z*�\��s��L��E˵���;R����g�z�(�X55�^c��cs�������L����tÌy6S�O#^���_86g$I��Ԣ��n��o�x&���b!:}.>�q�py�9�e�]ՈVۍF+��h�
�����]�st=�ݏ�f��{0W�(�8gc��O׵�������a'<.lL��r�C���r��x1r�	ќ ����Ţ�e�v�IHX@��I��vfN�.�A���	L���T�+<�!�k���KS_߼k���B���s<z2\c#Jѿ.���[����n.�Jg~�W?Z���|�`���d�e������7ʁ��s��%/�2�Uk�"
LދwCC�׉O;��ZF{u��D�������X��c���'��vT ��xU�޸����Ө����97�9Yy[E+�����ǟ3/ �Uνn�1\��Ң،��)ʖ ����{1Zٯ��H�gd�{����Հ!��y$P�gJf�0w��b�bɷo��$��v,}�㌝zNq��8�kzY-^��F�JA"i�����:.�٤�I����5����r�W�8=K�K,��<E��{~Tf^��ڋgW��(��De!�
���O*ڗy�*�O���G+m��q!�b�B0�)(U.�����	��}ϨƜ�t�F��쩃�����Y�I���RL��%�>\�Y�U�[5<L�Z�5�q~��c.��)N�RYRRme�����#?���A�י��rx��|BFN���Ѥ]�:�2(=!��xN�á�+}�]�sP�]���Sm��X��vd���mC�K,�a���I���[�R�!��ez��Fx,��:|����}6�;&�˃�w�j�����P�i-�i.R��.��4\3*����WA��C��H���>&dӆk����u0�zD��!t*�U��R�f�=+��^��n�9~ŧM��]�{dk%~�5&�	A���L�+T�{j�o,���8���bg했��P��mr[���(m��h�(�������0q!�ĝ��&�B�K���_["B�5���u�V��C�/9x-νx��Ԛ\�}�K�`qt���Oj��G�>���ݘ�/j��6�Xϫ��Kŝ��_�ld���zdgL��5A�`ce�@��ͣ	���A�W4�5	�6���U�kQ>��D�s�N���+;�E��W�{�H�\fĜ�i�JJ�¹l�3�T'��>_;#,`RQV��%��=jc3 IHF�ȹ��-d`��'6�|'�s��bW�TR�X��S��`�7eZ����ś�l�j�!���|�S��-�K"����l�,���c"�ؾ�T�/��u}5&�ٚ��I!2_l$^Ww��J��#�v3ۄ#��6�OP�T�P�I[!EUE14]�K���t���%P��!�_c�P{�M�0 ��ۺ�����ǁc"�m��R���xĴ�q {���R�{���H6�.�ҷ�6��ўiN�����W�H!S̋�5��3���Y��(�[�v�T�(n��36���Ƶ n�19�_,`��͇���9��+��%,�)�âħSl�h�
r�|�����#ӓZ�S"@�-f+�k����X
Ae@ɯ/���Ľ|���)W�g<cRߛ	S�0y(��x�@,�����ϩ��Aˎ3c�9�WG��?�7<�{3� U����-�t~""\�O�-)�KtD��?��-�ƾ��B�o��O�hP��d������� 7�����ð�7M�Gi���R��2=�ssz9�����ҌJ�lo|m]�^M[����ս���vX�琛:��� �tϡ�>iu�ͯ�V�w�s��g�mQ롶��*ȝ K>H���h�}����r<>\�[�:RfR��Q�jH!�p�T��v�
9F�
�iޓW�G���߬��}�1H/����}sƓ(O�X/����ri��1���ۑA�v����5����:�6�п8G�r��C<��Z%mI�絾��w.H�@Ҍ��l�c�x�#s���e���"�b�	��͎>XCЀ�[�g/�xfwЫ�z�mɓ �ލ�����/��*��F)!��	@!w.����1y�g��^ġ u�b��U��sl!K�We�y��Hᘭ��>t��Ωp�k5�&�K��� �����N/@T����	R��t�D�p��A[���BU��A�ϧrw�M�4� �e+~�aq;�'����1�z�`�O
�M�L��>C�Hu5�ֵS��%@u��( ��� )c+���	G)�`b��)���=H➼�7�V� ;5��Y_�H�L����ZS:˵8�s��i�쟠<�J-��I��'�֨�|�Iw�_Q9$i.͸��!A������
�󙾗
�Ţ�>9C�ө!�-�8=)ynyǬui~��(J+�7�'��O8y�/�:��Yڝ7֪�}�� Ü���Qj]���MH^��4�<1����I&�7���8%��}2���X렃���F�Z)���d~��+%���������z���/��@(�2��d�ղK�uCq�s��)E��.�7=��C���RŅ�]����i]�׏�Vp&]�8�9����U6�i�+�������(���8����)l��F?-Y��uT��2�o�Y�T ���ǧyZ��!��B�aY�`cH#PGi�*y�kV�	Ҟ�h��L��-�ڑ=6S���y������q��M��<�yXB2������t��d��lR��(������V�g�-198�4���T8���@%x�k�=�X�����H�� �6�*�f[*���ߎ�e�eQu�w���N���--#��ͼ}ȣN�b�Rg�rW�*@��h#�������E����Oi������jD��kۓ�L�=)�U�&��јgI$,P0  v}��y�1C���'�]���X��#��3Ʉx{�j{��uq�^��,R0k,Q��5t��+���)=�v�Y'��n>S�
{��D�C�xbU�Y�d�OlV�-����%=��? �)y�ck�ʹv��zZ�u?݄�pQ�j%сnQ��X*?����<W�t#Td�!u������J���:��cJg>EAM�cnhRyv	�}�d47g��1�\��{�w&������հ�?���7�e4D����	rCD!%�;�8�;�'� �C��O�)�4�&�{��q�*C��iJ�=|�s5�rAx�u4&�1&���@�'���Z����Z�Ϛ�Ȩ
V�����-9��j�J��x��_0�ɜ�_�}�VХcz2��%:�Z��<&���{Jw�+}:2�4��mz�^#:���#m(�<Ił�,T�~��Z�LE��l$:���g �U� 2���
3Qt�,��`���
�!��b�-���zٯ ?)s>��ԕx0��P(k�ZG��h��Bo]�����=D���̈O��,$3o>E8l�z��I�l�e�/���_�;%f�4?�uo8��TXr+ ���4� �U�ნ�𔴚��qn}���8��3�q|���
���|Gt�d����Q}-�:�<�������Fݣ��b)�s�5RLM�1s����Q?:��nb!�)�08�|N�~��6<� ��޾e�be[�8����H>D<�\��d2Ǎ�r�b�K��᎒y��k�>��UA���LRM�э���&c��LQ��2�Y�����1w���c �U���L�nL�.Xi�7��ca�ޫ<���@� S1�����c��?8zb�A�@v��/�5i��������oc���K\��:@�nA�atˤ\D�$��#ȵ�UL^��.�	�8.�������uX:j%\��e��)x��o�#/���k�Z�L�G'��ିP����[��,�6��؅Ҫ�ͪJ�+����Q.M�9��R`{E*���F��F2f��a��>�B�ߧ���P�� e���п'�$}�P"L�4��
��P�stP\�a�s6+\I�u���H}Y~��5"��D��ˠ1jTʭ[��Ek�Z�{GJ%�HE2�or(n	���/�È@k����b�U����򞚌U����oo�l >&J�N��׿�2u\���둇�Σ�U�s��E;j�(��*x�$c
�m�iڻ���ď�vv-W^���m9�=�������@��5���ւ�=��-(����P�>)��%�dG���:_�����:c�K�����N�E��r����\I<���ڨ��T!���!>݉	޺B�AH!���NXBA�L�)����d����S�gQ~�}~��
�/�$���@-_[|��~�טmWʬ��4�6N���[o=��,I��)Rl�܍�q���{G���'_mE�<� ԞRc��@�d�;hj�jO4��S�Q����GT��ԭm�wiiw��jz}mBT�����d�ʚT)(K�P�=���K$Ak=J7l�2L�wH�ÑN:��{wQJ4�BE�&Y�l���йd��@ue������︲�=���;������Ƶ����Oa��6�S�C����&�v����~��)6�|x�7"�(���'\�nM�M���!�]�7Reb5��	��L5=�+[�2� 8�fKɺ���`����aV�B��R�`l_�0"���8]E�-�ǵ���~�#\{���2�Z@w���iLRƭ_l�G�j�*s|K�.8-'OV�n+�L5��B	�������q*&�H��]��g�m�*�Sn,MaL�Iv�%.����cH�8RL~� �m��eX!�^N'�"1���"s�^���#2ݽ�%Ų,��^�S����C�y�V	C�M�@QQ&dJ96)["����@�{8�����*��$�q:�LD򬙡�T#�M}�0��w�E^\\'A �P��lH
�����թȴ6i}����St%1W��_;��)�Tbl�)��\�'KԄF�&D�z�pD[�����ԭ�_�Eh;=%}Į!�w=�괓n������ҨK��Xy\Ђ�΃��\�0�٨�1d0u\��bz�jL��h`�7�cb裓��e�j��f�x��l��bQ�CH����v4g'p��#Dg��(g�e0I��H�:���[0w�M���C�a��=3_Eɥ�=�U�u{m�50Fa� ����S�����Y��p��������>�J�г���{�U!{ꉅ��E��1� DV��<K�XЮA��$M��A�gG��N�@/����Nv�K���?3ى��ˮ�٣��x��쓐.�!�X7i�6J+3�{��C�n�!9�d�
��G.h���6|��e]{�Qk�9��ԥd�9���\��cR���>(��c���9d?\������	� c���c����q�H��l�� �5�p��g�h�"��z�/�&=`V����e�������M�"��đ�`3�!EQ¢S�˚أ?����6��+`-q���_�n!pi�OP=��+S�؃5�v���7�QV���|�[��x�k{2�<�pU8�E?qE����4VM�D�Y͊Si{`5W1��w%�w�C���s,�9��._Bk=Q������ìy��'qM4=�1>㇄Ө&�d��e�t�{��	�'�g5p���#ޢ�o]B2y=�e����ѷN+���1����3ǔ��1;��
���fD2L�o���<.9+5�R`��ޔB 1]�9]~��Q5�~P�J�y�e<@e�)"=������}|NK�P�ڡZ�ߴ<�gېG�M:l:�g��:j�W�ݵ��:t����9��͜�;i�� .��im\���;Ք�5��/�T�~�Pb Kz��C�7�^�a��l^��:Jex�Wc�����X�F@RÕ��i�!����1��3�P3�y3�{�<KE./�*��此/ȓj���h�HCt�YId��zy��	~G���Amm�8���u(/�B.W�Z�&Nj�?�U�T�G��z�&���x=g����ף�� �Q�G/��'�Ė�o�h#jNy �P�6Q	�j�k��4̘�|ʢ�Th��p���-�w ��� x�3��vB$�=.�H�2'r2h��ws��&�]���?5l�G�P�7$C��c;	"��?�c�rp�%$?(6��q���t>��U���"l�*�ح�oGD����e/�s��.��ݻ!&1�d�Ǡ�@�yt	����2�yҽ%��V�ց μ��}S�|E���KA�{�O��@<�P�Ax�`�?E�O�$��_2堠xM�E�Q��ϛ܁ن�U\J�͹b��t�
-�Mn�S}{0��VP\�T
]<�Cɨ�UE��H�֠!��\�]�g��V����ak��yFs�2)z��蝅9b�����ݖ^������'b�>	�L���se/p��o��hy�_ؤ��rD�Q�����)�%��+;����"hפ���6(U��3e�&/
 2���m˛$Qar�*^2y�Lc��tw{"G�
e�0�b�y����Q ��HR��.Ƨ�:��7B�B;H�(���������v�|u-�D9�x�+������a�9E�9Ȱ���$W���{�TП���܂fx�ĨT[T��]���_x�7?@0V��D�?�V��-]�V�zJ���ˮ�H��r�b ��"#����ਥu�}��T��'��/i�b$U���;�THx�e-�F���u��c�Mʒ�znq#�T�=g��z̾�h+t����vӝp^%.4��]{vz�%���W�H�P�9����k8`��8l�J��w��A�-w� �Nd��K���ig\e���#�Ă��I�����+|��ݭ��H��8�"$�A�5�ª�_P�<C�W�����hE��bd���L�x!�i� q%J�n�R���I�!b�}F�zʁ F�CĆ,[�L�!�a�$�2�JH���ʂ4�2�ޤ�e�ˏ
s�_����������G�ڠ��\��>���2j�N�����;O.�f�b�ѧuB	��1�>zg<��l��������0��>��C^`�iRJt��%����l���=�;���\�^
?���s���#b̼�p��p9�w� ��7��7��П��t�!:��\�֡�W��aGh�"����;d>4nz�b7djDk.b�ۗ����t��<��7��8�4�S@�����d�}�R��1>wf�����ߏd�� DN��}		B�g��r63�~�^�26t�&�<��W�	���ʶ���jn����=x��f��0�4�Ui�d[�o��a�iR���V�]3"7/��$:Hm��TO�M�7�t�f�Ri�g�_�u���av���������z��+Y�ܘ�X^~��N�K˓�v��ɺ��"N3ni�I����KJ+ps�<��;6F�zc�X�2k�P5ڮ5�B-�e?ȱ���.������H9A �>������%��iV���t���K�G�7����h�*�B��M�n�\��!���x��~��f�n�I���i:K$ơ;7g)�V5����PeBJ��QM>�s�v�Z�|$8)�١kF�m^�}9r�,aC��q�7�.Ϡ�Q�$�w)n P(�d����5/��Y�rPye=��f"�mm�Z3�c�tEsbP���Fʲ��7v æ7 S�*o��#�7)#_����4������0i[����v��WLP?e��8R����;(0��3��b����[�$��HP6�O���5c^-�&��4��Or�cN%�%@�_b���F[%5.����pC�
e�g(ϟ�sJc�_��cH������LLuD=k<ED�b�kz��k(`��%}��,'эԒ�K>�.&�*�?�-x��cB���+R}4 P��O*2-��$Z�������x������+�S���o+�j��X*Bst�M	�H��vd��h�E@(z?�nެd'��Ӎuz���s��O�޳~&a5M�"��h�j3�S�?j�S�n��n?��>��La�p��Y�ގ�����a��&W�-~�Yk���I���Z������0[ͮ���Ӻ.L���AX�>U�BCe�ܝdbh�3ڍU�(p��Q�ѶQ��R�
m,��a�x|��:�Dҽ�1Z&$��5��U�b�2#�Q���#`p�q��}��f/������¦�(����XA�R8�x-���Q�3IZ�e�r��@���ևD���kT|>�(q9Ρ$�g^����@̡�U��ڎ{�G�C��Gc�#m�l�,�����(�`��'kp����e�	�}�p�tN��#��|Q�[z�s� �e��멕C��M.�vhM�K�O�U�{A9#n��zO~Ǵ��z��D���$�5�u,�&㜫 ��[�ߐ���mf&�A���u�4�w�_��?�����A��u�s?�xJ�85��Ǽ���sL���d�=DZ$9�Lwa~'�q��]#�I��(:ط�ߟ�ϊV�h8����\��\�k0�l�ȉ��fOP�ӗ�(mV�M��#��� �G���Q�n���t~�ǭ�u�b��G�@�t��Q5kp�Qǂ��>��F��@���	�TQ�_ IJ�_ڃ��cH������y����R�a�hKwIF��G��8�C!&�=�7�ԟD~4��J`Ē+�y��k0"S�_|Lu��(Ƈ��S�k�:��t�TT�����ˮ�󢮽��*�Τ	����b�G�M�S�L�0v�_����x���������������iZ�D<3�v��F��LCa��so>;%�rT"��>�G���#	��I����VR�BsAã�k�\- H��mh�D��.�+Jݖ�@z+�. �ʌN$>Eg#\!L&���T8�x7����ږ�1H�������������'��~n��Z�'�aHk�k&��ԓ���Q���|�ۂ������=�卻�$Ź�BiFJ1��E�7l8����z�t4�:;�dT*�z9ŠWG�j�NM���]�N�,�1��,b�}�w˃�ڴ��jaޭ2��DD4�4��"Ӑ�r��B��)h4�+�l�h6��8$E���fd|@�7[�B�)>={>�U�����-*PT��aI$�ť-�V�>����&�I�&�I�!�y�ps�o�����Sx%��f���'�F��I�8v�}`%�����Bx�F'?5��Soi��r<�=�lM%�����Q����Z1��y��ؕ"_���&a���2n&�Q���F�����5g�֪��KH�n ��$Y���G~Y_j�f��ϑT��!e}	$By�9:��\p~���|2���ʿEByR �p��Sqg��*��@b�r�@��؝��6�*�z���,�E"4��+xG�΢�#9n�i��b`8������V�2X�Y(�Tդl����1^(��ؼ�,v�w�'�M�D����[/'gO�d�hf��:�C(2h#a�e��-������PQc~����lǑ��T�\]����݁�I����U�!�1�=�q\�jzG}�C]�3?��:^.(EW���,N�J��#�f'"o~u�[6XU�~�o�'�ɪ� -�,��C�n��7./�iQE�����t�b��?�^���A�{BL��W�F���ǟqk�.���]6x��
�K؛��Ӽ7��������E�Eх|�sq�0xi�tr&Z���cB��t���s�a�����.���r��6����ua��Sx�����]�_���Ýu�|�,F^���C$�C�����+�{}�2��֥`����m�[ޢ�.Sg�������U�����デH�I���%�~���MŸh��k諮��r��B�����E*e 8-����x�����������|Z*p:u��*D d��=W�c��s������┛������-,P������)��� �D�4�� ��븲
�"�z��S�.C4�m�a@�``�������S��-��7}R2L�� �6bA7~��DX�d�c�=���� �%�l*1[@~���Ð���CR���5��@N��Q��z.]B�#p��	f*���V���?w(�̷ҁ	曞VM�CM<V�� H�Neߪooy���frS�Xs��p���j��/8E����d�q(��c���\s�����WjT��e��5�������)�Y䈩ӏY������O�����y�?1G��-G��r�0�i�D�=��v�Z5�z���4x�c�Qgiv�e���r�`馗����:SP�25IWu¶�M��f���I栄>��8m��17(�izx}ua$�T���q��vΞvO����X`j5�F,����� t�P!'+Q�JnIx4���!e4��ޔ̰���V��^qc��xLiDE�Sx	bLq^�
�4V� ��I�\
GQw�8��/	j1���S�EPSTQ��tb��~㦉�5N�ٜ������4*o؁��q����h�k���+���LVo}*f���_&9R6��9��f��Ui����_��Fʷ?*����)]�G��""����ζl���i�05��ʇ�9�J9�M|�>�X�ؽ���F�� ǰJGL�ǤR\�W*ҩXB��E�P䗮:
����mq4L��̀s����s�Ʈ�A��� ��9�mt9�iu:�PpwH�R�8ۥ������힎:_a0����tI���r���p��A�Q-�Z�� �q��T���A�u���`F�yH?S<�&C��L�J4���/��ц��U�e�%���I��7Z���S���i?���PL��7#�\�Q�<;s����i�\�+PQ0�n��Q���h
0Qނ&ڈ+�|^E��L���;v��b��	�7��Xԟi9�g{������\a:7o�䌊�V�%|�����zF� ��P�%pry v�s9Z���i�M��z�쮑�{;l]�{;dK	/��Yk�PJ�<��Nڮ�]�_��6١�۫��¤�Y!������Ҙ! �7���Ѩι5�	���{(UG�!�2\�QW��f�$ŗҽq��7����`�Zn���5��,���Ej�w]���C'Թ�ч�"�h<�k���x`M'��Lə�#8���	OJ
�/���tEť7`�I%d~�mey�XFJc:�޸8 ��c0����s�!qP�%��J}$�8M�5��@3(7g��r:����ccn��h�4v��>�*�=�ie�2�n��ԍ���L�BX\C�ӏ�m;���������6�*�n��[�r�pv��39��=ܢL��6z1F�l�3� �^�	p�[j4l3�x��ɽ*T���Y���P�-s�~��lś�Ǭ��\k�W-�)~h��$��y�:t&B���-g�� �2è>
�T��&�c�k��A?�&����iж�A~��θ�¦/�k����^�Ĥ�)�@ʇ0w��$���	5�&U��gPs�d�>3��eē�e�-j�Dp��Zq���(K�����"�+է�y3{[J��5w�"�H�'#~<����X�9p)��p�K/��b,*�}�E�o`,r�Q���,�D�K2�̓�NŎ��	�ثe"�ʲ��cX�N
��;ē���pG� 	M6�(Y�;�����������u��0��4��'����C��a�ް|��k����"k�7pc
�x@J��G���IM���1�V)?�����p����Q�{�M=�GSAp��Q�����Ƶl��l�,V�I��[�-D�<
�tl�ok�>'<NWW��A�7�=���7�=��W�I�?y��B�J�OE2��os����J�sh��qX.���"�#�q��y_O��p��L�����=�B�T�K}��]�y�Mp�!�}��\����)viF_W�|����̜?@IВWD�њ�l���Șjr1XN\�d݌�����Q����I�$�L�r���ıE
pB�^_f�1��'�������I�~�³�����R܍GG���Є#Z�oR�ˮIk���2G�Y������l#bO��Xa�T�S���8���L�%�	�3k�Lr�^3��I��Q��;|��H�]�K ���d{�A�+�!T,t-."1,�������IW�J��ELݎ��.֐��;�R���z�iՒ�b�I���lC8�qR��T9�W,��Լ�A��Z&��
;.ڥ�u�U�rL�p(f>�DQBH�,�y�
9�Kfou��Q�j��1�I?���,�����s�v0��i��
�W��YJ�=�Ȼ��X�b�m�ThGj����#�HJu�2�L�jI(���ϒ�^��ynd�W]�F`=�����Qb�����9�]�7�Gզ���8�O/PE�����4�B�!�P!�S�f^�&rt	.�d�\s�[?�jY,"I�.$�򛲚��L:�h�g��vrM��!�}�I����e�j�<���Q�zܾV�FS��}^R���֛�E^�g�;ۘB�$|w1�Y�A��sɦ1y�-��&
^�}����&�κV�"C�<���3JL�~�"�Z��*���0�j����W�9����_��?A��?�1u�B����\�ǄF�L=�� �4�K�E��_x{K
?h��8K&EPb��W�E�E�^�����_=e3���i��Y��J�̋Q!��a2�����
�8�Nw�W5bkrA�?|lPċU�|��k��v0kL�BVҹ�����;T.���+Sl/�z�QD��
�-��Ι��o5��Ə�6���ID�#��F��,OW=2Uړ�������>Sa}"�lZ�t$���!c���enC��ƞ�Nֆة�D�^Q��^��P7`�?/��3c�x�y�����ۜCq�
����oZq�+�DC��Y�@Jt���|��3�hE�J"8<�K�w�������"�xJ�a՝��v���O
z�|�
��Jb�^��.�r;��f
!b�:�ʮ�=�������q�^�-{r���g����,���L:�m����*�s��5B���?��PO������O�ħCRz売P`�o�q��$�6?D�l�e�M)�QE@���q��Oն�=�'�+�O�c��q��J?�j�L��-G�����{�~���%P�&����m�b�5 �Q�Ja=N?�+4�<���˭��	I*�'�"O�}J���z^-���!��F�ң�lDF5}1�<��≲�[�HU<�[��:l��J�Bwz�D܋L��a�l&�og��F�W���2?up��w��;_����>rk$�����q�,�J>�����}F����`.��,����a=|*�����ȓA�Ԋ�yo
Zu�7q}9��)�`Ec`�c3�F[�B�/.aqx�h¡�rO$/������.B��n.�Y{h�цt�襯��W��4�\�חF�]�yl��r$
S/�%0~?�l�Nl�1��!�<|�2X��x����W용����eo�u��s�ӛQ��'37���r킁�^X�JJc�Qz5K��Ӊ��Wj��)a�Vt��{u+�9�	�+��AI�tIh��#{{�#��d^����%R¶� MMǜ�I���l�t�W�I���G��T�������߰�؋�� F�yװ��\i����|5�#F:(%��ۑ᷺��ۄ���>��>����tz�~g��a&���M*��/�
b�i{�%���n�N�S/"P�u���]^j���:f���u��KϽ��2
�B�9��n\*���W)��n5��Ʀu^$i�KwMf�\JK�s=B_�H�y;���zY�������X�B��Ө���'�m�b����p�\��m?�U�L5K�\f�c{}Z���Y|�H����]O�2:im;�VH+z�*����qğ�\p!�"����Q%>���,�ֽ��KP'M�:�V�G�����]�SF�F�o��C��7	�g��Y-�SG�z"��$A�*�.�:�fRF�5���6MA�]�>��Q<��؈��l0\�'�d���)��pD-�g �o#�6��"���f	u��0_�B5#i�go����C�5�[l0�,�D2�H�?㖮z�%!����0����#������o�誁Ѻ�^UPq(w���7�)Ӻ���s�|�B ��/�`�?4��+-`�;�a��;r���Qz���FE�(ݮ���D����S���[-�M��r&1��A������H1J��@�.TgC� �w �ᓚ���%	���;IS��	ٔ+��8�b��s:����Q���w&�y�����%n��1�
z�@�%USI�y�K/:@gM�����+-<d�S�}#������o�]#����+ZB�Ewe��N���b�<��N\#�c�uҮ��G��z��y��%��F3�r#Q�Pz�33s�;�QV:~M�7X�ǆ1�l��Fs'*=�j�O���U�n,L<�<p�y
�ׄ��n��ފ5�,`~����!�GNm��Īj0�������
uU�S��?� 0"�9z�3&��4�3�����b�$%����v{v��e�o�� �[�A��<����K�Q;_�!�		�fl��;��=�6�Ec��,����.ԅj�WR���~�ja���A4�bČ�Ce;4�uU�}�S�}~l�a$�&��7�	�FNۭ`�];Gb�O1Ш}�:I.��v(���,��j� ��$)�L�[K��F1�iz���d��	�3��&�W�ԉ��:K߆�l��黼O�(��Q�Z�IR���z2j�|��{j��4��&��9��{�i	�u7K��NJ���q�H!z�x��,�jͦ/�M��iS�c�L�K�=����I.iy))��r�N�e\xNW�\�7"�4Z�d�$�V凂�2����T��P�K�*��JGz�)�~W��(����a���
%�$G�V*XGR\�#f[��{��a�����I��6( ��X�%�N;2�e �XS< ��U;�D]+�����YS{��1b3+���y'�E��&��ߟ����w��D�,���M��������\�x��D�4���9�]C-�����
O�ci��y'g���oF�B#Z.�x0z�%��~Ê����>[W�%f4����́�)�Q����{�/8��f��V�	���S�yy�C	��(0h�b
��y��0>�}̔t�Q��c��F�C�;D4-�E��s!�'@�SPk*����_��1hz�'��5/��A>�oz�g�m)~����s3	S�6�нe�>ɥ�8>g��o7��C��+|�޸E����^Eq ����gX_���	���^�޳��B��-�w��K�>��'$�4�|PIӲ����d����~��V��+�x.��}~�R���,���D)��PJq�T����m9R��;`C�{�Cߟ��c��ͼz��?{"	������5��.c��u�AZa�{T���F����_%9�#]�V��(������j��*����:�|����m�~�A�?]e�����+��v�XO�D47������Cmb30�>i] 1LN�}P��F������Ћjc����N���hYN�)�n馜m�р�Bʨ��;�oU+Xx���s �{LU�$4�ޣt7 �J�&b�HT�������n��W�o,8� �{��u��!ډ�'���f�4�Ō��HP�����y^w�ko�m�$�@sdVo�T�"�fN�ER�L��|�ӵ�2rUђ��d/39~g�3��c�b=�3�<�܁���T,
���_�o��p<$�/!�����}���Rpi�*�8��@S5���C�<ʈ��%ݕ�D�	�0�P|�4��ّ�����S$[7��4��\�Lp��L��=�i�|a3�Aږ���ȯ�ǲL�ƕ�X�(M}�PL�HQ�с�>�Z 77w���s;�Tģ�(��f=>�D�=�t������<8�k��a<��(2��U~�B����h=ЏӅ$7Uc�Y
�^J��yVRPZ�"�|G��7fާ ���ٸxI�е���#�iPc�_^�N>"�E9���+���GR��T�!S?{d2(��=�v��\���4��~g���ƿ#�w����%�/c�=�}}�0~�u�a�z����+>�b���鴯Y�YCS)j��L^����
�t	��(�( l���͋5Ph�"����Kb�"kN��L��Ӏ"r�$�~��i��������!c�U�8��U�|����Pf����*9JM؂l��4}�궓Gs+�U�y��>I
��2�a�� $,�g&Wd�>�V�.��0��g�F�7t��"��3@�Ҽ)�/<wx�/��:9�-�y�&�>+�!*�#=UON.b<
^�|vg�ݝ�_�m^*d�������G�r^LUA���|�@��E�Y�5i�jXF�;�����սA}������4�F��eY�3=W�'&ݵ(�o3ޥ�@����։Q�"�%r�u[�������jq�ّ�4�+tv�1�:'H���
�x�ӆ!���'�DQy�y��v6�U�!xד�5�
dhC2�AN�X(�0�!����=3�d�ŗt9�dІ��U����RoeR��+��Jb���'G�Yx8�hF��-�VRԄ�O��X�8�E�Oh����$���q��j9p��bI��,q�����z���A����4�f�eX=��կ�;��4�*05�?��}/C:}�*Q��;W���CL2�[bi^�{w���T��߃(}�s`�h��z\Ƌ�9��M�l\��F���� g�Z$�Z7���1|j( ���8��$0zO� Kv�B�2^`���X��J`g3��+���|��W��5"�Q˷���c䑸��܈����2���VI��ߓ�N��p>���5w�'����|�R��}\Z>B��W�p�}5�g�O~�����pƭҐ�3�����>��i�ۉk~8�إ�8f����M�}�>}�2����}@_��iG�-0ѿ�z'�P�&�9�(T���4tlQ�N��ՠW:?�by���щs�(v���"V#20�a̝�ʊ1�D�Z��uJz ���9����A�@��6�q�����N
#Q���	C]��]�K	a6�i5�<~��U\G�N��mf7���zG`����%x����R�&Y���/��:!G�P-1�����}�_�Í��'��F)�3N1�2��o�p��5i4�ħ(,�Tv�Z�������M���ub?Udۯca�Ł���pN�&'�����F��#��	��\ò8�p�B��pif���ۡ ����y�lZ���u��O�����tA�csId�����W�m�� ��ֱ�	לGO��ɚ/5�Nm|�3�m<�G�H#�l�D�	<)̱�Q]{��6@��o��zՆ�N���V.�%PQ�}��J��l�_�2535\��^:�����w+Zf2ɡ���<��d����~�*���~6�㵢����+�S��M��F��?�Mt��#l�6�f��Stla�+k,��\��G��i�mp�jc/(�ɡҹwR
N:h���5N4{��� w�� �zv�~��15G7��cL-6�	nq�TM�*�Ȣ=���ٺ޹r�q��3�~�eWI��>��BwwL�l��o����u�����M2�o"$Ql&�q\p�g-�F�[|�R�!B߈�=��4H�+��%d��#��,��w6��:��B2w�)��:�ÿ�o��rg���!�z/�EEd����yj�:_�4����p�Da\X��CHU�¶�v������_P?���-�1z���[<5k."���x�ҽ�{)d8�\�0��<Z�zn��T����v_D��*L�9WN�<ՄS�N `a�/`�WU"4ǯ�!b_-��`m��wj��?lj���뷻���n\�\꺸5K<�8ď�y�2�9΁BV�٪:��������ǭɗ�"0�C�	���+[2�?�r�W hh)ᤆ���a
�O\�!݋�.k����� �d�g�"�a�:a�b���?����M%]���e*����ҍ���H�����$�B��@��1-��T(|��2�W�<���k�_ƗIh'�lPg�T�p����l{��(�"&���JB��y;P�pɼ$L�z��
�IEFЬ�>�tA�����R/>V�<�(#p����Hӽ3*LA��_r�&b�8?�:3z��L1�T]�0@�(���u�a꒲3���H���!�{��Pa�Ω?��_���4-@�_v��Z�S0%�)�����Y�w������S7�f�7q7'"��e�4�̗R��ѻ ����19^.��|�#�?��>�����rIW��	�:BZI}�Q�&~��)�X(�:n ����*n�tЏ��t�(V	��R�Q�t���F�M�è-��s[XU~aU��G�
_���DR$�,��v���#`�%|�7�)���x~l5��p����x��=��yf�
 �Y�j0?�4�wJ <�X���v����df�C�sHa~$CL穟��`K�Kǋ:,�َ/)��'����8���S���kI�9�˟�����sY�Xҷ6$l�~I�2Uh㲈wWť.�)�oFOa3E��Hl�`����w�/��O����f�7�z2En2��.<Ӹ�]^�l��[�1�x� �qb�Lm����Ѿ�^J}��?��#�����ڒ�9
��g˂V��Sͦ�n����d�@��Fo8���::�,˳���K��˳x�w�b�cy�,��b^��4q��r���j�&$<���Y���<������+b�"q��o��뉸: �
g��ڷ���w��ޅ�����V@�v����UYI�ͦtZ?X6����-d�i7��589�c^���~���c��z�8����G7���fT�k�J��%�#�s�i�DG����@~?c�R�'��O��!��s�9@���OXrn��T�8T�
�.��0c��H���0��->,=B�9$�*�MX��	vՒ^#��҉^��?h��ՉEMPN�{ay��˔����m+g�whh���F�`�#�l�p}��.��7A,���)O�(͍��I(�L�e��!<�!0i�ݻф&�����&{����)�g�q�{j�������uz�4�>r��T*�Uy:�Q����2ٕ3Gq�}rP�5� �A��Io�C�خ�C��S/$J���8A����:�//Ek�S�_����VE�GE#�C�xAm����笌^hcb6��[΂�C����
�@�f��0g����ښ���Q �)Ҁ���굜�p��8�Ft+ �T�N��f;�h��,�qHI~J K�#���G�΀+d�>ΥO��B���Q1!;�Ny���SM��*��ҏ<��j^��(�����~A�Q!����,H(����G_�9+/a�q}��a�
	�������qƚ��KeJ�Ƕ���.gJ�a��˕h~C��Ѝ{���>�6��tvwh�E���y.;�P%�is̷
2<��v����u~L�|�#PF���Y�C��Ȁ�_��F)�p��"e�u������?˦umn����N�+8��],���'�WZ���e�y�]V%>�2�m��J�?�u� �f�.���#� ��A�NV�wA]�܍I������%���a�<6ˊ��  T?գt�
}��U��0@�|�le8�m#l~��X$�r���ݐu<B����>�ѹ�m�=_�1s���*�Y�x�ܷc�PG���4bFY�a��LϢ_������{� ������G�_�)e4���_}}�{�A�sf�Z�����Ꮼe���t#rl/|U��S�< ��g,Xc���˚$�PK��EY�������HR�I��Y�*Fw�A�"對�߻�Q�zϒuT{��GEV];.�}�pj�jd%ܜ�!���<�q�׃+�o����4�6��޸�]c96i�L�b�8fu�o�_�g�@�����},���_��m�+��њ�V�b�"�8��r~6�����6����t�"���iLYWdH-�^+<���A�'p[�dG_J��m�:��y�v�oxŲ�=�Ebr��0��n\���IC3�W��=Y6{�挽�C��0֎la�(m:�Q;�Υ��K��dOï0!192��ɼ/M�F��~�0�pD�+6�1�"*�
H/Hn��J�n�)xv��I�D���)�V�8�ґ���x�?�(�i+/�co�!KdrD|�9���r� byj�Rl������͕�u`��&\H�#-j�F�+��%Į��9�,�����n��蛡k�¬a҇h�e;!1z&` ��>�p���쁶om-$U�~gͧ(�ؤ'����Mg���
�!^��KJ�w����l�m҇�kV�v6AOHU�,@��>&j�9R�b�����K�����N���[��;�
b��,�y`��phZi�L�|E- Tg�<�ԧ2K�t��]�.K$�w�^W`Vx�Y�٘��!�XLrAf���E@��`�-;�zi��m�Ǐp.��-&�!8!'�̄1�;�H8��[n�%Q�r^��t�1p]�����?��m֛�?S�m���b��p�S>r�]��1�z��Nb0�tI�D�I=
A��.�s^⎭��j_@O&
?=�﷘Њ.�g�SzX�C�e��n��EN ����h��?���19����t)f'v�A��s�bI��6	:16VI����s�ma�*����]{��Kk�[�X6��3��GďҮU�O%��O�
,R{VŴ��AC���S�U^����_�"�=�7/�N�価a6��e���,?���+��`	F�]�V�
��I�����}z�(�X�E����>�Z���}pM����9L(D��e?Y?=��ehEy�h�:7� M�1[�{�VEa�=�ib9���~v�3%�Q}���	��v�I��g>%�v�'�+�c��b�[�3�&���:b��)�����I�4�*©�R�K����}�(�8^��;�<"��G��f�>S@��/�����Ciy}��3���=�N����ݰcq��~�C
Pke'�!?8��\�)�rDb����Fɴ�N��
Zز\��>��9b���+�_1NNvn�b�ͱ-���ó�B��4���@\L��\��/�&=�N�8��"�k%f$���J������Ϋ��\M++�ԐS�*0�Q����E�wX8'�?���L|[��c:F�!���YZ�����j��m���5͸Dgmtp7*_�_�����Z�h�����-�9=�FY{�G��7t叴�SW�M�]�]"�L^X��hS���`��(O��$�[ʘy�0�W1�%�}٧���`��I����dLk[�_����;�q�q��:M'-���Z�%p��c�rSy.a�Ѓ�Vv�,�6�3B�{A�Ȓ�ecC�<TI��!��j5^N�
��������	p�t;p�V�&��	:�dʽ�z��O�$?��X-A	"�*i�����aC!=q�����=*G_��Ѽ& ���MoOWnWtaxAO�#m��u��Iu�޵���zÅ��۳�x`?�P����.%BTƓ�A��84���v��=�K���	Ѓ����R�yA<�e�[sը<����8��̵��_>���`��ڇ]���W�߿�	c"b>l]Y�|���j�yg��l���U�p`ۿ�&��Q�n�"a��Ҡ�Hզ�&�#��nQ��aZ�_~�����-�K�M��f�h�|w��k,����h�}��f��d�Nѽe�6�d��q
B��V�Z�^�OG���_(M��9a��R���::����]7j iO�څ�"q��Eh�3:��	r�zhFC8'�!ekd|=H�Qwj�0�f�K�臤���;y�NJe��U�b�[�vm{��w�LF1Q�<�?��y���