��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x������jTe�)�D�b���A����1v16�|,J6l��)~�S� �B�`q���(]�s�ˠ%��L@��z^ߴ�E����\>lt܀��|��>Y-��=��v�r@@����Q��2��^ԭ>=h��^$��f]vY� $za��"O� X��R��ȿ�u��v��\@��
��^(9������U�M4�~�&om^���O�|�;��9J0����E�{pY��W��AHgI��o(�s�����SL<�9K�	���-R��_�l�gI��9M>�5��׎m�C����E��V�e�C�FU���n%{��
]�^
;{*�>Ԣ.Q����ǿ��z 0�/��	c�� �(Τ*�?.Sڦ${#f	&��I9�z�u�4[cݻ�xV��PI���yu��o�����s�
�nVX6�n��-֐��&�:n��'`o�҄p�����"��/=V�ⷝ"���;�~$�9i�>�"������"��I��q�1��]k��������&�+��|��4�`���S��s���R���7�sYOC?i�Ï ����ʻP!��ߋE�k����Ԝ?��A���]�s�E
Ͽ-�Q��\t�0��H&�ȱ=��Ҭ��,y�#����Th���H�ZA�X�֗EY�}+��x!�4;����{tR��g�wD��;�&{xc�����&�p ��Gj�e�G�j��p�98(O@F�vϚw\&��ỶfŲ����q6#]�R�����?��.F�3m������*m�!D�S:��1w�NO�q9���h����aK�,<"������/x�:��V��n���g�:�k�>�ʺ�6:��H�u57����W���r�U�'>ރ�=�<��V64�Gs1^䝣,�ў��X�0�Qi	�a۠�-� ���xߢ�y�[��0>��{�1Y��'2u3w��i1S>�X&�m����);E���:`C�W�>$�BF�-���6�L�g�8�,�7(�,�(����0E������21�Up$p�Ȥ1��x@
��j5���ǪV=j�5r�j.�G��IФ;�/��BJN*��O<nPJ,���}��{܀5���qi
�0�_���>�JZ��5W��� �����!� �nb����:Ōk���O��<u:���C� ������Y�
*u��	ݶ{��$�E~��}�o_�$�I�o�̔H�=��Z<��v����� �Υ��7J����3��Y��3�Z�o�C�s
������{�'Vǒ�/�t�h�	�5N�Ĥ»dt�$݅�ʏ�JG�'!��� &��2��H��촿�O����Ŋ�����|���?w'�_�H�M4.��R!r�vr�]\j;��F΍J�ro�%k�4=pM4׷m���8���N��C� �l㘲��3r]�jSh���ʺ�8�ϙK�Tu��x@]�
��d��*���pT��X�R�&I,~x�k��*���>#�s|CR�@�fc�J�P�l�� b��U��kE=�H�0N���(�'���4Ɲ�FxN�h�.Q�"��m�y��T�=6��C�Q'���z/�6xuޝ��������Ku�6�u��Şwg�A�Tv���������5JI��:՞[���	�| w�xm��I#;�����VUi�S���
����[fB�#0o��O!!�y��龎Qt{Y�Q�����F�K�Pt���瀾Y�Dj)�yn��>����'��S�Lc8͝�_7�g�Ēk6��)�务t�<���ɢ��L�����@Q�������P/���t3����2��"��F��Up~R*��s���Z�e��>2u@��N��o�*���Tg��r�m��@��Sn��Ɓ(�㑁$8�'�M�V�*\z��Ww�e�y$��#k��x��g�A{D� ��+���E�s3H֬��\�4�i��7�J'�TEd�b�vN�0$�|��F+��&� �N��%�٧���Mc�ȐQD^17��(]��y�$�i�>����pF�*oKW����-��30���}�<��)�T�みL�
U�.�lЌ�~Q��v��]��$�[�d�i#�Q�/V��%����M�� ��ܻ��9 k�=p�*G���J�뷊8��i�������j�cۅ��ّ y4qPFt;�<M�M��4�̈Y��㴃����֢�(��=�3��s�Gd",�d��=�v�aDH��T��o�H�g�������mC���pz-#Jemd��)ݴ�sVA�\�M����c&z��z�Y�����F:}��6�u�A�J�MEu$>_��i�\�p�w�����������_�"@ղF[X5D�PJw
��ԙ��z�%��a�$����$����\���nu��a��� �G�{�>ճ���8{�l�bscC����Dg��<$�J�UJJ�w����)^2�+a�鰩�X�ux!v���������	n�L=���|�p]Q(������9po�ЫJ����`�6��Z���M;��Dt�}���' �(��)G��l��G�f �m�*м�*�꿗�=�W��k��3���e�^h�p��7�?��S�d�,�r��b���vR2)j.@;R���1�E�d ȝ��m� x����m�D'F�yV@���K�3��Q��ig1��(A`,.L��3�bo�8Q ���I�΢��JmV�>�0�T�Z�1�o@E��Oi��AK�3<��o�O+7ߘg0�<�	 V���yE9ڪ�n)� �����[T�����Z�F��<��=�QH�\Bm�η���B<���z�;��_���҇Z�:�LU�������G�P�L6����':����*�c�c�������@�pْ֤�ێ�JȚ�y�kTE!L���˷kh�A�3/L&�@}V�����U�ʴ�f�K|������u�a{�u��T90��v���y��Gn���?9�B���US*���f���H��-�}��Z��w��顜'7����5��W�N�)aҋ/�}�1�2�K5p�$���6$0�`�a��V���#7OZ0�e�HW&x���Gy<iQ�m��\�3�/��t0t�!��KR�Pg��"�|���.:$��h��u��f��xj�Y��q0��4x%:��b�k6�/e�0�k�����>�MR2*^-`�m� LjH�/�,�P`�S�*��e�
�C�˩�[^��I"H�ee-N��Y�������~h�g�=� 8�C�3��?R��ref��ݠ ,L�>c"E����%a`΄�~��ygl�{(�{4�7�+|(L r��8!��Ì�$o���8D���^O�_�P��̆O��A��p�=�!M��?���	_q��eqD}��?�������S?�0���jid�X�;�҆�<��)�ن�Z�e�i��?�$a2 �Gw~]N�r���i�h��Vpf�����:R����F����A�Q8[�K�n\��h����/�v�
En�{��y5���&���'�9���gg�C���2�XR�B�fQ�S�xA��C��Z�4
=ͻ�VU瞃�M�3������у]�)>4��B�<jlW�$3�0��݇��: jLsN�ލQ'���k��d�'b&�F@�t��h��R���E�%I�9�bF��L���l�vs�=�mK��qʀE�Ջk�!�n�n����`zqe�uF�SR�<���\�}{��xG%}q�*�~׫D�܊(��o�jA+�+{EskOEy3;^�r��Y����Rn�
�-,I�i�U�Nx^��&C�g�" �ˆ����;ʷi@4�mUm�Q?�G�k=��t���lA�|}5����m�%�Hw�������p���r��?Nk����.��R�D�|4k�Р�����y�}��H3v/Z�%����E�\D�迦/�_|�bw���&��b���xF6�U����cL̍��״�b�p�;��������� ��Dp��l�wP��P��3?�Q��g���6�&d�F�y���(����J�s�7��y*��j��>�c�{��LF�q�C�,�s� s�����������R��y�p��t�rf����Y���B���U[i����]����v�`�h-a�$�o�@��:�)V�����<��=���/��U��x,�d�V6�������	5ܙ�l�����ۦ��N�۟����)b�|s�u��������|��H��h�A�zS��|�{�_��5���[Ҟo����S��X�0�)�O��\}
ܨ�f�8-xd�8s��E�Ё,���4���!��ۼ^����إ?��H8�/B��b� 3^���p�D^��c�+Ǣ����,�	IoM���v�G\��{wnu �t��6�7;� Z�GEr��]����0D�)w��J�����3ڶ��A|�ϴ�f3���rB��^�/�P����)S˨r&���]� �-�Y� �{b�r����%VI�ʠL`$������Cx�w�?��Y� y1u?K�5���Q��#��'Sv�P�~�B�=�r���Ҕ6c`���R|<���0��4[��1O�w^����@ه�c>�}��/��r.�})ɹ��x��c�2�y�L}F�t\3���(���ə�GX���ѧ�-��8w֮`�$b~�[�6�.�GU���;n�Unmn*:+Q�T�|aG{��}�p�K��و�daU�Ei�֮��ԡ�ơ+�~��%q;�(���b(����y�/�%]|�[}P_G��*R�A���0���>�ڕ5gz��C 0���h�}P)��C�7M�g����η��(>{�ZX�����0I�T�@���C��xj�q��נp�k����!���3_�J)��vLzh ����/�����쀻z���\/�ǒ����z�Fj�����˰0b��U�QL��ԥ&����+���_1��"���c�;䵨�w3��� 8�6D�����ˌѝz5q���[�
��5;޺�\�7V�(ꥆ�F�ڋ��h��d��&<�:��|AL>��_�*���О�X�����m2�,�4ɖ�m�����d��J�}�	1�w�A���h_֒�t�C(+��fv�
�����V�l�Rj"��:�\�����u:NV��{�z�z�tW��-�>
&l�0��Σ��hCHAAtA�~�����鰐�'��,Q� �ˀ��bV3=�1�>��8b{Vv���
�8�$��1u8@���jUw�7��B*+W�@tה&���"������/���4Usg�e��%g;�������jų�(9�-Q�OLr����b��d9X�j1����Ԕ/ٱ�,��'�&����s���k���}��߱���Y.�-r~w�V��0�5c':��'�rv�`�.�����/�����ga U
2��e-k@,sIt��Y�٫�2y�w\m9\f���a��|۱]��0>��@1s�@s��e���FT�[��NO-��,ֻœn^@�=FWuLɗ%�oNW=:>�9W��IpU����k4ߐ��	��t�.�j!L��}Ǝ�� ���CͰ�����cZ��`�G�U��!w��L8��2P@�e>��o��}I����z:�������o���Ө~���Q�+)�*��9S#�����;yy��K����k�I�A�N����p���1~ƝX6)ڹQ��7"�k��)�C���I��Mӱ̷�� ",��Zz�1����L[@9�A�-�B�k�+왖�$lG��Ci��|섓!9wv�D
���T��wi�k:|d����|�]P(H�-���P�c�~o5���M'C�F�#]=���jS�\���̹�_$j���>B���X�ovߩ�J0��i�Gcq�p\�Ǧ@�߰:�&^��J�$M��G�|����F*����i���h�G����7�He.d��~�߬%�y��`�s��_l5��z�h�x�N���Q]F��!��n���ۀ^I1h(aH��8J��
K�Ƙ�>lg� =�I~=��oW�x�`���:D�&'�iV�R�F�"��
�z�gn"�4���`��S�VF�o�{�mEli;�Gmm����#x�ܮ-��"�H���*�7�?�"� ǺVH�_)�z�b+�cH��)���ʦ�����L�4~'
��qa[΂�/q�Ul���*e�ǀ��6yRq]�i��	�����ؔ�.R	�"��E�����8�w 15�����&F=(`}����5e���y}GZ��s�F�;�z��E?Q�b����&公��|����0�94�H+@Lݍ�W4��M:^�؂�-����g��;�b8��~& ����|Q���3n��t�+��շ���c���锨��{<�n�Uf�����R��с�R��9C`#���]�[���q�L���H�)j��3���>�%��޾��<DK̯h�mp�f˖�
z���#�1Nj���U�-S^��x����)��l�މ�<��Wt!�����y����y���u>�����h���{���9OcX���#���|�Bj�!�	�w ��j@�*>�Y��cA�4*��3�n�~s7�㭏���+��s���{��a!���p�{�+���H�T�?1?mJ�� R`�G�/岼	�G�n��0���'Ct���P"��1�)7��vUǲڀ�@B��b�W��������YT��Uz�C�
F>�S¿%��R�:^���� J�����'�
���Ob[�r�����:�X�*���L{��Z��ڜ[��Gj�$�a��酩d��*���}[h�շ��������~P���aА_M�,�\&Ip��f�eT>�"3J��y<�=�H�(��(��<z�����;H+2��%k��a-/!�F��s�;�;Q)G��F�,A�{gtQ>��{���Z��a�A{VE���R���TA�<2�4ٖ�����4Z���%`#�9Ū?�6S�+�����4{^9`1AW�o��x�92ry��)�뻱�ֺ�ݸ�S��¢�m'�
��ʢhP�F0��?M�E��(�JK,����;P����e�w��R[P����LU�c���������`����z�D�0e�O䤭�2�)�5bz�F�2��`d&�G�|d\�}A8��ώ�M�''��Bp}�Q�<�1^�#*u�x�-���˪��mQ�|yc��M
�3�:��ؖ(e8 �鏧ej���?�n�NΟ�,&R�9K�@ݰTE'=ܒ�?po[jp�病K�k�h4��b?�-�� b~&X1/���}(	P�dN���'��|�1�'CP!A��jz�։H�Ž�o�������������T����
M#���K_4�V��B�s�����F�٦�z�ƃ��ks���VJ��C=�� �ެ���GW�����W	�X:�bW%CB>Ȯ�����'���y�u���AM��,�&<6�W��b��X���㎏�,���UN��[���l�,u�I2�t��en�ё�n
�J���2�9	��s;�ʫ[:�g"2��Y��$���7�G%���?ՌLC?5m]���0���-Ɇh�@���gQe�ӫi�^@|�|㸠�ި�{qNa�Y�PW0�<	EjK��:Iw��@�]w��jC\�N��O���\�A��c�����:�9z��Ӷs5�<�P��~.�w�^r�g*�	���s���F����^�b��as�v�ÎwC�yNهzs�]�"��M�~�DD_���7�,�n(��_�<[a<�@u����'e{5�[�����S!�a3�����0_�u�=z뗅�i����:M��HNi����D,�̉��kN��_�C��#;���I�t��"��g(٬�����<jm\&�Onj݊3�x��e+���U��V��ϤmgtgUT1�}��Q"1P��ad�*2��%�R=�~�@��^��z�������X�i�l��װE�~���FB{��d�P
��W[�~eG\@�+�������^j���n�g����h8ΩskV#�49D�5ǆ�I�1b�H��,�}�8���!�i�K�� �(U�Hw3��j?NO1��6x�N�Q%�Zj��ӗC�7&�<��I�r��<^M�Ñ��?���qY��vg��&�lӝ�D?e����P����G�^�::��y��7��c�$-Ɇ2�X�6�ܪHƔne,���K�%����	o����/��Ut6[�T�5v�ɗp��
y�`�<.ѿ��3%��������n�\Z����N`���|��fG��חa��'`N�SG�C���_�'%�}o|��u�Jd��*�=�O���i�����i���r�D�(.f��нn��xx�l�$�~�����)x3�5���";��ӾK��Ͽ �����	N����N���/B�;�])vb� �٤1�V2������@l����7���se�����"���_����G8Hw��.�N�TBrF&ӖS��o��X!ś\��q?��3N�}�C�&=�>�f�Aq���ۄ����h�g���)�Y�d7!�����<g>�%/�N��Ǣ{��F�yڄ�k����+��Ip�C*&
5t�T{`�fT�&΋��iD�[�Msb9T;�S%�vKN��h���f~�=ă�~�繱V��Uc�á������
��}|Mg\I����.ō��9�9*<ˠ dx�!�,��m���p���f��G
��#���87
q�\�ȿP��y$yw�̝`�IZ�X�Y�oG��/&B�.����r%�����o&��� �d�#�)�В�7�J�9��x���њh�m*ϋ�t�G\J�zO*&�C�_/�7�giO��9��/�Au��._��4R�+[��������tI�V6�E/QQ!����D�%�ĩ�v?j?�[`�s�h��ޥ��*�|W��b����k���|$��Gf��?f�gR�b�v��#,�L郉]�%��N��N۽x�"�8)G8D.|x�^�?e拖��8iJ9ڳ���ƍ-�G.v�s�7���x/�H�ėM\7H�O|��¡���_�b���M��7W�ɔ
����,Xw� BU@��a+�b�8<8@r
 1_��i�UO���zcҹiG�_��P$a*-�zޙg*��Z�x��]Ɉv�Q���y#_�/�<\ID:c�5�����\>ޮn���bI��4�}ŋ�K�B�zK��]LW?�I6|�-=hj�y�t��+HYRp���nBj9d!(ނP�mՃ"JO_:p�j.A�f�Ff�@ z��Ͼ��,~�![�dJ�AOj�#oj}�S�V+�����z��DW�V�0u�!e��@b"U7��o�vgc���Zp�֪g9?�}w60���=����ut��!��j.*k�7�C��TN+�Z��3��`W���W���ܳҀ0lðv�fpP�����"���Iy�\ʥa�;��O�k�_YD� j}y�]��|�2���k���`H5�h���F��[�BŤG��E�H�6{�^�D����>d��� ���Ch�&�{�ߊ/�`U>.̬����º��H5j(�/֠��l>����
���&�o��,8JF�i�a��%��g\�BV:>[e e%�n�2�H�$�����7V���y����W}�r(j#I�TT�%q�z��iy�o�Ԟ����4�?װ�5��:��U�ٱ����ݣ�nc���GK~o���M4�y����0���L���� �v&�!�;)��̍'y�Pw��J>�����%*[.��N���g�� Ò��h������Ifn8�F}��N���N���j��i�n�A��@��A�o*�H�x|�L�Y���t�K�?�q:j�4�;�ٗ����A	��;���7 C���c:+/Owij�>�������!���j�O�/c[]C����e@�8}̶���[��eǍ��?��(6��*9��ͥ�:�NYpyqU������oO���������Ⱦ\�qG��0� Ș�G�0�*����y�ƻ��gx����FK��1Rf.���ص� ��kcN3����z�ڈf�O	�/�-�upH�*+"9�g�>K���5�\BY�=Zt��W
�w�˻W���q�R;��!͂�C��3/V�F�;�T�K)}����V�5n�.�΍X��䔍��ĝz�<���B�FU�%	,t��_�y�UUw�mze��ƄS��ʹ\M௢�?aΐ����$���f�xAa��E��������Q�o�;�h�,9(7�U�����1��GA�dhh��ͺ�%�U���ha���:&��m��#���
�y�:25N�Hޝa�����E[���z0$��?z��6?T+;���ۆ
�/7��Q{Y����g��\lV�:��'��j���vx��HF�aZl���;�4#�eܚ0d�f(��5��v��6/e�4��~+�s?�[�$y���>D@��Ҡt�r�Xʮ 3��L\���Y�.�O-Ρ�S����D�y{����It#�i��~cpu��=I�+`n`���،G�=��7�g
��w��wn�f��q��T���\����A-���ի����r���ώ�j9���m*���o�8���4����ds��;�?�e�]���z3"���x*а���g�xt�hO��)�[bWųT�k��4K��2�-���Y�@�؜��Qܮ�h�,��^���xX���-�2��̶�Ɔ�C��<p�l�3�R(U�/��90��Z��(!�2�o�%�Ϩ~s<�V�Qp���L��b�2t6�O`��T����H	-!�H�Tx������`g�cтT��~(@g�yHU��Wݤ����0��f��~�ɪ�j���p���#���uJQVk9v���C-'5�Ǻqh��E����[3�������]D������H��ؒ��~�[w~��_C���V
w8hm�wJ[����BW�b����K�UG��S�� ����^�^���`jC��3����ߙ��2��B�;��w�+���q֗�jG��_���j"�;(Ҥ����o/�l�?j�!(�#e�5#0f%��?N6�����7>]��$��ǵ�-�`����hU��\:%ZQj�bM�n3)+X�v�l����Y���m����9Z�p/�_�����.������[�LW�m�~l^�N��ehs��Z*��c�6e�3�Q
0C����Q�o?�l!��{w�}���2�n����]5��z�3h�s��j��)�;���m�)�dS�[_/� H������3���l�3u���x�
K�\K7�GL�;��Lgp��*C��Gl����H$�h�����0yGVDpq �! g��>W����ҟ��r�r�� ��}f��{E�kO�1pw���[�差��*�ʐH��%Z����P������#6�-p0*>b�E���ͪ4��-�ܺ�!*�D�/@	�iJ)e*2G��[�g��*&���&�p�Z;�O�m�������/�s�q����Q)��� 7�Bw�x���O���a�.ֆyS��ύ������tޜz^�Y�õ~���Bc����3��q,ߌL�vg=�.�+��M�;ɖ�-�ix6��RF�q4�s������QO@i���̓ե�.�)D*w�eH���'�}ɽO�v�1�A��EE�c��v�6uɣ@��#���bĜ�a���?�0-@[��N�噐�E��{���a�b+�&�I�3BRZu��d�HHA=.�%J_���2Z�nآۃ�c���t�:�����zĶK��4�K6ϡخA�Td����l�@��A7�Ϊ�m}f���e8ͻ�j>-m]uS|h�L2=U'�^�=���0y)�?��k��r3�[��"f��>ĖW� F�B���,�w���?��g�3�N���U��:�ډVPuEhM�Od�^�h�d=�3F��$���tǙA-�Yo�k�nL���iam�c�T��)ی���'�w`\�j��i�9�#���[T
��>�xW��?�,DC��Y�d�@�z�G�3���qjKX�#��;5<�Y�8�ivl�gͯrP{RHa�*u^��@�Un�n0���v�Ҕю��Ssm��Km,	�8�`�����B�b��S��i�RK�$��"�r�9����]Xx�� �y  mP`}N*/�B��������ւ���Q�P�����S����ȧh>�7,�a�d�^7j"9)t��w�թ�އݔ?c�DoM�[P��e�/�gM�!?%w}�-iW1�iAZM��3���[~I��'�G���g��J�<��9��������Ǭ�ʉ-Y���X��D�ƅ�"�9��n�Yʪ'PX`�uׂ�?s� �)�K���Tpn5�;l���)��czbt nU^B5,|}��aڗ��\�
�
�w�3��%*a��a,9A{r��nj�0�w�L���w�3����D��2�lR����b�~♡��'~�k��f_$~p;ʿ�������q�	@ڠ;:�m����#e���G�j$����`Be�I\$�x���������,��P%���ǿ��ߥ�|,NߵLũ�m(s=zC�I0�Z� 1X�s*�C�����V�R_�$F�����:�� ���DmS.v�4I�8�?�	fh>xO$�%�\���N/sTyː��'�vG@{q/���
��1�đ�߀+�U���8�rh,i��Ky���B��wlTΰ�:5�>�� �ts��7� �`�׹��o�w`�@="�� $Op�O�Ɓ�7v(0�\q�©F�iɛSޙ�-�9E�C0�x꣦Z��`���j�5����X,�\��֛[���	6Sw2�����Tv"�́U���DI�����Z����ۈ׳W7\h>$�V��3YKh����a��GzK	�n��f`)@;�6����8_Qe!�】3�G�N0�ϴ͊�s��w��/[/#�}7(���_�{�).n糘zQYq�Y��@,/�E�'/O4.��sBu=�J�������׽���G��Z�[*���s��c�a������7pUv�j��%���/�p*�V�8+��Oe3O�	x��,9.���U�}�cӳ 3�u�Y�2�?Z0P��R[��G����.D�����}����"Gw��g�_I@bi�9KkF�>,�脌���0п�GPed�����wt�Օ��9�VD�f������'�t���%I��O�L%��rǵI�����/����|$Jɯh�9�K�ms���L�.���h,T�2@���9?�5z�W��S��u�צ����.1��|��QѴ�|�]ط��4�W�P� q��u&�`�w�}'ny�� ��1Ҵ�ʩ�]Ek:7�5���fU���dʜ�_�/�e���Q�7��@�kW�`Ca��?*5��J��������
sN��d5AC�y�����b�Ih�ٷ���*�+ST���9��
��	h�mZ���n$�Դ�a�ɕ<��o����N	WP�K{	�{�^�,m��O�W�i�(a�ˆӹ^CH}���MQ-*�Uny:~��� ��1
���Y{�rA�(��_(쵇<@�=[��N^ý�:0������L�]�VZ.���5� >Y�n ������]{&�=��z3�a.ɾ冭^��c|���%=$���M�6����%0��@�<)��QJ���R�4���s�F�W��%������+&"�.���6���e^���0Y�B���4�K����<�$4\���c`X�0N�U�<8��#ԟ\����!�rغ��o T�E������hR�w�/���v�uv%�P�0vcW�SdǙ4�~RQ��h��.^<<Ȑ��qZ�] �<���b�����$0�8f=��f�;l���P��;�7��� ���!	���O^�����1û�u5��d�:�}���ԫ*��IOh̫��J��q��ٽJT<	O]�%�
��5?Ǽ\f�*�M��l��=���C&�)ˀ%�,0-&�2�I��t�d8'
���]��K�.�SP�z�P#������w�I��n���7����ի2Q/
(@w�D�h*S��Cv(8,���R�>Pe��˔�!�����O$�čad�hL�-�?@/j�3"F���,e��:�D'C�t=����m�/V�1`�0d�|�#��_�u��i�z@�N�Gx��B��0G*��D��I $���k��lt���p<>�G�m�c��/<��8K�TG�� �U�/�j�h�W��^f��k ?^l����l®�zB��6/|�K鷋��->��G���S�7�J�J�$jma,L�C%�.��h�e��NeV�(ȸx�	��zd�&�5��,�� ��>}ފ^�ޜS�jG�pN+X�hI����}�?�K�䭊� ����;A�z��¦�Ǝa�A�O�>�o�(��ٟ����׶O�tA�N��â/ڰp��䱴7���r�E�*�P>J�5>��k��i��6��N�>��@ϰR|�gB��ġ��})'���S������f~�h��"�4Vx������@�:>�]Ϟ5�����!�!d9�z�������| �8�������rt2����]�q��5����(�J�p-Z�c�a��>�0�Vs�x=����������T���� 0��(�b�Ɩ�m�s�{��������s�V*"�c��幊Yz��<�
�ν���0�ݾ:Mo|�8��泫*�Zf�+P��xhW`�;�]��`@�	���x8�H�3��\N/� ��8L�h��K�0.K���A���j9��G4��3�A�,M!�G���PDK��j l@C�'k��{��T[z�I.��|F;�ʘq�*��q�zb���L-�9�zY([w6�U�')D̊�}p�����E$v�iOX��d���S��!8|����>���c��]�Cm���v�݋��ģ>��<{���Q2�P���Y�@�ib	-e��\��V��0���+�Йx��9�����N�?ݗ��.gozsъĨ,9Y�'���L�ᓰ[4kZW����9�FU\^ �Ŏ�&2�����bkGPD�u��k���@�F�BM�����S�r��l��]����tnG��m�ےө��R
b�f�R:~΄�zRǘ���K�$�9�"�mIT�p^�.,���d�/�H7k��@�NFW������\��.z�?�Ѱ��h��nt�"b�\�A�Di�K�Z� i��:�ս�(��OH�=��p�hh$�wp��<n�t�Z��4"�kJ�~��)Pp��@G�/���&���}�̚X�����l�`~�TuHp.�Bj3�y(y��ΐ�_�� �3f���Jˆּ��^̣O�b.乪��UǶu��b	���M$�;����Ry&^t��A�y3�_A'�'��O_A��k���B�c3�0�]PV�"��)��3B��M'4T�A�����-�¼��x�ؐ�}:� <׃TUzX;4]x����+�>CYSt���	-/��ٜ' (��qss�]4�"��\���CBdK��G�6qY�,�Ǣ)�HF�5[ꑱ�۵^�-��L�8qt2k�bG�E�9	a1b�
�߀9AEޅ�|��|"�]�v��#^~bE��R���3mR!ʫ����b���Z�9�6�^~Q��C!�8�����5���vD�VYiCZ�'���s�#���d�M��J�2�d�D�{�֎v�/�p�9|/Ù�c ?��wV)d��	@���#�T�~��ҁI��Q�sZ�"����"�u�Sm1���Qt
5}��T�gU&�r%W����@��0g���p�� �:�.k�y^�$O.���
��H]	'0l��Xp�}F�R�1�c�v3wu�÷���^�A�����03�w�DZqI�l$n}BP7d�pE���m��X�%"�]�.�,�	��uUJ��p��K$��d�g��l���{�T��XJFE���<2��\�K�*r.�����4�$J{�[n����~�Hj�A6�	2&]"� "���a��	�m�"����_�V��4�E����%%�$r�c�H�ƜB*ƗCi���/hi1N��X�E?"L��ҽV%F	���_.8�/#ގ$����>:ğ�?k�]��)4�CzP�G����uX�5d��+9��A��Ӯe�ɸ0��g�~�戦�e,��0t����g9~����W���v�ye�!-q��e�'Ut��{gnZz[����eQTj90#��g�s^��t��pBy�po�8
�Ù,��G�h,�� �+d\5�����(�y2��0T�������'ُ�5){�#���x������5�(���Ǚ�U>Hr3��/H|S��#?2�����96���!pmv�.t.�KTوs�F�/����Ղ!1wGiN�o��� �lR�ϯG�	[՟$�����>�fk�=T��������
�'(؈-�\O'�O]]��׫ ���Y�&�aԖnyeWPg��tQ"�v`��MHK�f�Z��� a	m�5�Vr$��~�ŝ3����L����߷ap�����a��Y.�#�y���[͌X�i-U�s��`Ξϭ������W��xwi�}'��=�Z3�nc�,b�Hr��C8������Jm�P���u�!�e8�s��<x��@���%�pR�����@n(^&�8�� �H)!)b�Ԏ����A.�ħ�h�"L�
-1��8�B�v��mE--����Jj_��Bn>�v�<�W�d�+�އ�x���҉���D�l7�����V��If&�`��,�e`�:���3����f���A�{�	�71�uE�d�C�3%��5�Pp`���8i5�c������0�F���w�-Z�����H�� )��&�M��H�mTz��mJ/ʤ��$�v
C����y�w� 
7H�^IM.�Q��O�Jr*���F X��׽v������ی:��JY{:�F��^|��hxi͹���j�r`�k���a�U��ѥ�`.����D��'� ��I�z[�G��EV�	}�@�>�u�� 򟮹��^#��5Y�m��N9�sjg����
�5Y��]2���et'盪*�h�]�N�6r0�P�c7q��o.="���͛��=��j�EL�nj�M9�)ueAsw������XE 	����C�3�w����v�����WU���Ơd-�ڤc	�Mvw�X�}�|u]� ;����{����Q�3�^[b^m��̀T.���2u�2�A]HC��y�Q7�}��j:V�)����C����w�)��iD����љ�36{zB��g����3�?,���x�����P�|���+ �Ҫ:W���e�VQv&LWq�M�7�Y{�BR�pL���X���!�zy�ͥ�F�3���/�ۥ�v���Wۄ�G�&@t�q����kg�`��T-d2;�5wʄ�	�y�_nQ �ljG�C%���(l�=g�c���6��Y�- U��q59�����/>�h�����G�?�XfI/{�2o��{��W�X�T� y]W>h'$��Zd*IK�V�����_�2��?�J���Y�G�4>v�1=��n5�;�kZ���18�~�����=��)���}�@��Q����@�t�T�=W��@���ĭ�>�^�6hv�NFo�2t�w�p������8��+ =��1��`6X���J�e�2�z��s��rd�
ȵ��J/��-(!�AA
�*h��6!�Ip��C#��`�ǍLa��E.zn���A82�/C)�,p��,}'#�i\
<y��n��ߒ�B��'��`Aq��,�J�Çʦ�{Q2R0��~��?�B��ǁ�vzMX9m��´����d0SӜ��p�)�R#��9���@A�g�A����A����k���{�L�F)���r�Lm:�D�+���i�
�&���K0 ��>� �]y��������tKye)A�s%�#�b,(��J��ثⶩm'm��y�D/$[2IS���j���,I>EAG5�|��o&�
[����([wkECY�Y�.�߇�h�{-��W&�!�^#&[	9��,B�S?*>�l�z��!�6`5��g�S1�x\�1:�[���6z�<��*'�����~���{�8��,x{u�_w��͟c��z����?�5�z`���L�z���ͯ���4-h;�"=RN1��1�j�=X����A�ᨪJR,�v��#>j�C�5i0�m
�;����YO���2�p��+�&��M�l9Ӎ�2�����K���9�I���vgp"����$�r����:�S���\&k���	��!E�j��&r���?d��KL��l�]�Dٜ��	��O$cɜ}���0��'\.2��C�s��r���#����ގj���`��:�w��U�k=M7T"�䇿������v�!!�.��F%0Q��-4i�i�g~}��k|�Κ�-s�?��2s~>�L�)� .U���X5�1סl�Ez��Ԯ��� ���W�u���M�b�*�4z�w#I�ml� 9�p��*��-����9<�Q����}��p�c+����$�&��V�S���Tk���-B���뜴��h(:�ƃ�!T�^=�w�!=n��lҎ�5�2�+;������n_�58 �6.��l� AqpTY	�)�G=�nL�qs��9��ӪXF�&�SL����Č�o�[�2ٵJ �X�x���&�ܻ��b<�TBq��'���[��:�HZO����9��a���Cf��"�����3��7o�㶌'c�Z?�9#e]��9�>1�:H�e'
;�+�x�Ci�j��Y��H�=J�uM$'W١u!Z��/�����h}�HW��5a��x#/��|;��r
ک2�\�2�^�y���u/��BmFÀ��y�� (:n���� A�:"��g~�-�F�eO��_ �>H��
�v�qݙ��J�ڦU�K�F�9k^��u�IL�_=1��}���
fN.s{�u��k�SD*�T�"e�ؓ�����~�	S����,�c|&R���%�������sX?�k���湐�_.W���]��@�v4�,������}iY��߶��j'�#wH�M�aO�3	�ANe�t�(�H	��?�Ex�ߢn�8/Z|/�j	Nd��<o���֔u�YQ�7�M	iJ"g����WR�����yNj1��T��[�4W����U�MB���2K�woo�5��d=G��]I�|r�穪�Jg�,������pt���/c���a����:�t�U�b�	�\�&��=l����קD�M8K�A����* �z�]h��G����2Fո�O��2�䘹Q{�X�$�E�V�4m5�L#��X���V�0��+��22��>�tސ0�߫��^�����e�04��Q�����ȥ��������_RYV�=g��}�=��R^��z�u�#��L����`гg>pV�
!��o7	YOŕ4��qx�>������*N�l.;�ٵB��X1ٳ��!�=wp�%�l�vw���-`@w��ś|"��\9$���I}J.CnĹاߖOk �jZ���mnh&���a�埀ZlTưl`�09�G�\S�~��6�U!�/*�A���k�r��a��ֶ2�Ђ�Qh�'�m�'����s=�.B�v+?�H�>�ܡ0����&1ns��R��\� ,������ɂ��L��.vy�f�{PV��DI~a��ӎ��jv�{_�����K����t����#�h	-רPX�S��^� �d�t���_�l1�F�H��N �H�e����_1��;1���7�L�2$��`g�0$I$�{ם3Qz�v�_%LF,��C�&#�G�7�.�KEF��ld��g��Y��`�oRS9YvA��O4����P����� ���y��2�9�FN3;T0��L���bpI��3�٦ڰ��ۛ�h���ç���g�ж�o�FR��_S��c,�N�H��9�V���[�L�۬b7�ܴ�����0�%ϫ�zܠ)� ��8��a�Y����ZV~�#Oo~km��ӟ�b���u$U�G�A�?�=�*�
Q��h��0�,ߵ�$�����\�1�4�Ŗ�0�Bjr)��H�hJc�u'��'N��� }9uW�Dά���n�f`I�m���!�O6ғE%[I�~�L��oC�6J��Y�*g6dZ�Ԑ�����A Od�{��3gj9��,>�{A�d��N`u��aH��?�+����f�MA2h@eЫ��6��T���mRGR��.�v���@�΀q��n�"��WcU����f���ϛ1�J������{s2.1�s^���`�q�!�uϧ��O��+iA�?{�(�ɺt��E����v�2��i?�WmH�7̣x���_̟��$�:f|�����婢�|�c1q�����H#0��������G��MҠ�<�����H�P��%�*�r�ʟ!�cݽ_��8~�M�n{ր�:C>A�ͮx��°VK��<��n�#��D��������g�ެ��W���^��F���p��rnY�$9
�'�-����t��%iC(����еT&Y�'-�O���.����g\ݾ5��P �|{���^�m�"��YC�N�
B��Z6��ͩ��RC�ܯ�����/-�D>KH���ٹ�ȼLpM1��b�届�r^J��*H��)�U[PEh�z����Ȏ︹��.*#��@^�$M��ZUq�'���.!@ICR�� i�0b>���r{�3�gQa��t�V�W/5�-�׶�B��S�"��}Эe[X�L���<e.�GP+eoAv�"`��go	E?d��,��&)U�*�J�9Sm;�楖�lQK_����E5���jA?JX.���^|y��*��1�_7v���؉������[�oOU���?n��Ŋ�"��"W��Z��!/p0�`��f��Z;�Q�;�P!,a�w�礪�M��o�-_���0��,h9vy��K}�n���<}ֳ���1�4���@�^�`oA��a� �+��M�v�Y�:�N�����c`����T�f�U�܁�Kz)���D�e�����k�u��VҪ:�(.���P)ȳ��0�#�h��u��ܿ���ޅ�LI�-�F��g�A���蹐�)іҨG��p2��Q�&�.����rw�z��Xg���>����b�q[�:��0���������>M�@��x>�{_�����("I"Ԁ���3�s �������9v2AJ��ǐ]薕���٧�>n��]��Q���XXid��OF����ߔ'�N���{������5��K��*��CN>���)��o���j���A�C�m!^X���ƈ����ℭ���繓�.�\HgMA��Ak+)\����P��p<�q��v/`��u�P�n�pG���h����\�㣺	}�{�a�'ӛ~��t��`�FӒ�N�@Q����[�������d�v9����ÈF�R�����w��ì�2Q���
�~m��/�k�8�4iM�_�@~ʿ|>��E��J�J��d����@����AП���ǿp�u�3ӟ�*�ɀSe���0��i���D�Q�<�=������=��M`��u����-Hi���ҭ��<�����<�l�0��|I�L�MD���;�W;`8�Q�QGj1g��������j+��͓�ٸ��_w�9uY6`��i�U��;-�U#�?��m�@�.5�1���ɂ�*12#��Cx�d؝�̄x�Y�3�2�9��'��Z"��o��k͋�$A��顱	1�-�m�S|�_h�
t����i`�BǬ�1�	��~��z}rI|:��i��;��g)L�T�7��bш_�hϒ\� J\DQl��!mQ_�m-��� ��m��{]T��-lO�ۂ�G_��}\�����sG��dt�鉩Z$y����}4��4��k�U��F��8%�)�n�_q[d�N!̀��'V!ˁG��=>��\�z�ֆ�mP��L0���ջRN�ҧ�`�`h8jp�A��3��yo��ގ���4�E �i��`���b�`�
���!�B��W�x�)Q>q,��)4��9�w��b$�`RWTR u,�I�e�Z�i����ơ�����#j�����|���O�@3�Pr�vB��2ĺ�dΛ�`}�r��֟���
���S�^�Ap�g(�@�"�5D
��߼���Q�YY|�WK�/��,!UY [=�pj����
h�wv����\v����t�\��-n֛U�$G���/$I���ꏌ�� !��,�w��Dd}���˄�������P��ͫ��<s�d*h��/�?�yآy/�>��x�M�6�3*�����j��:V9�'�BC�"P�/M��&�)P�Ua:��΄N�j���W%ّI��M��xZj6��|Q���t*t%t�P�vs| ����۪�E�8�c/a�0������y��y���c�H��5l�D.�![&���d���`Py�����.-4q�K�(��e��L"6�+������Ha�(s��0����������C�"��#l��IW���M(|���>�R�?+=��G	]�u��HP�X�z���1;������qz�[�T�܀/
��OQ}?E�b�(�:Ueɼ�&^	 >���zz_J@mn����q��k����	9C�W)Fj���t�IӖ��?�%_������w��AF���	3����H�{|�@KYk����6u�U��/ɗ��W]�NsȞ�-�h�{��v�����!�|7J���H+;E����h�F�3X���}jӉgi�FM4c1<G�x��@�\5t&��4�7H���p?Y|W��#�R����ؿ>l�rCi!?�A���k��_|*�Cj(5It�3����S�ub%�f�
b�
Y"��u/���m��$�`P���4��B�Q���Iv�)��!%�!w����2�
���� �e+�����لuH�\$A3&���NB�d�5�>�Y5@�m���5x��Jǂ��K�����y�+T�%�>���
�(�0ͭ�La��NE �%�%V͌Y���}c����g<�1g˪�|	G�n��N��x�4�{%���p�V��/Rja�����eo����y$A����[�����'�\\���v}ĵN̟P�w�+tb�~w,����~/ : �S�a;T)�0>�i�e 5�(��y��D��]]�AVe�M;�����J�%!��$R��4y�p�A��9���G�>�2D^�A�r%��zI�&�A״&��@�c�sr���ё��J�~mp<�)����"_�I>�@��J�/m�>��\��2�H��1�is��y=���Q1�bӧ������p�����7tq����]
X�Fժ���lU������	(WGz+�}�IױA������C�36�6�3)&���ėŬ�MZ��4�����͂����{��"N�?b���\^3n�rX]���rX\���"�t��T�p��ɉ�^3��7qD振E�K:{8�7��z $8ܬ�[;���֌�Y����5��ƹ!�̱<*d�x`�����C��Wm~a�k3�ӢCd@��"����))7�loΘ��wO��i��*���~�#M�y�$�����ŖQ!!s��+̭�QT��9�!R`'�}w�^?brRQa�5�Q9+*�^�RD��8Ք�ۿ��:�W���G��CG��˭͝`aj
�>yRqsod��� �\o�
��cs���R)^צYF��օ�zlɀ��q��=�&16#�)�ճ�Ԏ��u�T@C�K�`�D�+��#��R��`R�T��\I��A�X�4��=G��H@�T��h}��i��C�b�����}W�|lH�Ņ�6����c/�rn���0�Jī�4�B�J`W���OAǫe��Z��M�C�әZO��8z�H$��7RDϘwzM�;ՁHp9�]X3�cMԥ��pU�ݻQ](��_�y��.�6�BCF�+=�7o7#W�:"�W�Quf�4�{֟b����$^XsY���S�fy)����.d�-�����}%ӒKϫȸ'�'��J�{p�vS�fN�w>]�wG���C]�2#��P�h3ǚ��P�s�{/1�FF씡2�C_<�B��%:S=~.�s�+�-�+K2->����%��a1�i�p���<��V���0������O��4��͕u��+�P���>I���e�F�eE�bb5������w�pO�Q%�%�*�4�3� ݣ����m�,Mn�T�C)R�4+�(�}Y��x�Z{��pD�����M�H��p�^I�k��(���yV�벓z�L9 u	������Lo�=���4���A?��H�˴ֺz���i�"�.C��]dgjb�i���~,ͅpV���o�n>��!��Z���O��gI���F~J�xT�`� ��b��n�Р̞��B�r�.>@��/B$�>��VòmM��)>C�FcJeC<��F��1r����ZvV�5� �>T@�8{���h+�i�N�%`k�d���i������c��<�e%L�l�
,a�~��H���������3�0�t���^�/7��j~Z�Ԛ�'�F"8�=��upxs4*�x>(%M��y�l�n�	-;kTUf&�D�$����=)��Cc�Yh�&�Pp��K�������v.zC̑PB�|Ѓa|D�����K��`�����_T�rNF�]h�$��9��m��8;B&.H8g���@������&�S#M�Ĭ�VF>S�.�t�0�E��>�Q8П9`4|��d�q!�'�#� Z�}E�F�6������Wݺ�y�9e������@)}�Wκ��z7T�����ۢ�����tr��'����>DI.JȂꎽ�XjO���p3�����+i��R�ڳ�`���8�[��Ԅ�T��lo�{Dl��(X�M�BU�sL���?����
^�p�)^�_���7�@W������ϩ���)�2]�@J ���xx�Y��'+ƫ���(�_��R���R��L-�Ж]F��R(\�������] t��/E��0M�P����D�'w��o��4�&��� \�1w�&��p¸�F�v�f������g����NZ�7�Py��1�zMN�>ɚ���&�9�@��86���fX
� V�����MM�t\y9�P�Ev�y�i{�?rst�E�C��Na�Q`!�|���'�J�Yo�Z g���D�����"e�&^�zQ��˙j��8m�eI��r��zly�6Z
Pt}^��r��ߏڐ���Hi����{�x�0����{��O���[L�B�7�a�
uǔ{3�*�T]������LA����7I��ǨZ���BG��s�.�܏�H%H<��c��������mWw�8hm�X3 Sl_�V<*���' �".�B3�V�vzZ�צJPN�<�����/��soŏ�d���u�|Ҫ��l,;� �pH�]�h�+Ǌg3���4��I
w|[mq��5(� ��Z�*�[�=iD���#Vp�����w=w@>vo][R�H7`D���3���<ҡ����fvpeCj�n;��J!��\��:��Xs�/uv�%'�Do��ϙ{��&Ѩ�o�u��iCO���mո���^3���a�o�2��qP٨����[Ǒ:F��h�W0�GC�3/ч�߰�a�4PP�5]��Y�@�K	\x�s��$�eѻ^7"��>D�u�>f��W��+�q2�����7Y8۲!��������|:�5>����7���G�g��qkޥ~5�coc����	�['�T�}�4��yaP�K�Ա~2&��siK]P\�s}���7�w��@�"������u�A�gb=�]Z���#�������+�����R*�P:���9�Lh=���
'y/'���(�!����2�xn����<��ѡzŪ$V ��q�<�^}��k@��yp@�_s��B[أǅ�� z�>_TƊ��ٴU)���Md�m�7�����1`{f�$uk�XK��)Ue	U����ڌ��n�Зg�E��/�H�x�>��ѫ�b�}!R��#��WT��&�(fL��-C��xc����^委=��&'C,6k���AxZ�A��/�	)�#��hu&肰tV��s���밿��З�<�[����*��R��i���^�����[7=��so/�ĜZً����1�߭X�����j���}��z��=��[N��O~�	%JLD0������$F�I����,�����6��6Fa}�5ϳ)����+����� 2�/�~�H��f_�x��7�M.�������) ?iwUl���ǭ9~אGA=Y���5ҭ�Fo(%;a�ne-���l��	�W�H^����Ԩ$���ho�(�.<[ź���9�p�d!9i�E#Z���0�pG�}�%g�7�ڴ���H���#������k$Y�x���\�9�~��y[lU_��)?]o;ظ������V�X�\�Y嘵.Hp��4�`|%�h�V��ق���j�r���"u����W��A�
@t��k�e�Pi�{�hk��Z�瞙���9�umCZۖg�1UԒ�z�v��7�J�WC�����+��jv�c����H����=��ŲM��иWT8ѵ� �N�+j�O�( ��-���ew��UO�D�LeJj(X}��'�I�c/��p��
.D��m�  U�ܚ�TJ>�@R^7E��u.�W��xQ��(��s�q�0T�?.�%/5�hh�tk�܏�J�CCW���9D����y��d����P��I�g8��4����M�?FF�Y���c1��/�bAiE
���emx�����]���@32�*�ͺJ��5p�Ǩ�`���0وMA��zP@T�P!��m�g��O7=��y~W��V��L@;�P+�b�J�se��EL�_�^�}����RvG�����~�f�ȭ?J�����8�j�:A�GA�oC����f��7|���rw�~�Pj��Fd��G�!�����9��HP�ƾ��H��C@{*�����x�4E��Y>37����J|G?L���3a<�}��n�l��_���/(����ٖ�OP�PU�� 릂'g�)$��~�.�Ǚ� �V�Zĩ�#�͝�x�q`���[M���Q�}�D��"3k�6�����L��59�;��`ڹ�T�g'�U��������A�GG�"���ϛ��7{J?�:��x���}�v���;=����>��@$��|+�859�zq�Ax��cWp��zL�(2q�p��J�[O�{G� ^�_cN���,qV4������DÉͲա� r�W����=�ž:$�j��[���kfƷ4?8yK:�k$�O}�D�Ĉy�F1nb�;��C݇�!������+x��{�I��+����"�[|�K����`*-my��1ԈgG�*�׬��%M��{"x��dϊU�P�6.W�ʾ!�Cn]�^h'z�:��Z��($6,�˺�Tz�&My��<��:�BT�>�6oLj��b=$:���u#ک d�����c�,&˒�I�a3+�M��7�)|�7�v��D�+ix���?�`F�^��3Z��F|�b�7G���}�:nУ=m
y���5U%�r���$�Hu~ޔ<�V�L	���96C� �"�)�[�-���/��P�*8g��޶�/��h���a���` ��d��ځ8�w�͚&bH���hz�4ßoI�3vtAQx�:f!gv7jG��KR��Y+,��ѶJ��������vtw����� �L@��У�*-�zGr+��O�[[���L?ݻ٥�T�����d'.���+�_7�y������0�|�d��*N���Q߶��
�R��^��Y�ʬB�0ln��ؤ���ˏ�YP�&�r�?�����,� L��k(���6�i�c�D��E�2�u���\���F'�]��Rz������������|za���6��&.Kɕ���ؠ�̤%�i�ک/GD]�@�p}�� ��J��:��`Wa�>,L���ldR��^\܎I$���^E�w$����$�?�ч������)	V�ׅ���~q@��öV�ő�+�*^�
�k��|�l��]Z'�	�R2�1O�}�}z������3���@��:̛��&�N��+!�$R��k�<ԯ{�Y�-FKha�HV]s��D,���)9�$�-�U���'�,j���fT�LC�a�
��v*7��IBA�� [��g&W�-�J�.�
��R�_���8���<t~ه��J4�Cqk?"Q��b�W���eeq����_�q�{O�{�ik�[�&�.�Z4}z&-���@O�a��7�&6+/Y��v����#�<D)R�N������A5�#�e�:��Q�t�-�4�I��7<��~��bq=�n�'�Ƃ��E��(M�4S�״����������q�F��zo��ȥ�c,2�L#�|�c2�ɠ�ƀ$�(G��&�K��EB�ֻ�X�~�lӥ��!.YPEZ�V$�P$����h�c��h+�x=�ӄH�L?R*�����q#����'{�ÂJ9Gj�{"E%��bK[6FP:�}P7
cg����G��]o����.�;(��[�#��%���)�d�ɯ�Ɯ�Ot���zaR�?�nN/�UP:ޑt��*(�O]�մKR��� }ٻ'U��N?Gz~��`�k�
(�-�
���_f���3��Jw��1h ��v��AI0�0�����<$05N��F	�>Z �G�=1�yܮɦ�s&�����4}����we̜5�O^Y�.|u�[������My	߆m�W����q*G)�H����	�I��q;�"�"Р��#�"Vwe���OԮw1i�����{^kAk&�#��_.�t�Z4����÷�H&���m(E��Z�>�0c����]-A�5Y#�(y�C�%"^�#jQ��BAT�����A�'͆���Ob�H_����(��/��d#A<rO�43����zC���2��M���t���h��Z�y�˼:��{;���������(<�AC)�������4Xl*���t�i",�;�A8q�Q��ƪв i3���SS�0��9�0� ﭥ��5�k+q�M/(���T�k�����[�P���~�OD����땲֠�ۿ���N���K�[�u9ۖ�~���1!)�m5�&�_�&R�wC�?�����y�H��U5=��S�y�b����<�홣�HM�p�V��F=�t� ���[��a��G��ȷq9b�+d \'�@���7Ò��{<�l�x.���(b�R�b���f߀Ҧ,E!��_{�`lt�ul��y���"�T��l��,� �#��ԜV��L��i��/�A��,	K�o��@`�|M~��8��H&�qh�>w�2�L⮒S�ɽRu�)gߢ��W�+Z�/`\����g��0f�|�K[q�T���Pf�Ϭy��Hū��.��}|�:��9?�������oC�Bd�1dx��՝��N���1#��W�w���Qƪe���F���و��7��%>�?6�`��rM�J�\������$���N0��Q��=Pҟ3��?����&�S?�����T̡g�Gn~N�YO�x/t��/�Qv����B�x�S��,;�\�g�e�dD��t��1q����T�⃄���"|���]��{�	��uSҵ|b����4#��	�f��J�9��X.�G���I�f�X�)~'!c�KNA&'ө'+�[�}u	��9�j�k�2�����m[��0�G��[���|�_�I����.�� !Z#�����,�%���զy#G�=knz%���6�p�1tr�];%��0l��:��*�g88�X�O����W�uX���r���~v&`��]�	�`��������
D��&��p��1�`Y�Ck
 �;A�_��ý�5��ۭ�у��^��S[�f�RT,E ��O�L��\s��:�a(K���VXO�yE�A���� ���Vܴm.��B]ωNN�5c ���U�I�9�f2�$����;|z�O�����敆 ٟ�X��A���`X h�H$ŦRv[f��R?P��=���~���9ߟޫ��L<̚��?�吥l���瓸_!�>h>������:�a�_Y�����2,k���)���Cu�6k"nR��`�`3�?�Ew��;�$����~����]Xon��>O��
�[n����D'��Ȓ}>�W�B����lύ(�ru���L'Ǻ�+<Z��v�����h{�`; ֌�?!ڽ��Z��`^�8���a%�����,J��{�<����t�����i��=6��D�98�.��"��Z'��.zUHWj�}��r�(�����h��o�7�3+��a�!a�u���'܋3�u%	������D?�bB<m\��b�����!��Q��������R�)2_�M�k�G�E��e]Ae;vv�U����MK��\ޤ�i��B�U8ܝ���f��;I��8+��DOp�A� ��I�Y~����=$^u�(�ZF��HY]�D/A��^�/�cr�!�mT#�g�M�C��Fk2���]&=���z�x]�]ø�ZS��I�O�iݖ'��-v�P|�j_��\��	�7&��E��'��)�]d����	.+�zY<s���� ��A����DRp[Y7�#�?��5h��3k#4
o�o�$(L[���S�%SleT�e:	������ J�_%ؚ�T���P�[�M�����O=��W'�� |��\����Ƽ?���_��� ��q��*�(a��ve��7b�e�0K�)���
ŭ���=����nY;d��D�|[A��(�4�r;��B��v��lo�F˫ݩ��؎��8xۄ qy��+Y��̍>�/��(B"f&�n|�UR����`j2����'G-��>L�ʅ��g;��/}cbq���Se��Y�3�M{�$��@]�*��ԑ��Uǩ�O��N}#�N|n�ջ��F5"���i����/`F~ (껱_x�z������%6�Yp��q����Z����8�G<.)�h�L�� ���7�kZ�TB2}��Oד��y��4�����a8v�Q���S��ؖc��z�[˪;���N�5H&}�6hR��2l��W&�2����$���h���͟;�Lǣa��wqg��uD�_3���'����Z��U�W�o�q  �U$��ƛ��p���N';4ݪ����.���5;���?{&di.蓻��=TF����3Q'e����2k�g�G ��[_3m���w~3�zx���F������<߀[ȏ9�v�G����zq��*&�ξ��h]�%]��x���a�:<�1��=q��3���h�Z��U󷕰�(zѹ�g'�k�;�n��(�Ɖ~���Cмf6��9h��
�0 ��2�Uq3 _�X��Ħ��H`J/�E�h�����u���ؿG;e�3p�Ɩ��4��+{w�T��vJ�&4+��˨5� o� �A�v����/�5��
c~�!�^�9ph;�`�N�Q��
ܢ<�[��:�WI**։���5K�Y�tb�����+p�~�N��t�c���J�p��ҹi���r��<ܯ���ۣ=�~���;�D���ÀR�^w�I,���G�v�4X����n�9�lCI�Z����^Eh����;�Z+ǒ	���w�dn��%E��]*o<Ľr\R �1��>��%���t��U��}�J�����T�^���O���`&̸�%vp7?Ix��"[Y��0��h�������M�߽��n�U�2�PkXϴ-�����^Y��!~!fא*������L�V���39v�߱On����	�ʵ��L�i��1��N�[�gMs�U��\�?ͫc&����op	�G �yv��]�z�ν]{�t�>+ �l0�u�r7]�r�S�a�-�j�I��gsMk� ����r���ӫ�u�x�~�
-���7�9�t�y�4i�*���F4�s�u��hpή���D�]�Mc�dd:Fu�
�m�:d�]�:s|>#����SH����S����؝fHe��A����)a	��I;l��������]�aT��n�O��d�ш8��%:��{�>L9q�)ڷ��ً�*Bt���ʼ�2�<�>�@t�C�d���y�zehI]o���q����\Y�	"$���	R�����폔ͭ�{[y~�D�o�!�M��L��nk�����{k��`/15TF�&vx�Ve� a}�<D
����)	Bbptj���cD3,�W�=l�B�B#֑���!ww&�LR暀#e��h���x}�@c��!f��W?_nF��5��?�u��3���3�ٽ�}��U�O]��@�%���1�o���zH{�5���J:��!���g`���F��Ӯ�W�덕������H��<$���埈ߟLT�ƥB<e�$��A�v_�o٢��>�s�� ;A�0m�z��2û� �ĺ�V���W��fX�#�E����^%a��S(�Լޱ�w��R0�N)��
~����ظH���PB�LN"��5B��J�T�o�?�I4��.
ȱh(MU��8����Y�����z-`����|J���8	�9+ןʝ�4>=��2U�r8Rk�~���� �a���{x/i�O�K�E[Ri��I�7��ew�4����D�(/%bءP[ɬNK߅5z�;�D�c�M_G�RocT�yb�ᕅ�Ϲ�͋��%�m��^|<ae1>ss��5�_�`��Rb�Y�"�[a�PXb�����'D"+�&�Сt0㲵3ڒ�2�)V��Z���~n����������%ԯ��H�{��c)	��!a�L��P�W���J�4��ל��	Z��[�\M�.JE�Uy��E���,Il&ςut�qͦ�G�0J1[+���v��*@0Q�|�z��n���<޶�r�m��ȻW> y)��9Pa	\��!J���KN�J��R>T���atN�T��E2����(����s��S]�9}�7=mg��.��}2�ٯ#i�|�7p�/����!�$���N��4BƔ��u⹅Rw#F�U��.���{��%�i��,��Gj�;.���L��9Y;�M�XW��1ݬ�l�f_-�3+�Z(3�)y)Oq7B�,:�
�-s2��z�C�j^_c�֒����Io�����]xYY���s�!.�'l2_
Ih�"MF���b8N��]�=�ho`Q�9�x�⼒|6�C���K���RJg�� ��*�Q���d�'$��
�*,��ɩ$��4u�)�\�xv�"��nW���Mh�Y�Ү������t~��+�]ܧ�o�c�)���} Z*�'�l�RA.q����t�O���[\&�@����8��"M�#��f�L�t���S�}MCr Vx��(S�/b��P}�}���	zM�&����f���8	�6ݴ��k#/�#*�L�x#��v��&�M~�E��xTe��������W(�^��]c�9������1�v�����ո���=pq�l5�V�$�� O�>��_�>�.�2u]U��M��д~��oB+L����v�	�W�'��� `eh�]p���f�$J���F�S���Wy��	!۞� 7Œ���<<sYv�Q�G�P��䋱���M����V�~T�;����|�9����-�t�Sm�B��Ĺﶻ�c�~�p�2R��T	�^zG^�e�����j��\�Ŵ$ĥ�D����h9Av� ߂o:����fX��=�l��1d9JO�X��r!J;����+�+�E�!L@]V	��Yk'Z�*7lB�xZ.t��o,�"��c�� ���f$}���ptn�BP��c��� ��P�q��m��Qy՜��>P�feI��t�f�@5I��Rc!��:�KQ#U�nE�y������g(5���_V7�H�)�jEզ�2�
�2H�0�!t]:�������*�P^RDx���e�
U��7~�s!h�C���.��IX�t���c�������{���Z�mj��z�;�ޝ-`��Ȧ��_��l=|�[��(�\�[�?�ri���1���P3�����Hu�H5�	�h�W��d�+�ֽ�tA�ْ�_�u��9��[���������N�V���b�?B/=���~M�?ǚ���?��O,"[���,w�y�ɥ]�:�����k��b̧�^���e��臍jy���ם��F�`�b�������
��C�WCQ1}�ͤ��o�gM(�y��Jӭg�Nh�'Ro��ڣ����辐!Ϛ3��\�)�a>WI���斵�T���~ {�)x)Y�V����#�� ��!B�v��Q&�M������US�%w6H�=_"�����I�Wӳ=ʻ�x���\�d���좦|{�A�Ճv�`}��w5gݷ5	f&�nxE-ݏ��6&Z�Y?���C�/�����:2�֋am�.�#��co\��?���k%t��"j�s�x�Bԏ����ay��{��n�#���rPʄc	�JN1�T���@��S� ���Sgl|9d��	�ˈ����ane��u#��%�+�D"�;z>��S�ր�H{�B{ۚW�ͻ���XWC�D��Jf?�͞��">a�R7R��Khhex�y�Q_��̣��|���-@u�Y�����%X��[����i	M�8yrc��y9z�U^aQ��r�5>���$��xI(C�.���I6,^��������P˥u���b4d�Uւ��瀣���:/򯪅��o_�ҡC��K���J{��҅���
C\;Џ�����P}i)y�P`��Ocfc��=A����w���G�D&p
����Z����h�ψ�vh[���L�0�r$���3�oڀ��>�[�!�G���b�w�(���t�2K��C�Ѫ�͟@j�O2��l)/ONM��g��1� ���\����:�R+:�@�(�L��B<(ћE�n��m\eTl����MO�XE4R��`cA� �H��� ����
t�(D�WpM�.�~R���C����u��Wu3cZApPɲp�	��e]�F	wF�3�^:Q!��y��nF�gS~�3��IH�jTе��Ҝ������=Z%,}�6���g��D�X���^k^�yWY�� �+�%'xSA|SR�!�g��o�B�3/e���4djp��/@UBUel��V�mt�W�%ƒ.桥��<ƶ/*�%_4{H2�|4?�?:rbp���#��^����{���8VND�	(e^�\&��x�0���bS`'R�;M���XׂpǮ�@�Yg�d�*��$@r��Rk���B˕��-d|iu���]��X�+�R[�  ��悹O'Uv�������(�xo@��%U��u]\��%j�8Q��ټ���U]���Po�.���v�+��2�a5�0/��� 1���iH�'����훞�E)�&�����#ڒ�����p6�%�|�3@��z��޽���<�D�V���T�Î�����99��a�!��"VK�ɝD�)�X����,񖾼�Nc�  G�����G���6�3�\�&���ch��_�S@�h�f�!C��Bo�P�Y?Mf���S��^bqثE��п��ݰsl����Pd�ǨTr�����y��M8	�_~@�S��|��7 �w��t")��wư,�(��>���VeN��|�բ;�GP���?H=�@~�|
�/����k��ʖx|Z�M�d�� Q��g�����ПwH�ۺzR317+ҁ��0_��:Ƚ���ϧl�R�r�R�W�l��S�M�{�7aa���tr���xe��cⰩ������^w�5HtUnͫFV<����A����2�SB�v$�(P���
=
�H7�r��"�"�G�W.$��:��xoX���{h���v��(B��ס�"6�e���^��R���o�i�vC���4�v[����3�q����?�a�������2��(OY�!b���DJ�������c�f���t��t_��M��(C�P�ҁ��f��n�E<'`N$���R�a�'įk-/0�=ƿ�{�u����\�F�>����H� ����!�F��������/O�U�8�F��j9I�=�o����rk�#��ĸg/A��#��e���49	�F0����^��g3@)��	z��Q�}t�ݾ��>d�m�,n���v�5SAS�؅|��+%�]�E�q��w�t�xX�ơ���prSO�U�Φ�RI�1�B�|��0�8@�i��A?�Zs|n`Ș��f�a�x��
	�z_h*�2"� kp%b#)���`E1����Q^K��ML<%(���+C���g�T��z��I=��B�6�>N��L� �5�?JQ������a�g�xxm�3|���UFPW��w��`�5"��ք���;�
Xo�~Nm�����PdwX�hl!?l��b�,(�w�o8'Z�7�#��@�؊�-���RZi�r��j>��_��*�qt�	$`��6#��ܓ�?Lx/\�j�^��9#p�ʆ�fJe�2CܝJ
�B������>aGzT]�x�;��l�!*:�f&q!#�
�X��*�L+���G.�k��#r|�R{���;W��2�uGi�7�&~B����y���9�������T��p;k����#U��Es�%�=,���B�V��n���b�E�a@�?��>����X�w�M�H3@��ڬ�fq,�<�#�}y�Wń�	\l�9� ��װ�գ,쭎(�l#}x-��?~�-)�:**���q\Fs��C\v1$�.�\`�$���4}�z�9�7
QU�a�r�Ϲ^�U���;�9r]���`��v�qx�Wp�eW�N�D���9`��VCx��6������6b|b1:.(	D���[��,"���w������ ��#=��,nF�S�-w�;'�&	�����c�-��Ա?�ޫI���q���#Fȏ �&V����M0x�u��,4�zL J���0{o�Kb�3C��fvsA��Y�Ĭ-��9���䪧f/�N�����4+$W�;����Q�`�Mл���� �@K�%�kJا_���AE�ߕ����C�i��\�gĺm��˷����ˀ�3�h=������Vр-��ts�
�����Z��5�|��By����Ɇ� �d&�+! �:�c19�F;�q� ���i\UҞ
8��8]��%��#T�p �a#G�(D�ɉ`X��y�p�g�Y<��j]�U_Q�8��H�l=[⨀k*�ZW����IwWE��c��%#�Sk����	�c���E+@|T��z5)gY���N�{OU�g�@2��K*Q״�Ų�e�Esa{��b��#�"���L���(
q���YH���^Z&���`�ӬN���"�h����x9H/ћn���w�hG�B�j��1���>L��V�EO�[j*�E�'�,c�d�W�$�^Jt�I���,�Y'�}�̐��gb�M�V�s]7lD�M��t�B:�1箟�&��d��;1�.f���T��2�8�%���B��UcĔ"Ϛ�N����>ܼ�(��I�G��9a�mf�9W��Z}��";�}�0��.�W^߅��Q:j0q�3�h]A��E�5�Z٘@J�q��O�l��a@*˜�Ǜ??�	0���C���s��dG�E��W���I�uUJ�Ԍ&]yM:7���Q<��@<gok��G�3�AW�Ÿv��[Rl�ψ��ĳh�P��������r�4� L��c7��6"�z����lk��q9_.	C�;ip���nh|�7HI��Ĺ�	y��~�OB�Y��_*c*(̽0��,��_:�=>�C)�^+e G�v(���=~������P�ym���,!+�î}5uX ��B�ne�T�Q'�[��o5:�K�.��(�z�V�i��f.����t����HWK�\�S�=}ʧg��ܮ�jo�e�#��ٱ,,���Op&	g��s0�.D�2�mtZ�	�cKU)Wɥ��ڍT��L|+�7Ĵ�one��3=��:�?�Mr�i�b)#W)mK%fǡ�g]���j�葵��i� b�&}���D�������7��	[���cӬ���:�r_S ǧ��kvO|� &'XZ��;C��Z"!P��H�D#bd��o݄>����6]��wwIX�����S�y������Yo������Bm��)[z�����xw���Oh���+�r��S�ܥ�4�f)�iu(>aAg�]�K��	�6� Gؑ�O��I(��_7�I���x����{u��hq�]�xG��;�>f'��#{�ׄ+��/4�w!Qւk5�=r���#&���ۄ%a��}�V#Ѧ�sg'2H�� P,_�,�� v��B~=��?�@�1��܄
Ƅ�5#$���d߽�(i��Unǂ:29$bp��AS0�J�?y,�ͳl�98��7�5K������G*Wr�.{��h)�� �9��hޒ���fسǹ:��g�E\
�opct+�&J�L�3�};S��H~�W%y���
�[�y�ſg�ap�����)K������,�_�J�|.�tE��i�v#�auB�4���"����	־��OA�x� X�h��s�։���~(���(�LQ�"+q	e�3�OݧF8-G0��u ��1L���r���r���6�K�����~A���Zf��>��;�{���9�iK���Ì;�4t��Ǻ�3mL��0�Q�2��+ܱ
��HI��$���x�Y�������0�����Q����������P��[�G���Ĝ��L�>�7&r�t���a.j�p�>�=���c�9�8��g���O�M*YJ���:V�Ш<DK��?Ff�����Y4�M.f��FL�Y�!�<H�) �*3�ἵ_�^1˚����el����s��ށ��t!�w�6�"�|
��"��1���ִ٦�K�=4˲�_�(�Sd���p�3X��)�M��G�U[Ʊ���.t�������I�*y�&k�)��C�/�B����Ѻ>�.-N�1o��Ο7�"Ӓ���ǰ��=-��2ܹF����Wyٜ��lj���Jλ�a_J޼(�����TkcLW1�*��,���?��g�|��)����ET����i`3pT/�5⬙�@З�1/mS���jѿ�8��?��Mɟ�H���eN����R��ؘ�x��
�=;?�����ʚ\aյ����XX�Bp�����;�e(:����3+xǪ6|y�D���K��L��dAL��_O�ae����@�W�h/I��<87�<V%D�G�3u�rn�̙�ݐ䋐Τ��� C������H��W¸�w��~��}���}�TK�!�_V�������~��;�gw_�=_ǜPO`����.7d|p/��q�b_g�1���&���v�Q�?�/0l�'Š.��{��;N��`��S�%��vD$CS#7�ȏNф��@-~;��T'�T斺�'�NOl���i����!'LG'��R$n���U�?�Xm�(m(�ü��nH��= ؓ&y$s<�t9����M�3��5�gg�N-��@�����.9�u���Dk^�+՘��bz���%�V������E��0Ӹ�^BV��\;���.:�1��XņhstwPxB<��p�bͅ��-��0,����pr�$#	��P@.���8�>�d��$AM��:�#�v�y���5���U"u(���������+Z?+{f�6ȟ�����
m+��v��8v]w��%O�)�`3�I��k|���:�R�/���cN�������#�����$��#gj4);�ύe�:Xv�V;�}�%��d�6}U�����v.缯�/��E�Ҕ�������L+�[�I�~O##�B��V̵2F���׏��Gp8h������k����������QA���[�����%.��%	[Q�Ej�!U^���s�Z�Y��R�s����4���q�����p�&OR��L�6��L�M]E��ُ6r���'�8�HSH���U���!q�fX�F>`4�n�|
�5gުy*��H|uӴ���V8l[���)/��+r���^=��ߢ�km��I��:��c�?b,��:ڢ�IҀ�	7�(b���Q���g�}�P�h�ݸ�m�_q�^�b�M�K��	��l$,�\hu%?��{᥾U�+���@��u��`�,��L�5_�n�@��.��!��W)�S0�k�9זf4�?9� j2)w[*�# �"�K��o.M����T���WH���3db��:�	 feÒ��U��D���8�x�(o��0kp���a
��b�교t�R&C���gY�{�Ă��|'��qe�PV�.3������3��8�_'LY����Լ�N��ԙ���%��( �?�~�x�G�Oٙ�^��5�LL�/}�0t��q)M2���S9v��\�/��<M}2au�g���!��I�Y�q��!N���  ���fF_�C��YX����P��z,�;⌨_�; �%肻�O������6ߎ>�V@C��S���[�L�of��ޱ�T��+����{!� l@�];q�<{���e�,�{'08��Zj2����I���4�.�%m�!��{�u!{q�I{5:XL�O=�!��!�n�e��Q�G��2.�F|\$��d���>�	���U�!ݼ����Q�ۙ ��,��IF�k����3Rх�}K��P^DSD�k��d�������x�P�ٺA���VK�Y��*�pGU1�Lc"���e��p���F�$o�C����.��������{r	l�N-��(P�����x���(<�L���þ�y���t�:���j����Ţ俾��cV�ʠ��Q��>v�)�|纕���\��K�<V#��#�V}�m�9D5(����R !�cmms
m���_R\|�q�w���:�z���a�r��q,/�Q��g��vW֗�rd� � ��$�'���Ժ.�	H'.V������	q�4g����!�ە؄�=�2'�\��ᒄ�Y�l*����:-f�C>i��yK�,G�$�TX��������Ɂ�?�l�G*���RWe�#1ҔA�	��+ 7�>� <��c���/�8@cz�ŭ��[���2Z{%CX�!�BA��a�~��뿝1�5�Hb�=l]j�qIv�����J���-��<��1_C4[$T�ލ�Ҁ@��w1�J?>%����g�H(h�:Q�Ӣ|�_x��� �#��'3\�Z �w9��.5-���I������M�jv�r�A��m��P���~F/NV.�m�'�8�ͥ���,��_GP�̲�`�J\ ��wnM����2^"�W�B�v�l��ϛ����e*��{a��w.��=�ʈ�%¸���Wq���|A���������8�k�D��wȈ�q��=���� ~s��
M����zv;Y��p߼<��]C:39���ڤAgR�0���ꋶ*sѼ!kD��F�R�h���)�L5��e3��G*,B;ݞ8S�u�1w#zՁ�V��A7~m%�	Ñ�?��[w\ζLuMp�4T�"���>�O���~_MR������s%�B��|��h��!�hY2q���AA���x�5O�͛��B�E�~A`gi5`/\{���^Y�n��U�,&�ꯒc�z�V���E0ָ^�b��u4�T._+�(tleW�(�8_\�V��9v�vx)��FR�����+�
�M���[�}�v�|ݾp�B���ucp�L�B��Yiy��C�K��4+k��"4}�+pN�6�^O6-��r6����"�A���%�G�H�taA�5���]%v�}�f@���6��분`�����#�B3����ҵn!v�9w�|�2]n0wJ�m�XD$�I��-5�9��ɜ*����
����Զ�+q@���3i6�]A��7�Z����Х�a/�(��NOG��dp3#u+�V�j��*�9���}�.ȑ��'u�v�W}B�Á� ����WvX����}#�k*0���+�0?���oS!��:��o���~�(���k$�3W+W���A�'>q�13��p�D4��G�;t �'�2�ۑ��?���*�0Qf�ϙ�PY��*n/+��ԾT3�,p��,�#M"0�U����L�S|��#�ےA��-�A�+6��;S�]AfU�j
xY�fR!�Qn�>������{�duy�K�t��2D��7�?��aoĭ{%����m�.\K7,�K*Q٠�:sc�&�8��&=�R념B*Y�d���|e0 XN�ÿ��S� �Pfs�7u�C�B����w�0���lm3��&�J����wGhi�e�v�g:?����;y��
^��4�{P���T?�a�%�����U5���r�Ov�}���y5\�Ɍ�@H<(5�ԗ�c�&
��r�m��r��O���q8�6Al��gA]X��2��G(ۉ���\m�@�
����\t�M�b	�ʏ�rص��s\��V�
Q���+���T����j�Ǔ�aD�Q#���F#k�Ȫ��U؏���P ����GGx1���g ��\�����a�͐���X�K�7��SQ�6GD�=T��B0K`�X����r����5"�4�M1f,)8�S��7���s�]�]�K`�e������&}#3Oj�̮X�B�����A�y��?�|�"���UXPIi�47f-0����i�+m-4��F���=����И݌����[�O�n�S�s�<)ʊ�N��V2@mqW�c^5l�%K��Py��S�]6�[/��[ ��b�� Yl,��K�5��.7o'X��-� �p�蔝���9���2�ZM���!x�W���i)e��ea���JfY�Q�~��rXH��I�E����5<���8�D�*��4���:����ob�\
U�*��7�
ȁ�f@�U�ŷ̙MyG/\���Ԁ�~�U��İ��3�Q̎�sG�$B"H�0�'֥x��p���o�J�����zX@�1�Of;���h�3��nƹ��6�
�Xo�(�WfF*�"�5(��Y�u3d�S�&����>ORp#m�(/�Z��Ɨ����q�lk't'i��޼��;�c�f3�7��ӤF�RE�H^�Ok���q�-��c���Ph��:�����Λ)3ٍ����AR��T���|D����<j,����x�E��ŏy%�[�a��e��1���a]aR�$�@e�KT�hW.ܵ�͎����#���Y�%��h��`pG|�����V�v)Iދ�N�e=h�9xǂ�l�f��v�,���l)���]z+E�j��2�'_Q�ͨX.��Ypup4� F �B��� ��tv�)$��5e�ned�J72�p;�����;���F�Gi�`\������<*bYq�Y�"*̊aH��m%>�%0(k���,
�����E �+�'�q�*�I}+6�H�k��k�Cܕ �,�7�g���.'�Xs�_�Ҍ��0���k�_����/�8�;LCl����ɛ�:Yf�,�݈,�v5�A!��l�u��6.�8�R��o��;�\V�֠W��ӜO���u��}��S$D��.N���ɡf�%��v;�1kZ�.��q���6��ʭ�W�_E���(��`_֜�������ur����8R�ϋk-��k�~� ]�S�$@����ұ�A�'״v�	2��s�"�� �"��t�K���ݹ���]��/qjg;s��_� �������%��j�J�"͝P+j(?��;�f4Z�f� G�T8�� դ�֕�fM�'��I��nc~�`�m�>��=]B:Wu��f=j�*�H�f�#�h�0kp7�Y���~�M����<H����F�؁S�g�)��h�R��O׀ڪ��1?�<�O�L��Y�{���H���O}�t,1v;�6PD }٨��$�A�8�Tb��A��#��.g�q"�j��d
+����*��00T�Z��f�r�_@8�4U9�X�V�QB1�ΚV'iI�G���x3?�$8#��� ӽ�p3����"�3�����k,
���l���K���=Fzd�֪-)�����w)$�XA}<���5�H[��>W��삆(�5I'ܣ�9�=� �X��z�D�2��>](~VjM�sm��T�iJr)��$\<������ &y7�L��v��Yy�'��*eX��4�����H�����v[��d�R��Y�S!����u&"�g7`8�<m�lz�.I�:voA�D�5�F� >�ugn��)r�3kK� ��#,Q}İ�3|�����`�/eC��x�8m��'۸��c�;�=�ҵ����o���m\��9�w���P,|�.�[j�����������8��lJ��vK��#Ԃ��rjg�+�.���-��yws^��V����@o��^����lr/~u�m�f&c?^]��h�J�.����+�N(Q��p�|D7_3[���r�J���~�#,K֯6`ɑ�ꈛ�p{��/�QQ�[�M(:qWu��b�A���+�o���1�&�֖Gl<�����̰k����B���'���� ��a,p	��ܯ*%�V"p"p#�J��a��{�n�>��C.����m�	�����t2��� -�v�/6��ʢ�Q���o!{��(-s�Q�I<���ַ7��$q�g�`L���k=Ek��������E���}A
}h�W�^q�/X�R����`�'%`P��6;�rU:�LQdJ�:dy�fw�vI�9���1h��N{2L<g��'g���u޷��E�{%{�*��3���k��W�5e24�MO#�y��C�{�����l4�xb�w��q��b*�FB��dg��Ed먿~����MY��^�W��W�#d�P�]Z��|�!`Y���:���"�L)0��ݱ8�C����;�����N�Ű]�8y)t�͡ɀ��"r�C�Jb�ɸ����rjk�է�#�D�|>��=�z��3I���H�qn;���_ڬK�F��oFM��sN�?�U��5B-�	a��p4�;|	���$�7��c�"�	�M?�c�[�~;�<��RɌ,s����G����V�B��|�M��*G)Zâ$m9����HM���%��;�&B|���'UP�+�:z�̱i�σ��4h���惒�Ij�D� ���3oyDllD�����fW��F5�����q���[�3w�ݙ�Z��3��fY�Y��<i��w��|��^"#v|u�Q~��ޙ�0������Ϡ����S�VCGHd2����8��O,�4+�jZ��x��R�(;���"Y*�c�?b����'��mR;/�;���"�(�ck�E9�?-l׈��ͮR����jb? $b�v�$龤Y��V|NXC���79��Hm*���\^YHAT;�]?.eH��a��<��=Y����������"z��*�X^]a|i�E3�8rc��~��J�o|��EV[fgP��:
(�}Ņf$�§Y�[W]���8��0� ����2�J,I�����9����m$�Oה��H����[�=���j�	���Sd�����n������7[��Ki*�tW1�gd�ϒ��Cf��P}��%�'E���vS���Ef;6�Z9��dôپ��y��_��p
e�$A_3&"c�H_ߐs����/���]0�Z"��i�����B��0���l]���:{7��x#n�j��-~!��@=���*��	h��\�ِN>	��h׸#8h.���!}ԢӤ��WBq��@
%#�
���^��XϠ���ކ�<������M|�	L2]��-|?X�p����C�ŗ�����D���ld�c���R���ݢ�񵲭�>��1�KM%�q�BV5�t�c&�<�b��E�a�Hdנ���c��RC8�-�Ƃ\����TaT�.�SJ��S
;�*©/t
;:~Z �P�w���bE$�f���~��U����_4䂐7�W�	�%9w�ů�@4��p�R�P��[��&��R�8�C�����]A�����>r�����g�=�8���� 	f�b��b9�Dh[�Rm6`F�0 �f�:��q�?Uֶ}��TʸB����g-$���t�)s�@v�L)� e�Z�=?A���X+��Q��'�F?��fK?D��>��xÒ�~N�("�r?� �����2��e�gu�t�z��m����l��6s�,_���/� ���a��M��^��\�L�_
��	��j�_���.d�&��X�n�G��>H�P*.�����UO'��t%�N<����2��I-�!���O�����N�� զ�s��g<qc��L:�����	?.�o�D�E�4g��;C��g�(;doŲ��ݤ�ai�3g��B�2�ݛ��:���ˈ1� ���d9p��UN]Y^������I<����*jex�S2B�I5L����Pb[)��?G�Q�k�4Z��1w���\D��Hf�<�?��jb�;�k�
ښl�A1�����"˔��6�h��	|�S��}a�kJ�Z��B�X�k�Z�n��~5[�)!Ýh�(����]����_�!�������_n�*���tV_x��
��]�8�)F�&�՗�.µ���������f�N�ph�������K��1��F�	���r�L��A���� �����X�.R�$t����<$lW������"с�}W�՜A0��O	��!wd����x�R�U"��6� ������>�Q�_zg^�F���F?���h�����b݃���6 ���i|e��8�:�LR��9��AUrL0F�/6[�!䄑R�c[���Du�*��b1�.�=�9�a�D1XI���'# ���!�g�q5ᠲ�����Dz�ȇa�֛���u�a��`͞(@~���\{ɗu�nf4��Ψ�Z+��136�'��R��#i0�PTWkd��{��k��q�עv0���b��u��r����̕,��Jh}�#I!^͜��`^U�raq;�Mt E!S���r��Ot��Uy8T���g�!�K���p)EH�K���1�8��>~�������R�}�����Irg��)H��42P/�XH�cB<������0�3y���	 &�6��Y����Ѫ.��Q���~�'���'*�#54�����4-{U����"�%�o說3�Y̌�3��sk�O��dr�RR����ua��_�f4��P�����Ӏ�?����)���6I��b��p��_{�
[�\E���:fִr �����!W!���I�y`�*$c*{�<��oc�� �4�N�)�$T����6Ą���dE�`]p�Q���9X\Ƨ;"+}�il���������%�Ziz��eJ��Z�^�D���d�Q7#̝�ObtBj��BrG9���)[]���ب�5#F>�<�`�7�F��->G��R��X�[�>p�\�&���*.����)��~�>�>��jr�j2u�w*~�9����4������3Ia�>w=��U���<t��O�OԴP�+�m)�ڜe�&�rxk�#�]��I�Դ�A�m�� �|�� yΔ.��*c�	<�Ak~�����鬷{��]p�Vc�� �����ϐz�(g�YC[`�d.��}f$��<6�k����-��nH!�_�/�\`�h@�w�_Q-x�qQ�+�cAP�9��v
�M��{{lB�	:d#QHpy�N�tiC����d�3��$��S��xd={k(����ڼ�y����%��Y�I�4�t�[���}J����P��a[d��g�;_�A�K���<��F_����XM? F�d/~��(�l�Y0򟬜�O����]y�i��4W8(��^AQ.t\�v��N����4{&�!$����9s��7�\vyewE��Ҿ�XĀ�*`5���Tȏ���S�V0��c���D����r�YDMU6`y����R؇��[�|�H�0^�&��w�f�x���gR濜.JWu{��j�hsY�V�W@��\d��w�,VӋ�@��x���,��qsч�(��A���+8�InR֔�F��<��Dը������M$uS����?<���2�P�Q���� ���с���1�ۨ�L�����T�����E�2��$}�&����BJ�� �ڡL�}�Y+n��{��h���>�5�����q�\6q[��+�(o�1���z���,��/ļ�zM �oV�KVU��%��_./m�:@�	��e����h����)���'�!���"B�������F�gk>�����k�nLh$�Z/r�����.�~Xӹ�4�A�g�k��4H���b>��mt1��3 �4�&�.�wF���̀�vA����'�i{V}���m�n�?��5���p��â=8��Df��G�T~�<	����� ��2 s<K���y�>�;�9�V� ���|fDe~�!-j���TP7��~�lb�Y�_�@�2�׳���	RWo�$/2dJl�J��e�c
��%一��~4c[&�']��m��#v�l������Q����=FG�T��萙SR����u�`j�hÓN�y`>��mZ�a���~\C��r7����|�9����8jLWd�B�Rb�7�	;������T�Q��
m��{[��ǅ��	.�$�{ i*����?��,��F�eΖS�l'��Z���$��F��G9g4�f�Cz�C.צ�0��Uqﭭ�N��'݋�~�s�,��N[s�_��nQ���h�������?��m:�#9�_o����S�}5y+s��� �ة<~��O�+�[��l^ĩ�M���">{��g��ij����o�u�>-S�;-�F?��}�TRB�C�6����'��&Q@B���|��L̞D$ǔ���L>}��Et���g4g�vZJ| ��B�X5��܋cFE��;�atƉ]R�r�l�D��gD*��
�# A0o�P��07t���w�/�V��s�љ_/`�	�,�K�݈"�BL��ą4��H�Ā�c�" JN����U���N𸦦�2:k�xD��K�6ȕ��������A�J90�#*'q��
�3Z[h��.�k�4P֡[��֑��e_[���.�����+�����xuH!�nm��IP�ŕ�Ll�6�4D�"\V�V�J���%=.+��f�q/��d��j�����8��A�\�^�n�dtS�Vw=��W>��Y�� ���r5����2�����L��c���:F�� b�r/I2,�Rz��<���b3�{���<J�����TI��i�b�SI��4�b� ΰr��m�<WA�X��R	s�*	�W|�s���_��a��C�M�Rp���a�״�olX����8��k���ς��9�,���e&��V�Z�"��:��oZ@�_/y�{�J1��=�9�(l��~�)�8��c3�
 �̨;c
�1�h�e��S�EP�j죶�!ߒW��{/����#��A7d34��6nA.�3��ys��CT�S�x�2ଭ��"��8�#��L�b(���ۄW��V;xX�2<� �Z���	8I��ƍ,G��'+��i�t "�Ƹc/�>���e�������M��A�;���랟�4Y6)^GU��e��<� �"�Η�vܱ��fN�t?`c�:>��e>������[B����߀���QUǀ~���>c�q�;]���G�9@m
�$����'�jw!�:��X���'f:g�H3�~#.�_���<�ľ~���C���q4�!�}B �S�,��9|	�����Ϊ~5�A��� 
g���V��'�w�C鳤{�~���C���l}e�������k��0��	M%]�T�j�P�2v�Ғ���1�T�W��$�����fؔo[=��|�4/7x��jc<��[`]���!)O��]"��Uf88i��||i�=Z~���ӤmW��؅��K�׉�z=�ʛS�0TtD.s�
a�����I]0���;��:�JXp|�ɻ�.l��<T��I�5���K��b�c����G� 2e«Pݤ-Ey��NE�K��}�qg��E��̨�"k�j�2E��bWw4f��*�Rr"��;�H�P�
�W��H�C���+�l�zv9�����iV�1���>����R4
���X�|?�m�j�����`|�di�Z_{��*��ʖWr�ƚ����@D�W}��a�hG��%W?�"*{>N'F�m��8�m�x&E�ľg�G:�8��|��.����;�~A~�"���ͪ�� ��床�����a��¥�@1B��x���yoK,���'����%�L��ߚ�^X!�N�Q	�����a酌���Y�౴�pQ �Oev��U��طR,xF)V,����9���j�'�^dutK+L�"