��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�#&��#�RWG�a'hj�hD��h�\�\Ʌ=��R�^�} ��@��z9�|b�[m�X�7T_��s��'�m��#Ԧ�P�_B���������
�A�l�9{U�-�u�5+#������	b�J�A�`�6~ʁ*%�E(�x�:5��]z��j?*���GA�m��`�x�C�������QY���h��z���.����O��f��#,x.��%Iu�
�n�S�p�NU�����=6k�������i}*�2��G�)Δ^�F>�i֍@��F��l"Aj
?�.	�KGeV�ۧtֆ���ȷ�!� A)z�+-5���ɉ��aR��`+��j�Z�E~w����jMO�hF��ǟnd�I������{p;*SFN BT^��qپ�ʞ��@~f9K(�Rg��VfCm}������|N��.*�t�a�ѣ�jrs6x�h�{����u����S9�*�+��s=_&[�~��t8���R�Y6��l�?�f�S��g�p9w6�����*�X��gi#��%�M�j��('"g灺3\���MS%R5
��p��/O�B ZS�F���r)������' <9tp�=J��lZ��\>-�C�~���:z6|g��4�u��9J�i���R����(��6��'Fj���L�<w��<L1A��pD�w���F�P�^Д.G�G(�ޭi�t�@٭|�2��b���<��5�'�� %Z9R{e���t��+��eY�9�\�͟�E)���/����m3:�#	���RR�_�H��Z�z� ��i�͒��1�M(6[-�L/�6[ל!)k�_y��Ŧf���uBɝȣ�X�~��]�`P����]��Q�MP�y�ު
�NHꧢ~�g�-���H��EH�F�Z��W�> %�N�FAw���lQ�~��e<��Y}8�Ļf�Ic=-���,�N�d'�՚�g*�l�G�k���f��g�_G'���'�J3 s3J�K�"Q�f��o����^j�]���WНn^R}}s��;J� �8�;�뺧a�&	|�8|��v�mI�����%0���8P:�4ԛ4X���XBh�it	��m�@mZ3{m���N_(,���G������{���b�o ���阾+�3�`�����Ë��@A!&�4��Ї��l����1���v�'*�@P�5�v������9��.�l��?"�\uw36w^�($���kk9�c��)�m�:�/�,�3��^G*4ҩߍY�(�Z����9�_�vj�]�ۻ!X�6�E�vUN�`���ߑ��w����J~�����,����[ԁ����T믪BN�d[��_6f'����Lאk4ykɇ%e�b������yX�
��q�f��.��ps6��)�?2+���;�n4x
�o�el9{���K�γig� u`�.���(�Xw"3�
d�߰�噼�!����� �oX�ayؒ3qJ��"�ahǘ�aظ��qH_X\���y�"S�$�6�e��o9����<h�F��!n��ő5 G��`��@f}�����_曖m3��@y>���c��I�!��K����7`p�!zw�����H��DF���u;�
'v~�Z���4\?V��e{�m�3D/����)Jf�g��W˾�\�f*Y�fi��UjG&3\�~^���O&D���"�e�wOP��`�Л�L0�hW�0�&C��L`0��D4��M>�U��UNئ ��u��+�o��?��_����!G��qO���X�%�Y�{���:ЫN �	H3P
MuD�l��j������-�N]�r�/O�nD����=�Ƈ+],�b�B��i��5��+��:��gi.!"�>�MD����>l�`H�v���
9�r�C2l�zs[1H^�QѴ)!�M�X��P�j��U����,�S�X}�����JU��q���*=ߢ��Sgg]�6*uo��HZ������`b@�<���	���kt��O�|p�A�9�S<�ƈ���s���nBw'nb�����2N7��5_�O�`����I��T��<)��yc<!�F;�&�TA�Þ�ȑ��E����f�E��+�Ӧiy�hO��§�~:"�}�Bs��n�����6���>�<�%�M����c��d�;��mp]�K�f95�T^�=q��)�,�t��D��+x���EqAO{S�'��R&�>�<f��+�iu�;q)j2�cH�b�]gb^s�ۮeӤ4ӣ�f$.<��(�3hT������_�����	,\�j��$���=#� <�2N�'׬鐅�I����m�w�=��e�)������]|���*�k6o-�4�'�*�o�8�/P�4�,��h!G&Hٞ�&�#�q]xZ}-t��w�9��
��t^.�>��G��ؘ�_����Fg���q"���/)f$TIS:��Z��.U�dv" �H��Z	��+}�}S�1u��uYRv�N�ʂ.��8��c����3;6 ױQ5 ir�Ȁ���*:)W����@]��U��sD��6���uG�<�4�æ||�]�k�{�����G��'�u25O�eh�4��M�~_�~�>�u��V��H���p�C��oZ� �Q��of1���aW<�|&�����]�=�eB#b��ɟL�q���V&闖O{ �G�3�$�Ű�Pu �.��P\h~7�S�CK��$��0n8����5#��i�=���bt^A<�?E��X>?U����s1f���Q�z�(����a^^@��a����m���Iu��oXe۶NK3�euv^����
v���cڨnĠ��� 5j��T��2^St&?�`���ݰj�'���~&�:�꒤���J�8F�.R8:���8�M�b�C(��`N$ЃBR��{�^9ؽ�����hV�V�V�Y���hw3N��Ŕ#�2:<���`�~	R�ND�'�~k�J1(��&3�%���{�d�cQ�=����&b8'��N��zu���I�cE�ݮ��#�f�Wx���.��%W��!7|����x�����HT��RP�G`�[+9�SS��&�������I0�,ʤ�A f��A��� �#�Dr�,-立h�xP�W~T����Z���DǘJ��ݺm���r&��b������)�нA?�+Ol�k�o#�U���&1�\��2�����m�t$��cMz��a�3>U�
�I�ķq>�D�qG\X�gN��d9KB^�%!���]W#n'�����9��E�]�wȥOE����
��>�"f�Գ��q�ѿPp�Se��i�
3 >�ȏu%�~6�"e˛)|�45'P���_{j�dm��*�a�(ƪ]�&^���<?9K�v/ 
��r��TGUV�f�1�)YǘS:Ƿ�Ӭ���th�6q�g���+�,� �gnrɣ�SG�S��ŝ���VPk���w= ��O��=/��1���a���p���&R�N]Q'�&^����GB��o�A\irI���g��>>�S#A )�b���E�u�x�\-A�>5��~P���{�ғuGu�-f��N���0�'r���J:��W0����g�ߥ��zР<?W [QTl	���^aҞ�z�jH|�ѮO��}g�}0�u���$m�$���cJp-����PެReD����W Az!�U8�	���!PǞS/�9C��s�9x�*A�\C�ԞdK�#�y�z�_r >]M m���U����6w���H�qK�4��϶�u'��=s��\5�����-�e�L���h�[��Z���aLG\��t�J����A�`�Yą�
 c�5^0v4����G��pe9������I���$�a�(�z���DN�������Z6:w8���:9�<����Ä-�%PĬ���iv��g�	��\`}Jyk�$�
���ð��!�f.�k5u�����=QPR�����2=ܵ��j�F�������a)k#�,��-��DU�&wY[L�XL7��� h��+��e��f�h^����a	(��Щ�v(�1}�Z�IMT2��}'{��:��f���'Ms��kD�]
�5��I�f#������4����O���q���@^Җ��n���F4̑z� ������2?ǪE��i��g%zI�� ����o�y.���Z�W�׹@���:,���P�yQ�$��ԃ<�`K��<B�S���ac�Mm���U���l{�M���W�U�'9����F� ��<jod�P7I�b��ڝ��t���͕������ݪYcf*�����{��0.�Ȑi��A5���Gr�g��K
��<UWӖ�,��n�H�T5��m�f�"�p�p��?�HG���pal ,S/u�&o�K�]2�,�D	f݉N�l��l�	&
�U���F�A��5���F�$��0�g��m���_ĸ�ɋ�����$[F�:g9�;O�e���k�7�"�W�>|���/��ź���,����au�^W��x���������e[�VM��P��a���ݖi<�s�F�-�x�!0 �ۧ�1�-&`�'�R���or�ᓃ7�������7*P�n���UH=3s�#6쉈���{)���/7_�$��j�������D�ZB���,ǽ]���W��_D �c�Y-��xu�.����T�@^)r���򠽌LT#�|Ϭ;+{�?�v �J蕢��x��5�G��vE�_v`qØ}���@����9<� �Y�(v�/�U��=���g��%���Ӻ4��pz��n���^3��@X��-����ɽ�z�N�f`�ag���֑7n����Ah�8%���-��p�\i�O���``�aZ��ގ���;�M��q��әu㫽�DM����j �����u��HW��#C�f=��c�s�!HѴ��."'�������G��Վ�Lہ���2�(X���z>�_�*�D�,���q4�/���n;�E��a\���[��H�$#̲+�����$�u��Zڳc��&�{�i��i�L��;��zZ{���Ζ��% ���:7�;q׹�Wc��G����8�l�ZD�{D]�~�w����K鰚3dԗ�ħ^�G9����Y�VL��e�6��ceA�#���;e̋����%���Q�}a��St���I��ݨ�h�$��;�8�2,��W�o��U�u��ߺk���<�����w7�ߟ�S��<|�ScO��X�/� ]+��v,�D��Bd�B��ً���\�UC�B1eȲUv9|MjE��:2�+
~�&����ch�r��cX�tY����h������>�ڞ45��($�

��Hwj����o��ܰ�LL��H��N���>)G�Ί���J�95(q��eF���֜�0!��-e�#H��.x`KPL�L��PE[쓩1���=�Z��V*�6�gMpXi��\�7p���xM�(4�N� ��j{�R#�����/�A[$�^6�������a㎟���|UH;ҀX�M$P����,�{����j�
�����0Y{���)L���~�چ	Y����2�vdҍLG޳l���d^6H��AI��z����IO:D	0�tT��{v�����7i(�6b�輯��
��,��]=�����%��3ꔙ��iP#	���A�S���$(J��+i��$�3��W���i���!I<��]�Ai���'�(u��:��?��b�$��z8��k���6I˾Y�nOi�Y^7�B (�rl�Nm���9B�c� �nr�zޫ�����A"ng�yj�H9nu��r�d�9#Lw��p�"yWv�'��F� �2���,��vE��oo��d�jD����� +1#�j��� F^v+�����Yt/�K�le��Kւ�����AS �8��PM!>�׆�ew��ؼz:�'����[�����3�[�c�(Zn���'��;��o����x���f����
c����ijό��C�<�$��[��l��heA1*�-�Y_�$Hd���"`�aN���O�*D���_t����7R�覆�u{�������֚O�1	���GH�qĥ��3�uO��\����6������@���M�o�+)��Kڭ����nIX����~ڢ5�'�|	��'v����̄ObAh�(�xN�<�����2���SQV��l�ix�5|t-t=~�t���?��w����u���<Po�Y;��*w%^�C_K��R0E��P��g��s�䃓�DX!=Y���`c�vMRD�-ܔ�_�`^�`�vNqY�ő}� .�zk��r.���΀Ә�w/}���3�
��F�K6������ր6�Ti��a�6�-U�J����`����=�з2�H���0Cű�~V����{'���lo(ZJB�.�#��L�Xӄ�ש�R�Ϸ��oW���G(W̏)��!뻃�N��f=sH��`_���aj��uzk�e�Om����Ue���ǟ5�v:<���fMyۅ	��O?U*\�3du2��Q �ٯ���o+�E��iQ9�L�-��'܅��N�lU˳������R|lZv`���`�ҫN����s�̓�7T N���W�)�s�{A{�X�=��P	lG�9�>�r��@( �
�9X���Ց��{�T	�#�2�@��=���sR��d�C��<�kڟ>oX��ͷ��h������8lH�b����C��rëǼ�|����+���+>�GY?�S���E�ZMz��c�y�|�a;+��d�!�y�g���MD��*�k��[���(1�'1�'�Co�U�$ږV5vk���p�>��?�!ķ�q��m�b�V