��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�#&��#�<�����-�l�dD�i�Ս���yws�tu��e��A��!Z��7'j^�,� Q	r�ջ���*]�D�<q ���m��$<�ܚnf��Xj����&#1�K��@�1�S�ϝ��J$�36�)��f�3/�%�QS�G۫"�r�R��*D1�����>(�.��7��>�K����9�ذ45���\�W����b�
�h曃�{!ܵ4xېHF��c�;%HV�I�r�z�F3Y [����Yk$t����fұ� �,:C��v���'�\�$��$"�[����ު5�+�a�]�=[8ݗͳiW[���\��~bS h�;��!��x����?���E2�!Ҵ�~\[���YF��:!s�Q�x}�&o�r$jOy�U�~�.�a;}oN����Y�I$�|BY8)-��<~��iZѤ�bj{.��O� P�l�Z�l_���ބ�Ҏ��j,	En�ԇ!�`.�ڗcQ.�੬���E-7`���Nk��
���n_;��:��>�%���"*P��XD������B��`�N�{��T`��XR}��㍉�&pc�e��_�\�ũ�4HK�6�,����9� l~�."�����4�k��@�?)��Z�g���q0��e>�CXx�SC-B��]b�u	������EE�
\A�yL*ܡa	%���y�I	7k���72Õ�9G��u�!:�y�dɂ�E&�Nw�Y��j�[��@����%���K��=ԍlRߞ3�<7���d����n}�P�j��M�ETL�����`���J�@x b���WG��a2�yz���!h�U�G���)����n4�?phG��Ŧ�YI��d�4��A>�u5;����q�E�WlK�_��ئ"ϙ�(,l!�o��J$�=�C�g�&:5Y��dC'�hu��\'RdI�Ө��N�[�D���p7H���U���%�F��[q��F��6+򔉭S<*�H���@�E����6���T'[�t�R�����V�{M#z#*����t�3���$F	۞��Ց>.�hw�2b�%'l�������V6�?���nnĢ�]K3�F��7Ȋ6H�G��bkT��x(Y����W�.}�� P�}�t��ʻ�t�K�L���.+�w���Ո�@*��@R�rR88Syt�O6�8lQ�ӋP�}V�FRв�ޙd�P�W�.1�!�a�~��o��B���X-��bRv	#����'�O��H;�wĲ��{�V�t}`��c�#���Y��!#�J���Z��y@&L���4q1�j�o	�R>k�?�W����/R����*IJ�c��F!�'�,J`�c�L�8ɱ�ҡ�ž��İ��f�D6��8։8�u�������w���������Ϧԗ�TLW�1�)���x�%�-b���'Њ0
Y�Sp{�*�@|َ�2'�@L����㰯���,>�b6Z�g2�-F�{3rU�l1u+�o�إ�@�Әm0��m�����)�'c"u�z?����s	��1�Uݩ{(RS����R"Z΁#��\�6�yGZ����3���u�?��ۖ��c��E^¾�m��Αʇ����{����*皍����<G�O���g��ѝ)�� ����k�"io2�l��c0��'�&N��E��"������s^�moja�%@A���v:�מ�u���_"4oK��E~/�50x�K���7��M�5���+M���=����A[r[{��+-*{+bt<�m�hcsYī�ƐZ�p:��?�$ Ec�z�7o�FӞM]�ۻ�����'�Lӹ�����k��J]GG��Q ������w��&�`1#�b)〈�ȭ<�IO:�dz��@��O>��� ��0�	Y.����0�~ܲc(+��a�!�4{�l���~=A㟭����i�F(�N�
��[/�>VBx
��?1����x���:�H;�_�i��2:�Ǫ�A$��-�F���B�ȗ�Z�V/��r{�%��~k98�ݭ)A��H���I�}��]�Ԕ��z1�]M�9�,ZX!��d�m7{��4OM�֙L�\����GQEq������胐�{����lY�5ό�c�uB9�x@Lk�7�樗Oj��5�jp��#Y��� S�-��m5�pbIxe�/�M�TY)��ڍ�?lӾ;4�b��}��rF/2y��@�L�Q�u�B��E�	�W7"W$(��%��`�GKZ�8���{�g%�k�q�R�7�rUD�������f�Oec�&;�QNſB	+�t����vL߼e��}���ak>�Ӿ�n-�-H�}:���آSo�x�-G1��
����m����2�������6�n���AQ�OQ-6KO��¦}���c�p"pK��"�N���"M=�~����۔ޢ\վ�^tWm���.��O��}�����S>��n�]�QI�W)�ޮ�*��Ӿ��)�zn�|���6�����Hi�X֌T��m�� �V8����l��B�U������0SqVk�ӎ�BO�����WWlc�YT�ť�j��{�
V@L�-~��x��gO�����8y6�p�~�ܠ�Wdr5���o�M-�%��ѽ��z����n�z��?F��,���xytڪ,��"'����[x+�%K���Īj�f����+�4�Vm�C��\|���Lu��$��O��؉��mʚu&��X�W��T"�]_��$o���ǽ��?G����}�2���[LR�S\Ɠ�G终b�s�ݨ�qv29gƤA�:�~���9���E)���e��?�}������r�/K����~f5`�zeJvp�B������y �+�t'���0���U`�+\F�^z?M�O�|�I�Ɗn��`�=����5���d��OƶF��R3(>��dd�Ì�w�ڊ�e#��[Oc��Hzdh ���{���H��Ka�f@N��6��VI���>?�¾,r�T6׸��A�	��UǠ�֜��(%��p�cr����f��9��X��$����kX������)�橅����Ҕ"����=S���Y����H_ C�!���-ӻ�&�Z.*�o�%ۆ��H��`չ���s?D�����'M�]�`�f->�'�X����C�It�q6w�N�`��	\d��L��u_��l#�Y�.\����o��q)�W?�75��ytJ�b�s?���o	U������ ���a�/;|T� �D��d0�i[���{V�,�ba�>�,~U�!��L�+^<*�~�e�#�I��I�W�k�%��� M�^���9���� U��bR�X�"��ð�.0�G"�;lq؊���,�LO"�@���9ا�Ɔ`�v����fc�؄��Օ0�: INR.����&��-���ۦ-��z�ߪC��!&��뭇�(yM�F5wF����v �# �B�����k�2����E���"//br~�(��`�}U+>��LBI��6f�*�M`9�0���N$���|��>@Nߢ%�
�	�^-�[��/i�-���}��W�)��$�E����/�)(]�������t��pM�ć�k�-��t��R7��,�Lk�9c�@C����ߑh��y �H>bC�V�~�
E=�ii���^.���0]�T2$�ʹH�}b�z!ܛ�Ta�CVH���i�wx�m%�B@�����Z.�V�x"�\��*�k{���RYc��Bd;�?B��;���