��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ�������������=��u8�O3G��#�}�xuI]�2�����Q��Q��������c�8� N�~|wy��z�H'6���א������>ށ� �oFr^ݩ�\�;mZ��%��q嚶	���X�ϡ*��s?���B��NL�۽7?/��|`4,��C�6��/�n)p�sȸ���i*���>�7r�{����4'"j���m���BsE-���Qe�jvbء�P�BTk�Y�|��y�@�ڼ���B���7�����Y���]TUn~���'7l.�+ȁ�����I�����"o�KYI~l�;e�BY�Zt�W���� &�0����{ 3�8�d�y��9�]�j�������9_��11�0�v�\��&*�$�3�0���L���a)Σw	 �,K������/$<l��֭���8}�����|Z�Et̃^��1{��24�g��b��Y�����{����F	������Bn��#-R��W�A�:���~mO��S�d�mKġ�!Ĭz��aA�L!y+�����t'�sM[�V�~��<���(�"�]��L�Ufs����n��Ѫ��]2ؤ͞��!��U�!��cT��ȬzI�nx����np�ۊ�������)��B�;�i��ܽH�y���f��h����vw�^��Z���9�"O���ppl�'���S'�vXf:-vs�ݬ�G�
��0��?ѷ�@��4ч�1(vLQ[�x51�R=M�W4���Pj\��2�He�䊂�
�~ޞ����RT������X�)���&V��~��/-�>�1��cI�����s�yrG��G��S-�[�x9�/iBl�?�� ��0�!��s*�E�L��4���|�}gd:�^_w�&-:�	��tFe��\
�9�#N�3��f��ZGGS���S�D�篹g� �� �Λ_CA�[���t��hƸ�Qѱ�����Vu�C�U�u�Oċ�s�vX��6�~*����;z�ff�JP0 �~g��ٷ[�Gv����`t�ɶM[���W�`^�#��N����Ͷ{�o�U��;����R��h��ƅ�{?y �Vz@%r���>��Ѱ��9� ��_�m����p���٨*�����K*Tq�6&Kz���ٺȚt/��<�֝>ig�q�?M��V�3Yu�2���\�Hؔ݉��y���pM�t!Z�cr�NO������^��VL��0��J�g	�B٫���8�����Dt7�_�>:Jkt}H���]�Eg{.�~�#�J�N-��"�KQ���½��ν�Q��]T�M��FWF�G�#˓�ּ9BٜLJ�E��5AOYy"�w�*E/{�}��`�(��b���f�Ѓ?��W!��G���=����?┛�<�Y�j%h���;���F����j�V1�{w�t��i5%#Bj��}��ڒ����h$�M|���/�j��KR�g9.�w�MN�s�'͘�*H�
�O�4��L2����BW�M�"	'ic��l�����r��C�>yQ(�S���yoB��rjЧ�-oc�("!R�>��� cz��n��b)�4o����[h}Jg����%L��H�{|�?�(��N�E��Kg��/+İ��.oT��� �nX/\R@ԷA۩��NI[=~e��� jDۚo��):uߌ�۰Z)pƤz��ûl��x�M�W�J�����巫�6�j�����ZF��+l�&τ�̷�������1JD��,"�'�,�"v��>ٰ�ځ�6�ǺDk��(饔�
�٣�MM=�&L	`��GٺE���ɡ9k�4FM�v>_z��H9`]ǎ:�	��Ŗ g���~�����v�ӂfi��4SAB��0�4�$�0�