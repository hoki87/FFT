��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ���������K5��iqn閒�XU��83�&� ���%(.�3��%nN���v�G�s����K�Ó�;H�����y{M�B���C���B���|X�wC7���_�[�҈}Ky*���-)��L��akt%��Q�1��տ;X�f`࿸���f{y
�qخ�P�^��Ak���5F͕'�(Md�z^e���A����s��b�U�v�<,,r�~�o��л���a%]Њ���e#��atR��_�(�c���H����8"�fR.�f�:�Oe{� M."���3V�֐9��-6G�7��G�TL6n�5-9Y�����\I�����4�`?�r'b�<�y����&M���=����Erߡ�Yt����_4I�~�׃ydo�:���_�}�D�7A٢v�̈́�X��[�d~��ȸ��%�ޭ�zaw8N��p����G�`��/��s����,�A�B��־75�H:c+q�$F�ŐG��~�^P�S�k�Y�K���/@�%���[b�t�8�OU����P[�ǩj�tv��ƶAEHC؎{���p�KR��^�P\�V����H"�z��S�A��D�m2a+H�N\z(�Ā��Ȝ�v�k˖�ӭ]t�B�:M8+�Z�P%�m�lZ؍����x�o�ϧ����BG-��
^� t��F�T>1H��t��'>�ޏ:��<֋"uP����-�!��׻ֹ������<D�[�S���-9)��jX>���{|�P�����Era��U���a�JEX��f�X2`E��~�-��I[|�7Jk�JU%s?�sJ��B��#�6��b�g���h�R}�(Bc�&40m|w�ק"�6��N��k�a�u��)��	���x(����c�=��¦�`)֒? �yB^��-�;�*Vc�%�Lǔg}^�;r����|�Q�v�^�|����G��Y���b���b�B�Wv���'S�r�=P�����bE��L�R o~�Tc}g���%���|�$��#*�ǋ�^�o��?�%��aҜ*IԂV��ױ�瀹�M:	I/~i�r�~��:��2J���O�g�@��ϙ"�FDs�b�D��=Q�`7��ߛ=���^t��@�z�쑹�@�Y���b2�?*���h�>�=w��jb������w%��^�;��>{s�Z<����z�7��[^�(��#*���$��h
�NС&ˍ�x�LV�x��?��}��Nv��\�UB�<P�����5Vk�ֻ�ΆEԀ�ME�Lě��8K1���k`8�4<4aR��|�O]���&W3a�W6����T^n�c���
?�}�HЁ�M�^7ǥ�\�����H�C�v68RǍ�����I@rc�N5�#��K�}ڬb�����JC�B:���6�i�i�����s{����P�[.����#T�k��xq�;8">G)�`�^__-tZ�rI�%v���zG���NQD���?Q��e��ǜJ�"�M��I���?+�q��rq��\(޼-�2�+x��Q%�	:�d��jӟ�eB��ϐf����A�h �sɬ���n�4h�X�#~Ƈ/DÈ����A
�ܦ��vt�։�����s�*5c�:ľ��F�� �e��]�{8[q�Y̦C��/��!	SO��%1�(��ҙ�R��Q	6n�OL���JR�R�p2�f~��x�L�yF�������_fj�
$�Z�'W~^������-�R!S��v�7�S�7�(O��Z�JR�1����#���>�m�J$�O��`�y��U���X�����;mz��^��{L���t��&Q�M�3�XO�ߚo�Nz&`�+a�FM���8���^�y
@Q�z0�d�7X�Ÿ����P���(�C�>�e?�g*f��ژ(ձB��E�]����>/��9����_TW�c9&�;0.�M��a�e�~��j����d�&�������D����q3J�DjY��r�����'�KԚ��^BGI'cL�:$c����qy���w8݄�<Ny�<Z�"䡌 �]QJ��=A �r<(*��(� ���WK�c�t}K!!��ti1��q*[�0�U����)�E6:_�߶#]�D`+sBW��/�E �T�Ű�PF���F��dm��ku��;خ��i�Kay?~����VK�֗%��=��KB��ă2єT3���A0�P�n:F*�_iR���i�^j��gFE4���&�3��7{����̶��4IdA�p�s��k��yP3�K�����m[d��H��[�����_R;Ug���Ϙl4N��goj:��".�j���_A�}y�o���dNĳfI����Xr����D������v�������о��e�{;�ե��$h�r�~�<�3&-���1�bEPֿE����+
����ҶgrvtVL�$���Q�[̙�>�Iy�w��3�?�pBEg�w9hT��*��u7�e{��<��T����H`�GYC��J�s�c	����(��Bda�8�}���)"��沶�o��Of]ۀ^Ik��z1 ��d�{�zw7#�qA�{r9����v�L�(X�`����&����v�, ���H�c�C]YZ���|v�rhf�ՎT'���W>�t(����86g������ a���2�6*�G�7�]ed���s2OIy{�ͦN��c<����"f���k�E�E��Te٤��~H�*])����$�6x��^dx���4 l�Wd��&N� <m�͜R�i�����s8R���|]*��u�h;kkVW��V�M���/�,Y*!b�{
x����~��ݔ�f�K�d�C�]j��6Tm�<ԃa�bk��0������ n.�>(��bKV��ЅT��Λ!��jGh�G��� �w��G�Bs��p3�����-X�D�psO�N�b��z����I�#Mg��kw)�ӄ�}��
��XQ�5�MX�w�^>=��nС�q�,5�K`�+��c�v���f�;A�l\O�4Nu%��j2Vj2\T��L�I�XZZ�6|+�|����AU�s���F���~Ek����Gt�o��7py���(�cU>let��{�q������i8��zm��������HJ�9W��N������.�?����e��k��U�?����C���P��<V
�3Ϫ���'�M�̃�H%��vfKK�����)�ҡh���rXD'��z���ZO$�y�)@)��݈�����{�E�����w�xǻޔ&�vnr5i��iAK3���X*n'ʤ�� O�3�iw��Ss��!��r��{]sѾ�����%nI��f��`�[�閉	=-tx�3L�!�it��eP�����A�x;��^�r�w�����ͥ;P�б�0WI$w{~����P������$�	��K�zG�Kb�v��Z�3бi��˹,B��H�u�
��Ƈ�>���[{A���D�q�����{u�s���-.����<� ����#�����?Qn>-�v�Δ���I�B�ݔp�2��_V����/�$)`�(V�Z_��^B��Ռg�Z���1��M9֞��>�>l�F�����<����b����]3c�VX����pr�x�05�t��5�߉���/Ǡ�N��:O5��|���u�_uƣ:�Y3�3�I��GY�Cs��(����E�������r�Q1��`$:�&I�P=Ĥ���p\	u_98jMt}i8�DA���2.���\��-�Ҡ�sGL�e[?�����y�]Ϣ{yi�e���J�0"Z���w���h�(����9fx4QPF4��꜁�g�H��±�*�� �=(8o[���r�n�F�}1I͛�X��8�b�f��XFI���9� �%��tcXH�g��(p�+���̗\�m��?��>N����@GdY=yȳ�$�V���Q�N�� r��e$[���iZ9�ո\��t�F94}E9pe\'�Y������!6Q�j��t�i�
˿|l�fK�h���r�:�г�y,T�:	U�?���Y },J�B����-&T���u���1i�<��P�/D՞����H�l\��~���JOUG�O{@A�pSm����>{���=���Z�g��?:Tn�������g�U�W���2�>��\�LB�3��D�re����dYNŋ��e���� ��#�Ӹ��{���( �BZ�;�8���V�<�6�31���Ҁ�診��gz�(V~�j���h�Ҳ8$ ?[�",MO����g8S��B;	s��Ƭ�Wd��V���#��sI�l-E눴��;�����`iU��S��RJ `�l�1u�*8��f�&�r�*g�U(y�]�)�#�WR�'�~jR�hnY|�O"����"/:=��=�A�gӡ���5$!�����Seٝw�GڦX/�J�5�� ��=dF'S��J
F�#C�l)�h�n�6�����w�?�_��7]��z�P�#q`�0��!���� �Ѝw�v'�y�cW������-8��ϥ0*��>�G{%C���=Rͺ�q�~�.h�[���sG["=��1��X]tt�* ?�6�p_-(V�{�9W2]��C�5mU��N�9Ih:٬P�Z>���w��%�M�!��y�E��Ȋ�=K�?K�j���c�2��+n���:@5~��>ŉ�����Ld��5���Jm�e�T���lˬ��9�/�V�
C$�� џl����4֊�N�A1�w̨�t�
ũ���89h��R�������R asBv1�E�]ğ���gR#��B-�d���]���su*c�pA- ���sb�Nj.��N�+����x�P/��$�]R��)�<��Q�d+Li����,�����)�������
@'�ݝih�%1߿��
�o�rw�-�"vQ�7�w��#]�VH�-�б"I��* �#I�){D9$Y�В7Lv_?c�	-&��]v�'d�x�S*����e����@d�<���tL�r��ڇ�|�2����q��3��'j۳�X�����R�_h�e����q���,�`��a, d	<�h��ߡB~RY���?��i��hvB&��B�;NsJ�>�_��ӳ�����㘰yjH��|�v3z�ú�j���Mk����  �(��1��5� O(���:�28
��fv)�����~�§���Xlc㽶�?ύ/<��Ij��>;^&e+�j�tJ_�)N�U'K�����x�R������K�i�	;k��:�@ՐF�+�ŀ�����1���Ώ9Y|4��Q�:a�����Jc�ʦ;C�<�MY�N�%\F7xެ!8Io�T��w��i�Q���0.�rյ�7��t�*��w!e�;�&����b,~�8�<A�@�;-����H�\�j�6��<�\�w�,�ⲑ�hq��{�{�"h�G���a�A�	~��G0�"�(�>#-�0�F�dJ������1`��o�NF¯`�{�f���x}�����#2���Z�jl|
�k���̓ssA�^-,DY���48`��tp�-�����t[��4m�A��Έx�,1�3W[B�>?���tYH��![�t7Ӵ�*��E����D�L7��e%�W減Q�{�k4;h)h��'(v�(�NA ��H����=w�`�	<;��+,�}���B\I(/E���k�&�|�4������K��#�6�x?�6��s��x_�YYS���,����u�IR�ԟ-M_e^��FO���
W�h�	2���t>ǅ�F�g�ϱ~�DQ}J����M�ٮi�\�B=�J�]7J�|�z���+@�/�pPm����Ր࿆�L��/�E��H���ku	�~]�������� �nwK�F F�8������I"^&J_Ӳ�����ب}�)�ǿ��#�@W[�������u����ޑ��vܑ�=h���`�:�Y�pqPa�,l�� �Gw��~���*�Bm�6�~��̧-�֪�!�{
��?LXHˀP�ھV���~�30{�4�0�W�����Y���ČY��_�>U���EfE�c'R:I�3UIn�I�S�X�bpNFOwh9�K0��D�`���ρQ������?Vj�i�U�o���|�xCO��vN���0�Q�^��"�$�4��ND۸��E�R�M\Ht�pR԰!��v���/[X.�u��/e��W��x�t�Hl�����fJaz�c�U�#x\��y�ĥw'Έ�?���{:;����HJ����}��ڴ3T�Ɨ�&M=��ZZX��R��o�v6a9o�����d���un=����C74��ӮlF|l̢3�W!�Gۍ�k(���#֕l.m�`W�/�'?��p�C!!�S����k9I���a�pk;`��r��/�j�!y��6����*09a.TO�~��T���,5�w����=�+_B��F�>p*�=*=������h\#��퉓.š�NdXh���B[$엶��C~���Y������D+��<{5�:��j��1�qBia��^'�RPk��\�%��F��P~�Vp�.�������r���f�|�ݏ�u���9��w���V߫⟴n�84!�G�P�,�0�6g��[i�M�m	%�*�-N��VD�wLǍb:�L�i��M`�	R�ɇ��0��3ʝS�mfT�;�58d���U�,�%�w^�g&ӛӑ����%�Pm0�֘@����r@�OM����"8.VA���3�A��|4 7�?��@M����R4s�1Yn�d,���S�;���({����绩�l�9�2���f�[��Hξ�,v1=)���w3M0P�&��V=�f�<'�w��bӁ��T��H(���,��!��2r���̅9-�8�K���|�%�\��n�|}9k�{��V��� k���⠳�m��d�O֎<K�ͥ9�=�-W^u|��/e�V���ܵ�2}���*��u����	��Xa�~���x��E��Q�� R1`jj��ݏZy/�}����o�	!�ҷD#M��M)0�����\����K�ٰ6ܝV���^^f�8&�9�E�r�Ѳ�� �q�p\�@�2i�LO�s*䍱�o S_�4�D#΃��OCSϖ��=�Ѿ�m.I�͇�%S�.'4'��'�9l�_�D8~�O|����_��=MP&���kX�uz5Q���Kf������"������MwBz z��-�W����RHw�� �i?��H/��B��t��x=P���0�؏��hՉ��lv�_�2H��2���?A�8m�Qm�n�U���)�e2�gJEN�������gj��c	��R��xr���b��u ����1ݨPU����ʁ��N�\�~p�=-�������y$6�٥\�>HV>�<����ꄎC|t �M���Ek�ūB��:�����,�z����;艹ӯ�U�Z��$�� z�AR�8	�>�sC���?�Ѫ���c�ڠ�OR5?���BC�nY ��K&�餟mP�}Y �r����͹��ܗN���;Y�w"ɸ�]��?��A�(���^O��^	�ct"�T&
N� �cUS�VX�Be��,*$s��l���Ŏ� ���(��
/eI�3�3�� ;Azq(Ô�X�t�Ί�I�P��̡���C����'3;�
�}�B���?�,퐶�_@&[��3=����[���0�Y���]���D]��W���ܔ�����d�8.�W���V	���C�����0r��g`�6i�����A&8�3�[i��`ʞ�yn쫪�Y�k2OnQ2����#J5�(�&L�2������Y����b�3�N��K�LI�떴\2����vHGaeV�x�#r��g7Gv9��B�m��&�%:l����L��p<�6���t�[s�� �E��4`S�<w�/�2��ͭX�ðY�Ҁ�ѭ��6u��.�8>V:
�������$4����{9p���x����-Qp�	����şz5�VZr�`��t�ή_G�b���)����5��6_�
38`M{�4�^���	�����A�Ч�g0�������F~��@���?��ÕM��-#�V1��Y�v
��T=���V���I��_�7|q�[�z2��Q m!��J0����83�����@/=�P_r]���o]��	3�4��Y��mln�A�#�����}�B�
a�֙�Oa�M
\"!94[<�oa�'��O����(�IH����D�wb����{��#'�.2����088��ig�j�Q(ܘ,�d��᳋iL��`���bAQ�s%'@�-�����"�����&8��;۬�E�c���"c �93NU�xM+�ć,y��*������:'W��x��b�B@��D}�Fd�G�,�w���f���'#]e���mԡw�?�Sm�_
<�ÃN�rA#rm+(�áԻ��1=�Z�C�(��N���ӛZ��kiu����&�����M�۳w��rt�V�RY��G�BpO4���z�ʮ��d:��lyu�)�I����(I�R�8���D�c�kM�_�rT��v��if����!� �Y��N虬A�<07*���~�v��gs����؟7��s�J�����F�％@�֍;v�`��*Gff���TTN>z�DJ>��X�����;��'�Ԕ+�O~�4��NǏ*��O�.	�№��h����F-!0�|�!�b��(�T��q�3*_��j��#�2��PM��vX�M�fɵ���e�����Ap3���_�?<��C�����?�MfG�8^
������Y��s%b�&���W�9�%1�û.�πۅMw`