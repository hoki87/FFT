��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ������������~��LF>�j2XE�\�oB�P��9�Tёy� �����b��<�AE�"G�U[f�U@FIp+D��~�C+ҕꏘL9F��-����D��?�K���T��TY@8,e�*yf�RM�Ð�;��d�|�n��7����	}�эz�3����bkRi�U��w��ȵ���]��L;2}�����0�W�_��cm[���b��v��ZF��D!K����v MՠK����MJ0�.{C�4T������/ �]{__�M؀ǟ���u�**!F��,��w�[�JUg�g�ؿs����3�Q?��x�o�� �m!�#X��'�O�%D'{ ���-{�*��آ�]e�������T�w�Y,M�=�1Q)��n��[I﮹v|	q���j�4b�,F&pi�PS-��4G0\;YOR�]������u��k9����[Y����߶���AL%����1;y��=�e!O�ct�[N���+�jTJ����r�SuV�{�j�)��MN0�ck��Ũ�������l����J�m�^�㻐��p$M�G��~E��w��,-�1�B��F�O�&ϯp˲��fY���9��%�xY�[�0�����3�t��\�ە�V?�%�	��4�.#�w�à@�^2с�.*�H%��[{[4J����gc'&��ӳ��>�hxn�s�B�
��8nB=:�wؿࡁE��fj�0�5L����U,;�s�g^;l�۸P?���2�-m�����V�⬜>��I�$�<�4�t�W0>i��R���5ñF�Z|���}�Ȍ$R؈F�X|��h��*d�W�u��(�#�g���u\E��$C5Xp��.��+d�뫊��Za#[l�a-���i�|�~��aQ�8�W�$�H�"�^L:G�	}�0���4�X��Α3��!�ս+�=&$���Z��WG�?`��s��bj�q��@�� �y�w���!p�y �@�;
=��I6F0�����qJZn��w��C���KP���.d;�W�~~kK���(6o���D�!=�r��uԊ��Z$����n�ny&�5�ޯq�~s��Z��ѿ�+5a�O8�����n,���Ǿ����6��mPA;��a�K����O����'�U!ܤ���CCB��f�������Zh�ᅛ��N�n�����-Ա��GA�;�x28x�����	�ZeQ^��O��ڑ2HVY����o n~K�g��-F{nW@탖��;�$Fg�3�&74b%�ٜ@Z���uޟ!�"CYH�TĿ�r40���w��	�1�qzj�:��f�\^qc�D�H���ߣ��R̾�s�����/�DZ�`�GKj`P���M$ޭ��S��8Ƞ�t�eUi��':B��z���w ?y�{4��t�ݵ�)���}}��D�����;=�dNT<��gf��)�K�|��Ei#��^T1�����:+�t��V1��+c��lr��iak\��p� �^BsB����L�x��u"F�v���ر�:���<d��s�SR����'����xsF�A�l�,l��4��ߜ�)o����pX�w��w���v�Gc"X �}����O�IɈ��7P'ݬr��V�׻��$��s�%����J1>�5ÙhH=h�)'P��O����up5��8�1$��ZG�:S�y��T�r��;oo�L��a���ۂ0:�T�^ʑ1<�:[���>
�ʒ�%�c=������v)�-��U�����Il��E`# n�,7�E���^-���۴�-]m�ky$i�ĥpŗ��A`��`�^g��y��]����0sid���K^G��.=�
�쯡��4m��eS4�lվ~�b|�7t:���6(�:�G��X�G�'j�?A�PHA�o)~�:c�X�y�I�m���sp��:v3���b73��Z?��wE6&"�	����j֗��$JL�T\Y]%eri
�xNu�--~: �dvN߼��N��T�8.��QCJ��[�u妖&Ҟx?�ð<Uo���*`*B�^C�4N���K�Ko���74��r��mD#�b+_>Lf�����%��	��x�*�Z-E@/0y����7��\�g����t�K#7�٘���_ܑʽFn��3��G�j�������:5v�f6�^�����^)�P�5�n������*���B��!�@u���ކ� �w��(���%��k���us8��N��Y�;K��;~ q��CLle��ڲZ�կ��ҳ��-�sK�:��5�Ռ��
*�:n[�0�Q�a mx~�)��Ү�V	�)�s�<n��r�\�+��b0+�}0h�,}j� ��I�}G�ϩ�`�"�r�}�
 nN��z�����q�-!  CH����,a�������X��p-e�w�7#��`"�B���ԅd�+橷�B�6Bo��cds�Wi�G��;;:ڹv{�B���q������@�ؾ����2|�Pos.���JN��@H01��ǌ9ϮQjp�.�	�Ҋz����/,L)�39��h,�j��y���dA�� >�%�t٩�!�G���2d�R1"͏Vn:�=�`���c`ܣ������M�5 �}�GZT�̶G����GGE�I|�L�(f��\_�H����+�b�)`Ύu����E?+c�YjSoꯂ���W��c�`(t_�A����a��F+�G�
���Z�g�8@U�	�e:	�u`��S��A�hk����4��(�������G�益C����muI?��&�3�T[hS��F�yԴ��3�y�V}
��q��s�Jʍ����0���Ŵ�]͠k�ɉ�u�����e4
ȥU��r�8�������H�s
��t��t2��z�j���!�m:���;0?��\V�g�t���'`X�y��>�7d3+OJ3X����O�:rL}H�v>��j�]>�haf�Y_~�����aC�>&1�mY*�)�W��S���^���"ˋ�(���6�4u��5�˨�C��sg��gF�R��,eOD��Q�6q���b�x���t*,Gl��֊� &�	�p҆��1�5�i�q�L[�'�kH���d��ф^+R0�9MK�T�G[eilW�6�{�_�UlJ�3/Q?�����"$X�8�ZĦqs��hMf��v����d�V����#����:��H�j���TF!�p8bm��I��5?�F�Ӑ(<cU�e�P�pG��<D�"��@�-f�T�.��U"�:� n�H�W��y=`��a� -1�ڢ�z�k�q�"�]W-( ���0��7��384��3�ۦe8��-R_�锳���R&���$���D�D��`n�&�6V����kqmbVئ�+�E��Jqrn�r2��ގX���G��ؚ�#��L�Unpa��/�ĥ�����&u�i������E�~A��a�,�N��&�p%�tWj�j������.z�����C�B�Y��,��n�P/7 �9��w�e�S���`j�[�s��j�0����]�yb�0
(���n7㓶�qp�VU���s������V��)@=�rN�J�Z^�� �1XxY�6tL�"������>�`{K/�ĥ9��[>�5i�G(*�,{��J�ΥJɴK��KL���%���+k�IC�	bS�������)1^c�C:�g+Y���v~H(.����-M5�b�?�C�	E]�㈸�[����w(+�H� ���Kt>�rlt/��p@2,b�uJ�0��	'��� ©��t8;xk�.�e�C���g)��k ��f<���$6������,������c�?mS�a��T���v�F��ԉo2���؛���+���j0�s8P�s�¼�g�8��B&�ʡHJ���BA�/,���&p����;��~wj�쵣����K��gףp�z0錇/�6(k���;au:����.�Rq����&ӆ�]�����a��
��P"yD�̓�Q�g5L�����w���~�����6��R���Jb�W��V|4�/zs�X$8�,�I!g�{ۆ$��~��D�$�﹍�N�"����U��LSy�������V;�W�> >cO'��ܿ�cף�wdq�7�Q�&�4k��q��\��V�?��R��lm������ss
�$<p�/<�ֶV���|�#�!1�"�w"4�f)C�����e�<�F8b�+Af���f_4����<�B�<0����<TS��>e C
��
�#����p�(�6�ڋ53��bw�r�
���ޞ�jg���Z���7«@�#3|��ŧ����<Z_WXh*�~<��O1�ϔ@^������|i��JԽ4-R	����R�ɗg}�|�C�yK�Y�mY~����¾MU�[���b:�+']V���誃>=a�fg�� ���U�U��܂���:�ִ\6�&#Rߘah���i���ߦ	���Q���?!'md�2�@�Y����Q�(iP!��G�ok�2������}�{&�:拠<U��LwTH���b�\����M��Mi������:D��rra2�+�B$
������h�#����ck��eF�wW>���<���XD����k5�f�[7�9c����6��%cM����c��g�8�.�u!вC͓�"��=Ѹ<��L���u9~�����R��)e����?�A��� �fn��5�5x�2i�0���ω��M�۾$ݼ���i�(�LX�M�q-�I3a0ş������>�U��00��-y��~�EKww�Oh��q8�eCI����]�eQiKkT��^Jp�DX��ML��;z>Yvk,��0�;��ZH�ưT��Et�r7X7�*:W�M_���cU��Ǿ���P>��"�$!hF s3��̓[m��d�[2u���y�za{?�N�%!�U�X]���y� q⧶��h;��ea&~�[�tH��q��7T���֮���(7����0�`����Pb��u�T;����<o�����D�������#1!�!�R>����H�� p�y#h-x��#w�,���&��g��QT��L�=��LT�e�߉�fE�J�2ƙ�J�W�ȩ���ۓo������F��A������؜��]0f]�"S�����]�����3�W�Ka���i�ߋ]��u7^|�Z��͘���4P�_��rH��' M�T+T�q�+��7VCù�I��iC좜�%�K���ŧO��k��..1��c >+��H�"��P�)���r��,��)�gG�+<�����?N[<@k��6C|���݉)'�F�Z���2�OVL������ C��+�����P~�,��<�Բ�,W�oӲ�QXX��:\����G���	[��7^�%�X��	�K)g��8 ��%\/Q���s���"J��)��Y����I��F�V0i��p�ǽJMl<�[+�൭�a����2�fF����"a��s����&Rp�z�\��������W��Gl�:��@��1�02R����ܕ&M0�`�.��*��eBQ��U2u�fD	�4S>�Pc�%4��>�F�G�;ne��.�����#L�)jL��.����W܀��0#ۈ�S�z��u+�i���+��ڛk�L��{��|��i^O��;�3�%'Q�� i�C�� �k]4���E��ڎ�ȕ��~�/�-T�96���;���wX�9��ؐAJ�^�����e�v�)�$ j�HW:"H���5�C^�e LZ�&��I �<�/�����nRo��\��7L�+�{����4a:xtw�%E}�@�7ȏ�O��?�!�y4�B��9M1��JL;7<�;�v�%<��_:65��` e^��i�z��@}$J:W{�)����NG��sH�s�IlZ�3i�����|��z��j�c��3�z���S���IO�C,��Z�:���`��1�O�̓�M�(D3�3ݎ:H$�˂b���	܅�s֎^=�q�ҨO��`{�7w��,y�����:��ue�5Js*�6,���I�6̴g��6��?�'�:o.)��j���W���j�=w�d�;v���ߏ%��*)�">��w��T5k	dw�h$XMڙ�Ǩ��mlx���4�G�~��{�tbrA��D����vH����v^�p�xN�^쑦I ֖��W���bC4�8 ��r��S]�m�� c\���$]ov��ܤ�jgqZRK�E~�Ns
�L ����u�R�a���l!G��Gd!�[����5�WM�����ި�1��,@�L��ع�&�5���mI��⚨扠t��y�3Z��WW�O%�i�1�F�'�Gf{]v�RxL&��&�a�#K����g�`Czq�D4~�`3�(��Jä�,�� �� �����M��J{��_vh��i�����M����8��o���}꫰��Z|�7P��A�vߐ�����|R~$[�*�P�'i^H+:^!(��B'�h��@��Q
D�e.d�kmۅ�ri�����j�R��=wM�.��G�v�>wR�6�����/�/#_�ǯ`�&�aJ����AՀ5,A}A[�@�}	\��;�6�\��e����l�@�dV��hvM��iQK���;!�h�B+x���xp��3Hd�''.�4x����A��-I�h�`�P�����|����cV�;<-�Ѳ�����!�L�����E`LEYOko��A�=�C�qp�Z�\��|���k�lxC1
#������ww��oq.�˺i�9%���@��$���n�9�5a�*��L�ه�O�VM�#�Sʳ3��\P�7����H�� A%y��=�;�̻(!��x��r�"��	��hF����Ԟ�|C�+6
�ɿ�6gӠ�"x�q�3�;h b��� ���8��H =7�ow�5`:?��u����j�[�ɔƚ��7u���g{�Y��]z\�}�<��rd�oU��g���e���<�.��f��oޏ ������9�S$�9��y``�����jϞ��S@��f��)�pS��J����$pF!��P��j��?� 0�@�Mu<%�ѻ e`����'���α���JV!q�H�D�u]յi���4��������C�t�Œ�V&~w��H2t���QYЖ�@����-��A�p2Z:�Ҡ��`}Ŭq�*����T�Ӛ��߉��M�?;3N+�~�K�8q���E	Ȩ��( gzyȈq�Q�[�a-Ӓ�����-@D[o�Ѭ���I���<qԄ��k�$APǩz�3�UF�pp�ʽB�4r�*��l�L]8"���*<ɽN>*k�z��E7k��#�Q������4��eQ  W���y����byQ�ww���(��Wͮ~(G�s������v���S�E�ZH�1�[����-�c�V�A>#+#�#�uȱ9յ�0P�1x̆����;YY�Y�9ZяOמ<��ح�\��]_4 ��n��B���4�|�A���O��z?�wͯ�� �ܑ6�vz�M���`��Q����a�I����r�����n,�%������n�nǒ�ȅ��	4U��jBro�8򝿶��!�y�SH+k���K�#:�j�p+=�"�G罋�s1������p:B���j�#�Qِ9c�fw4c���xԑ�E�I-A�\Q����\���8��x�T�2?2��gF�\�v*�-Ժ���R��S� \�./Io��L�]  �shg8�\g���8Z9�ek��xW�l�X`M�TΆ M�a�7ʠ�r�J4�x} w|ػ*�"�'h0j���ʡ��^nG�|�L+�4�ͽ�vo�=&^}*UT�o��H����ݦ"M=8m���e%a"��T���!�,�j��<w��R`_��ѩy!~^��B<�+8��	��}�eЪ��W�Q0�<�j*�gC$%M�B��0t������:��!�<!���;�KRV��+.�k%��4~"n �ޡ��XC���&q=���o���RF���|����/���01V����� �jS{��������9��
D��C�a(r���������>��"��>D�Og�e�UꗬNx����{/���}��$�Yn��e4�t�:��'@�*b��Ҷ�t`)�,o�4�c�GH-Z���[1��P���3���_f�߶�������B�xwH�9��1�}����1Ji�|_,
��%�9�^����c��'��Y�/X�ifu�/�t�G�Bu������ϢT�~�3C[?����cB�e�G�U�}�,�U%���h��c7�ZЛ{p��Kߣv#~�� �s�l�
��B�#�����L�_g����=k%<$�g�ֽ�����b��Q��
1��B�J7oG�����>ϲ.OƆWM���N���7ᲾP��le��1��!;�Bܡ�d�~B���׭24�p&��/�"���N�#�Kv�>a�[�������G?3s.zZ+���u�e�6O}�J�_I��o�
CK7M�vVYQ�D;�@�t	&ۍ��n��iչ�Ъ�*���ێ�\�@��m��};�͔��3��;����=�1�:|��P��1JS��{7�����K͋Ef,}=�N��[��ֱE��P�Z��;e����%��=a=K�,�Ӳ���S��@��
�7^}��Ap��´�k������vo?s�cT�h<�\�P��/�)�h����#.�_����L�ȸ���eU2�����~}Me�<��R����n]RŅpC����eUΓ�7��
ԁ0�C�Vw�P�j�����c��>�p��n��j'�1'��+�qF��r��?i�4t@6�S4�%�<w=8�ԁJ[��uv���et�]�i؃����
kI��H�����|�����tg������9sf���hȳoS�������^t������ef��n
��<y��rc��L�����U�Wq8f�����"�\|~J����9p ��eT���ӛ��<�;j^.!�K��e`��H-+�0�5��yՙ�1B.�"|Ȍ����orM���ٳ.</2��| ����1�eb�~��K�|�%������a]9]�\B��cd�Ǟ'�!1� evQ��:^�~8���?.p�aj�M�ߚ����j�`:�J�^��.@T��,�#� /+�������+12���-��N�@M�P�ɸE����QK��,NM�U�o���e�P׳�[�z 7�l��Wx~��@U:����'40��i/�!�L^_�M��0~���*C���V9e�����e���R1�8���g,*���`�3B� &�1�e@�Y�J���Tf/"9~n��z�ޕ�n'���	�!2]���|�Y�FƧ�?�I=Ya�J�U�Ƃ���Gz2�y�X�����~�x�Mp�P����0�K�fS���F&O
��i�AN�Mb���dH*�A2������tJƫi���Ad�Ƹ��2-��p����:̄��ξ�9�P>W�=���ž�!� 
.0�8�ڊ�cV��]UkJ���$s�I<�W�D�j�h���-�X�aR$����5E2�I)�3�k:U< ց��r�"S���$��gs�����3צq��nKQC�*_��pî,_h���x0�@=������^�g�?��#OoF�Zƈ�D:�s]�@��陿�0�U��59��a��0ʻx����Zűr˜�]��5���ŧS�l��ތ�� ���o�x�|=���nx�*�O'�Xnw[���1$��j��J���9t/�><�:�s�̸�������3��ߕ��턇��o���פsm{�l�X�_A*K�=P���jiLgH�]������]G�����_�ٽԠi��/��*'���?��B��Aʤ��4{b4�, t����"[�.u":�Eȩ2���9���H��T��qkܮiM8N�Ȟ�l��/9E�˺t�S�+��o�m/�q��1
|F�����\��
w2�
2��z���@�Ӵ#�f�/�������Rd�$��a@՗���FܚQ���̻�']�c�N�N�+W�Pp� ��>u�U�qT�-/��=Hm���{�%�\+�f���[iɏ�0��{H��|���$FnX�n�a��=q)�;/M>WU�D���� �T�V͵4�\��㡙Q/��L;D8C������}�N
� ���	"�Ձ���n�}��8���5c�^�|�,�7Q�e>RqE`-�S�x����}Qq���4|�Zz!}U��sd(''E�#b<��Ƹ��gt�a��� ;YWw��%����ɍ���Tɱ�S�߃���(.�(�1ZD�쭼IC����u�&�>+�������bf��%��J�Z�?>wS6	֘:��m}�_,�v�@�,�ya�?��	]Zz���X���`_�6���դ'.f�/�]ft�C�ґ��n"0����Pa�?9����8\�$9����W���7ݲ�������d��%.B#��u>4�g�����f�KA\;��=���G��T�Þ�:N�կ���d��I��s��ɢ߮����ړe��FW�Fn~a��1�6��E#_��9���
��ؤW�D?!�Ukn���4{�_ �+����(�ڔo��6ٱ([;��H�>��T�Z01���B�O�)�S\����LN.co�q���Z~N�kr�I��	�Y�haV�J�kTyg���O;o!/�\w}�E~(�i��U;�L�����5w||��f(���$�E���|����d�*�����G�ڇuu�ʉ�G7]����0!9�TR��v�WU����ۖ���%�՝�2�BV�C��!�8z�����	�h����״��6�G0d�B��7����v��[��w!s���wJj��W�#���%�h��3_�19����c΀��4<��Ӑ'ǋ�� f�KN;љ=�af��xa/a7��K-Y����V�U��qmբ��~)�"��_h-W�����HؓOb�c��M6�q�AF�{,ʻ;��L&�������q��M�W&;��������n���7�%N͜��� ��Q�\x���K����'�1��c3�Pը�ޓP�{'�ݚ�R<_��7��i̜�������~Y�yϝ�����`_>�IϩVV�;��|͎�c�;�t6�%Jb��_��)@.�t\�����u�tm�_��M]� ��7}䫠���2�?oJB�|3fl�:)���l��~�n��� �����*>#�MK�p!�a!`>s~��������]ٍ)��-~Zc�)�@bU�����$o�Tx}V�)R0z��\l۸;��mF��/GW��մ��dv����*��>�G�+G��x�8�ŷyC��w��b����0.�P9������ݭ��1]������CM���Os�0L��S.w��ߖ@M����;l$��ċI2SH�+�Շ�*����/P��qu?*�zD�n��X=��VO �*���Z�R�g3^���]����8�v��W0h�(I���k!��t�Ċi[�F��|b� ��CWc̡B���	X�! b>���0W��Zdp��M`F�0�����֢���miP���m��Q-g.����%�/��0�� ��4�U�!r�K
��hW9�M�}�Z�͝�u�m��6ޑ�1���M���9�-��!�n<�Y~U.�$��#?��:z��O����XJ����m=�%�!>������=���o��q1h,F@���"	x��� �Pkaf2=�m^m�Gۊ�|�`J��(v�.](�|��I�'K(�5�"�,ه�U �!�k1�n��r�����Z���sRђ�ַ?H��H�q0�J-����"������$�64��kMa���Sl��Ӗ3n�*����9D�;P��L$��+z�2ZJ�?�eS!���	�?���� 0��6����) �&K*�Ƅ�!f��Uf�q�T�0�����R��,�q��MǶ1[��b����Z��^w�.�^���N�U���;)��ͮP�3y�����J��x4��K� ��3~2H�<H{�f��]I"Őt���L���#�X㍿�Β��z��v�U$��}�ҳ�A��=�
�����k�u�pi�R+n�(�S��vA�i�X.�|4B2�|��Pb������C+�K�8wa��D���e�Ig�R��>�T�5�_3���'������H����o����5�I޸�����]�SL��=�Z�%�t0�f�rhj_�S=�N5d,�<y�vX���I!#'�%��Xg9>�Ӱ��p�}� �7[2��vxs�`��H�k,�����P��)f>�����CZ��?�=�d�\��bo��/Cl��"җ��h������ا��!@�bk%m%b�rs��3���~��_������p&y����#)�h�K��:�W��a�l�qv�n+��<��ZU4w�3�<�&0�b� O8_ф}�9���"�̸c�\��}�K��%�AT���a�2d0���d����O%��ƫ�F���
��I�ôؙ�zY�d�D�fp# d����S˪��88��&}�A�Y>L��>���;�\/t�aո8�.�x�-n��Xˆ�w��t�_e>��c[��2�l�`�Ԝ�*���ۻ�}n^&-��vR�����f����FB4��M���]\��J*{�M�ק!��<gC˕���a��m��fK%���)��I:�R�G�;N'7�,H1أ�E0 ���@�}?WH_{}�[z`�b<�������%��h ]rʽc7��'���n�MT��t�9Y/^!@w��g��fF�ij?ƌ����-&H��U4��<{	�����Ĕ�خw;Y^�3%��5w5�+�ʠ�T��N�	x�#B Kf�K�v���!Uqlt�E�V<�*ۥ4���� �m9B�G���#sKP���Ҡ����]��cN��+5�&GF��&wG̒�r��8���&��+�Ll� �*��s�i\�I�P2�:fJK�H�>�1*��>�����{F��''dV����.��/:�=�͊��V�\��LwhX��X?K\�j}���N���h�t��B���4�ʥ���aq��<��X2��7�O����_R� �I:�>�}�BV�� K/��W_�yaX����TDk�0�_�Ce{�O�r��(v�]�o��H (D?�s�_�w��Xd��S�b������r�I�R�Z�=%2��E�we&�Kd%��x6�,������d=��_�t��А;3gTV@|�NBx.U��
3U�̉�>������=���	_�Z2�fz��ܜ.ٯ��_��bs��6Jn�{��'��UE(t�"���e���TOs�=^r��4-�ؾ7<+Nu;,V����D�Gb )S�4��v�`ațZ�i��dUc
΋��%Z������KN��-v��ތ�X�g[�1ǧ��w�`�L�pW�N�-���tn��FϬm�H(s0Z��9
X	���ҫ4 6R��vK@'�R��r%�c/��]F�L`6���e��|��A�@�d)�F��:l|U/J!0�C��ף:���ǆV�_4��|�;s-�t'���:vX;媱�VSq[��:f��0K���\�b�x�*"Z3� �$�1�yg'o� �ʼ5N�Z�A��JΕ�&b����s>�]6���,�,�+��~)����Sa]�����XOpV�5�J�&M�Ƈdz����P���p[�d���o�b#�{��"�c�ZVP�D%�>:X�Rz�s�ʮ�4�r��4�C�{��<'�0$�/�f�/퉻E�+'Y��<�	\�w��"��2ǜ8d�8k��o�hsn~
Yc��/!�JY�Ė'y.���̳�>��f	��hp�3l�n_톴v#ĖB��~�w�#m�Z�,�vNW�ȭ�U����c�uR�����*<S-��0PX����bZ�֞��0���-�?�[��4Ru��B�:9
�[��&�n�n�i��܂��h��\k2���`F%J;�I5�.9��L�'��{��:�%9�%�Ųv��� Y�h���� |�Ó]g@U�mMsO������i���k�,i&�1x6����L�P�f�f^�މ�h �����*����7+X����]W'�����"N�`GO���;�F��[X�PvK����u��Oh �����d�՛/��F#K,%u�@x��O-Qk�ǿ�Ji0>B���m�7�*j��f BD%IBV�7Ț9G4C�<�R��n'���t���I�qP��1&���@|��*T�۽r!�� 9S,T2���v]Ɔ�kN=�0����h�a{DY8�_�e�������6]���:1b��ɘykGU�7ؤ�w�ϋ�'�b�������N�D���m���|�M����� �ڡ��P�~�!sB�y�k�@Jx��c��"<�gw˃�^��Q���`^+�*B�i���׌�MNǞ��@i}B�0�-���G��0�6rQ���B�М��ȠX-�E��f.��O���vf+�	�_/Y:ο	�$wlmQ���"xD���oB&�eA6a5�C�$Q�s������x(�ˏ�h-�A5��<hEa+���uL`ĳ�d���%��f��,QW����m���$|9�B����3�~�	��D���TwS�%��X�$$,����/�Wj�lpc�I�ň��TŞJR�P�e}�ͷ�_�&4gu��Mx+�d�����A����m{�5���~�4���;�eSGx#�"_6�L�i	d�*H$���.�\]������ (�f�������3���Tȗe~$�	JpG@�W���2�_�ֿ��os{Ib����
���dU��͠�S�C�L99ͷ�P��N(,B^�c��, ��oSO7HͱU.]�&��?�ѡe��͞DG��朻��3�������m��DBE��|�Q��2��5���Bo�U�r��TcB�D�d0y�v�!�'�0�4F���e��,���-*MLR!	Y
e�9��ч��n (ֆ��M��u	,\=q4�ʆ�]B�O*���'%*�^g}�����C���D�8����#"���mQ�	ބ�_-^�nW���@��nU��,���x� ��ݓ�m@d>l�0PJ�=�4m�K�<��f�/�HDMA�!�U�
�J&�Xl��*~/E�u���a���<E��+�7�W��`)���$�v5��2-�6�%~�����P�:��p���qu@���HA/%�����K�X�q���H٠	�xo]>��S�8{��0�@|�y�jH�Ģ|�Kv�vQ�c��߮�6�g	�L@���{K��ь2ދW�ɹ�����wg"fKZ֢��PO�����J�&c�!��]������D&�+��8��2V?Y�Ό�Ԧ+��35�I��p��r,?�T�~}��/1���ZHm4�x� ��.�s���O$6��=I�WY�Wn�MY�� ���h���$��oi��x'���F�)�h=���S���r�����o�=S��	�9|X� ck���j(+x�IA-,]�+8�͠>�D�=<^�	S$vlNQ����t}�3�@��"hW�B>��z�o�����X����!�[��>�_Lh�G�&���4M�`�ĺ�(�x�r�Ҟ��ͳ#'�-��[�q5�Eщ��E �T�%V�A{-æ������4�3�3n��t�,���g�)�u��7m7��2�g����~v�]�|S��]	�*�&��[�5��̝ݎYWJ��4+ݹ�[݈pc��(L�&>O-�VB)��4a�����̔8|U�=9�/%����Nѐ�L� �dݙ��0SM�[_����=��Ĵ�m�[%��<�2Y♂������P%v������/�'9��b^��������@7�����и@KNf�_�Ȧ$��"/��P5��*�҇ަh·���mK�H�F���v�=�a<6�.�f�P�����8N�����N��a�W!���5�3,�C~<Sp��~� -dG��]��B4��&�V(��ֻbpof�k�B⟿C᥯Ul�㺯���I��x���!��OE�T�1�S�gp�Ɔ���,&�Q��|������(d˗��ae��3"&.0�r*k']�L���� t ��&�ς`$�Aa��{*�-��"F���K,�3B+��� ��3^�p�#�J&A�0HK��[��9g���3N�6ޠv����L�+� �!�A洺=��$l98�U��	����Z
̻x�)�~�/�ԅ�鰏�x.��!��;�)�ڥ�c�:5�T�g��^��t.�1����F3�3�Z��^B1/�B86�ɂ֭�]��G��A1��
�Qp?/9ϗ	t����`��l�\m� n��^�{- �6��i�;�/zL���u(���A״Ct��1%|	���SñN^��ke}�e��٠;��uxp��G�����:���6~���0�@6T������c�K&M3/�� �9G|�x{��ь�X����y�/��Mۇ�T�T��<B�葪ܮ 8���c�e��dfΗs0���i(�R�^08�NI'�ÉG`�`�n��q�[oO�Y��	Q�ijKC˟Sr��~���|�ة�2�#����C����M��S?�`�AClYF�1|����c��j��A�����ւ�����\�+zN=��u!��x��V��|-r-|@���՛f��94��Z}
�!�x��v5C�Ź��>�=>�BS.�����(iGe��q}h����\��g}�Vn*䱱͙�B��(�
8���D]@I�A�!c �Cn��@ �,	q��M{�q�%�l*?E�C�am���Cˊ�&w��(��%��O��Ԡ�ex�C�$5&�О#���J�'H�da�Ex��o��Fa5�2���40�I� �B �u��K';������ޯr;}�SⱭ$f�����.Q&$�V�[�J��pԷ_H�*��8�M�5���80-.
��>�z��t	�Ɵ�:58	�OR�S#ttk�QwH)��Y,�5�NSn�� ��g-j�R�eٽ$�7���Y�g��k�	b?��:?*l7��1���- �\C�m^��U�7��=6����b��E"T�;ꕹ�9q��cp�9��*�)a�|Ɯ�� ʦ�Ùa���*�tC����ӻJae���u�=�zO9fqK�����p�:<��7�`��o��B2ïj���؃*_�#���5GMS�ے�䉊m���.&�0��͒��ҭ��q}�4g�YX�ؙQH(��1A�ɇ��>v�5���Q;mw�9^��65��8��qNf���Ԭ�ȒL_!l�"�A>1mǇ�x���G!75�Z��({����J���u�1Q�`PLLsE��ڥ�w�A(2|~n�#��H~�{��H�:%���Qـ���Y.��@o֨l1���JTh�5����=�d�`��pΫT)������R0z`k	P�DB�_��7��џ��[��Ƅ���$�aL#qc��N8��ZÇ�9w�q1y��Y0�N6A��S��]�����184+� N@�ޔ�¾����X��a�"��N���Mȴ��юj-�;k&�)I
��}����,YJ{�����J"�IT�������Y6����0У��RX�I-�!,N����o�w�Xm=�#��$�j=a+wk'��܅Э�c1J|��|N���Ж0Nb�5$qD��j�����D��x���M%�$&��H%�+�j������#'��FN��33�Q�E��U�B�M�$�}�lAM2�,_ `框|1,�~�_�Z�{z�W&ũ
XM�4P�� |7gY�idQ����Yf&�z05�F�!w�~Eƚ</Q���0�ؽ���Zv������mw�ؽ#�]���݂��%jw�hm����ʘ���o0�������X���� �8$�P�?b�]00�{�y���nء[)���R��򀐔'�sw�����
��>��yV��ɑB9���[9�_:�~Bq.u��$&��Q���^�ZQ�q��O���3.���b�����xBRo_z6v*C�f �<��F1an�6��X�Wz�^޴��_.��)h�U�f��m}nc3饾4ЈO���߰:	�@� �<=յv�&��E��x�3��a�D�,��MS=�-��A&�z<��Oʅ�v�;e��ǰ���P(E�I�ǹ��b%��XU?Rx�Fw������W�S��='��/�!"��r/Ed�+_P\�_
