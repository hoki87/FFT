��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ��������� ���n�0�ּ��d{�gS.�I�[�/�d�i��X��%�,v�H�lv�M�+㮵�ӹ�aB�3���&� �Ѯ��@����f�B�xd�}�s�������t��,�d���Az2��$Q�op��r������5� �9F^4Xeq��+������q�7�`��녡0N��j��������=⿼l��@���{u���Q=L���}�,X7ɜ�F������8�ݨ�lK�z��A)�
��$Y.�V��h�m��-��"/�ֆ�����pӇ�,�_��������vu!�� ��0)���(��)=/�X~���9�5�������L���Z�]��8�cU#X��K�|�=�5�-�P*v%����~,���T����-�ڵg����T���uG�C�r�E=���4�C�x�bގ��]�f���#o��T� ���:Nd[a�㷎~�%�������0N.�x)�~VR_�x㷻�fmظ��FCI�����N~�\5 i<�-�ly�]Ż�趫8 ���� T#���ƚ��`~�W|�Ft���z8��H��4�0��F��jO1
��\�t�.Gy��sRG�L�;%�u\���F�zy{z���c��_�)���%�ϭO�q��@q;I�|0��X���"��^�Ff����z��E��mY�L�=��>y�K]�I�d��Rt)��fͷPgBn�c��I
oك��J�t N�����C�d��H��No���*s�{4�߻/H���UY�o�N�L~�P�ޖ�I�`�������p��ixt_a�"��b�l+x����r� �_(�Rܚ��U��͟5���߿+�(b�v�-ڌ�Ͷ���8`G�)��CO8a�bxV�O��o5(��`�?��i��/��ogϜ���=�-�6O��P]yFs��E�U������1e�5m��6bTUL���x�;MpO�|F�����,b��s]�pG�Pp
�p�?������V$������V�X����̮I��ٍ��v��\���(�M_�?�r�����
��AT@ �?rO��͈rt>��FNٖ]mD�)�iU�5�<>�R��[���@�����6_�I=]�/n�>�����x�o�{��u�S����O�`��JH	�=���[V��N@��x+˭wI�[�E���ig/1�#�����~���oɊ�z�&�����3�1O|u({v@�R��S�C@�:��SJ�%=<��.����f�:��k��X4,`>YI5�&���fnE��;��L�E�71���gv��#!�B�S�y��ɟ�σˉ���m�
�Т�,��TD��j�0���=��4n��U�d|Ž�6�㛛�t@�uJBe�S�WF�$����o��%M'r��^~ �hXY0=Fwa�-��ڳ[,5�h5.�pYԤ��M5�c���y4K�ep7�;0޻MВc~�v��>Vձ������A�&J?*Y[��ڜ�M�!f�eP�[�w�����N
�����
�P�1&�Vh�#�k� >�Ɓ,Q<,E`6P���Fә��Um��R������j���>؀�@^�F�cB2�~� ���4���!*Z�R�%?��D��'[x�}c�^������6��mК�}-}y�Y�x��nVc�[�v�4��o{Í�u���#~�hk��Mj���q=P�F��*�O<lc)a��y��J��<R�̋$�����P��2܀3Dy:�~h%Pe�T�L�~4�*�V�@X�.d���t!���J�Z���]9���N��g�ҍ�Ũ�S�6s���Σ���4s���LW
�l]��gg!�5|?���h����К�#vҟ܎��p����n�W�u�[�7�C�xS9:UR�u���0�i�gE��J��p��gd��C%��&�؇�YV��5�b;O�V֯[�'�dM�p���s{�����D}�����y %����毵{���>�;/���Ca����	�<�"ݩ@�EM|%��Z^�!����э��;��yTm��ٓ����������xe�"���y͐��=iD�iչ�ٰ�tX㌤0�[�	^`a�c��F�]�QST�U�u�������"y���}��,R3=)���9�ߏZ��ܴ[6M>7�I��V.d�=�0�n��*k'��,��Π��3��|��� LJ'yʐ9��^��y����P�Ɗ�ɿ�Lʞ�Ձe���(+!ɷ "
f���4��$���.ˏ�w�Dng��"!�2�e�t�(*��i+�q���Hi���H�ǘbd��>KA�i�a�yX彊�����@�]�Pٖ�6�:��:�q���{Xq��[Qut��[r�H�④0��X�A��#������|�-��-�S͘>J��+,��/�H�QT�=�r���GQ� #���� /�h��5�e2�(��:�or��-TqP���[v��!`��:��3J��
��!S��3����	�B��Y5%��H��4�E��%ww�p��w�bc��M�d�-��`&e7a�ԡ_�=����bY,�ֻ���d�2qk�yn�ͦP(���cӎTf��m w��V-����#�9��&JA�J�)DY�-�+�T8cf��g}���c�e��p��I;V�{`kh?Vqs����L�y�5�鋲G�۫��_��ٮ��MU�G���o�ir>�������[P2�ӛ�5̮O ��	�ॾ����@o���)s��Z�hH}�� �da����]��!8Q���3��(9z���g�u�D�w����o�ѡ�ID6������W��	�^>��y[�_i���o�[P�oW�F����J��jHV��]�IN���MY̴���f��
��������d�b0��5���������]J��Û�t%���hnAbPZӬ�f��.!�»L�#��z�X-It'b@A_qrC�2|�֜��P
���������yt�� ?5+�k%4�<��p�q�p�;��_�3ȇ5������j�jV�ݓ�@�8��)��b�pG��h����4+.�>P�����V8d���'��u�A<���8G�">�qN���۪��9��HÆxd�U����(�߯�(I�x�4���^<�̫�K�s*
�Y�2�b��<���T��<��2�ϒ��U��-�^z��
L�L��Um!��I	�8�7�:�}�j�gQ�)��GђK�
4)�� �� ~E�d�)�+��w�v�������!�2�!O6.�K�_�N����ʦ� �,��yʒ�0�EV�]IA1��ڢE��LBl!�k�Ϯ*�cxfԄ�<��[����̳��n�?�c�����nT(�Y�Wv�l@�oG(d�x��>�L�Ouk
c�����J&n����.O�z3k��D r����mÑQ� osc<�,5�ε�N�]�e�z��*��ˏ�yF˯�����B�Pe3	���s#l���di��Rs!�Ƿ8��~le�h�$��9{��°�E�F�4�13�#�iA��+^����{%�,c�O>5��w�fظ�ݏ��A?������M�@I�������|{��c0J3��R.��R�ze����.���x&���1i�7c쇡6KW��S�eĖd�b����	lB�[��纩KNVk�#��"VdaKBQ./F�5%�+�
NF��w$ׂ����m�#�!�M	�ik^�~�$�%2y��=	�$�Y}���U�?E�Yv?W"��t}�֟�G��8��y
t7 k��,�@J ���l���<Uwy23��������8]]��Q�2��Nq�A��*�d�!��ڌ!g#<4�����I�u��S#�<}W�݉�KS߻XBÓiNs�N����XP,U�Od}"�k�!C^� -�v[����i
RE�V�`�<���Y�flԶr��0�8,�+��ƾ�Ll�ls�����~���U�ok�j���@��.SA��0L7$�f��%�F1Xʘ� �\8X��V6嬵���:��'f�Oݹ��J���"f�=��}ڭ���(4��b��2֮�L���0S��Q�*v7�}���Ŕ7��J	�齌�e�l|���x��H椣��;uW}[�u��ۈ��_a9+q�^���m&FN<��Q��K~ L���B�]�Z����^21��2�%��V�X�+�^|�o!V� [8/�T��%�hL�d��-��P{���61�����Q��s����Q����ZZ��[�Z{�0R&@};��L������J����w۸)euV&%���>�p1Щ�m���:!�N]m80c\Oi��w*���P
j��=�u��\3S��<Zܼ[B�ѷ�A��*҅��1-|\��4i��U�[�2m��ʞ'������┾g�B2�`U>&U��]u��Bj]}UЏl/��Y���bE!�_2��Y���*@��҄���3~@����W,���&��("��}��~���{{����Yck��i��3��q��\w[��@q�&\^���Q�>1�!���2�K��D�UA����O�	a�Q�U�^��(oT4 �^>���*��a��O�J�E5�W$�?� g�t����9�ܫ+(�\�hk�-�u_[��U*f�:�2�8�i�%�=��fMUQ,а�1���?���<��\@l?`�K�Cr����9��Oġ���w~�RP-�S�_7��v���5���s[��tgǯ��}�̺��;� ~�;UgY�> en¢�ˏ�@�̏�$�!͘yY���m\� H�ZM�9�ԖR�7�CUR��>���d3�-����d�n���.s|WƂ�Gx y�$%�y n�X�kݡ	]�?�}�0��Y��	�"#�J�g{�1�t	qG�	4��r���NͣE����N7F�wEB��y�|���$ݠC�,4�����׏P������l�'�o�nV��<4�C�rR�"$����A��v��(��^$D�x���v���z"�E���PX��VK��kT8V���<�T[�@����l�;Fk��o��4ާ��WI6Xy1��\��@
,��{���]�/�{Bּ3rs?�;���6�BXJ��p��1�{2�gT��.7��!��9�G��~��@��V�a��Gᯢ��HU�}��`J]�l2����3����'��!�o���� "k�䙲�c� �Pi�N�K��j�Y�X�Y�Ze�-Ñc��zR�;�L�њ٨��7��N�Y�s~Jܡx�2���Yf���ť�W�6���vn�42ߠ�<[:����Вe�Ȇ�J�q ���-x2�̧uJ�	]>�N;s���r<4�O
?�6h�`����D�N�7<�cjZB�9��	�פ-���>]���x{n}jQ���'�s'~ۆ�;P�CNa)m:���\��u�Z%�\qN�D�)8$ӊ�HU��dQj�t���a�Y���
"g0�7]�R'��{w�$�KW�S�|7U�|��Bp���'�`�/�����=�͔�7�������ƣ/t���T/t�fluiߣ	���BI�(Z�X�*ֹv�	Y�5'K�T(�������UܒW�8 p5�1������/k
���]�d���-c<j9�1�Ab�Xɉ�j���Zi�@���+��&p�����L@�i�Q������]ô!�"�F�յ�T����8��QY~
kp%�0��Y䋸�V�UJ���v4`�7`�*�a�R�g��Q�_i��Y�����JY���"���kH*���Ҙ��[Fr�y����4:����A8��0&>�4C�D1��L5G����d��D�v�e'"�"���a�)杍���v����wd�:�9�K�*�("����� �=k�|�JT�٥8 b��I�:{i�����4Wɡ�'�� ��:��G~�qv�2�f��=f�01M�Sd8�9D���O�۬�&[3|p#zg/μɐ�F���B� Q3����g��
���>{g��Mͻ͉��x�������O&7�z�~���^G���B��̳���D�O�cW�)9��,[�M�O�����m��b0��Ks�>�i�k.��K�v`gvܪzi�?c��(߂����m�x)�z~J6j۰P9"�˛uЗ�ݐ��t�;4�q��!qC��)Fl�ţ�C�Z F �~ti�����Ď
oC>�27�TT��.��i�/������0f$ކ�2~e����_�)�"�'Ƿ`�]Z��t3��ͫ����;7+k����=�-�ix/��eg�S�fc	9m��lm�<\�j�<��$��fO�̣����٤�q��c�T������v�C���<M�v�c�L�P�����e�`4$�Vr����xB�D#�=�>��*ڣmc&��f|�aF3o�ŉjPCˇf{��T^(R]�;qx������Kڅ��F[*J�� ���Pb�>I�a���my���ܵa�2������z�?)i�ܸ��>$a�4�{4Ɓ"а�{A�٬�#��֢�&���mλ7G���OW.hС���a.gj��VUA�(�����<�B
[��C�6+�ۆh>��גd��!M�;�+A;$눊�+`�d�.���9gv�ol�b-�5)���T�p��hV�z߆��n��rʔ�`�3�C�y���P1�E��'S��-Ye�(���*���릈�!��J;�@�Q�7�z�%�;`c����6K�:hF{��X�ES����q)��;��zƏ^G���Ǒ'}x4�*����;WA�AM�(7���"^!	���G[���:0�@�5�:�Z����X/��*_�h$T�)D9�o2�a�ǧ��!��B
��%�ӑ-�(�	�@>t���0��Z?jv�b��!�?��l���/P�9� �á��|&�Т�A,֪�b(�wZ�a&���>U�T��ގw�4W!�Y"\갞S��\杘�5ͥ������@. օE6��M3���t2��>=#6�*�yM�e��	ִA��|�A�"��ݧ{
ٹы��E��Jn��� MP���C�d�,��M?��^. +�A�����Waհ��K,����vݒ��}�Q��C�sx�ۄQ������˳9Z��_�+���?��ȮzĝԵ�����	!�7�tNM	���F�������N��%éJ6�;���մ��� Y���ʬ�<��{1���}I"+�R�v��X�κ�Y�i�*��w4�3_;�7�Vґk��
��a�E����)����>�Q(�*
�� ����O�qf�dk�?���JE�W��˔�?�N�Ez�a�ߑ�y%��ϴ��� ���h0i�DSqz0�a�X�gꍃ�l/G�/���2�J�s��lQ�j8� W�qz���ړ?��!n�(!���Q�i�C	J�;޵gY6\���mw�C㒨�x�@�*��:��HW���A�SΊ����gu2D&y�c��zO��p{Lt�y��Î볏���2| ;���rE���|I��^b?l�<��'�*��e�ځ;�;��V���A8��^_�h1u��s� ����e��da��PȉV(�(n@��X�fe��6D������VcS[3�G���2������i��A�	\P4A�u��.�I�����yL����s�-t�34�Y�w�q|�/���a�3 yF����5�o��M�/���%QB�C���g�^�z��h��L���F��w�7�ծC���r����obΩ�)BJz�8U�0�~5])��A��Jy~���"��l�(�Ht��8��Gi�� �9�-4�����nm����K1���LT+�}��}4ə(����9��
�C����Vy����~% ��G�t���;��;j����q{
e��d��F��u��%��_nr>7&�i�-rl�DvQ�6��@T~���1�8o�C�}����f�,��{2vJ;c=��2�VO(�@�Gݐ� �wp�,�(�f����:�'P}N#����U����
��/}^EK�+T�V�4�Aؒ8iɜ8R4�K�9�	V��Ǣ��l����1x�fd��-bT��G�VQ	2�G��F�> аV�i�Yh)��MV|.e���ے�B,ޔ�M��X��	����+$��7�h��:�<��V&��5�auǳ��f1����9����1������'{��w�2> m��>LvL6�i���u���ɿ�F�M�8����
zn8��k$2���@l�0��<?C,��z�4�JOmSb��	 �f;)�=�i�����:�t�"��x����5hT��1Z�X����>�[����~s�&?͈�/�%�����Yҫj��ڹ���&x�i�N�9r�����a�ԐBp.������n�8���Ew=����(���71^�F����6*���QRΠ�;Y6ǟ�TǾ���z�ξ�����tl�4K-:�����I�f|���=]ԝJ"���b!�fCD<��XV_��i�UB*�T�$s���@ph���	+�%&�c���Ζ���X��!��0�:k�@���!cSFA��{�)d��0򗻨��ME�;��*���@����)�r��>�75��ڭt�>�4�i+�"o/�m�;�v�c�_'�e� �r�:T޹��hkC�����3���%��1ѥ2��>��Q�4r}8#	ut٘�R<�y�N;��������C��}�|	K�r�1������(]���Ĳ�^��Drљ������L���֤�Vr4�׼[)lF������~�t�V|;�v'F�9O�-�dc���":�ui��ٍ���l٧���5F@�g\�?G�ߘ�)��+���?I��H�I����f�f�+5��("3+�w����lX��U�<(MwA2��i�W��SE:z��}��.e<�V�>�
Z�/Υ�O٧'L��W���RF�$�A�X%"�2�Y�V��?�N�g����`.�G�qЀ֏f�P�;��a\��[#
�|���b���:Y��n'>��5�'�F��I+�h��b��_��అJ��Q�m	�OR�U�7׭k_xKa��-n	�a$��_��^n��h�}�Rf��.,B@��E�&\V���O�R�ӷ9���O�+�R����3W[;��ǦW{Z��l;��������0s�57c�����h�m�}'�`�ћ:\m��v8	�-BD]�5������P��)}W{ȓ&���K�5�J%`���.y#�����G?/���A!�;��IX���q`�o^�3 �&{M�uba�iUI �-��#&�Y�A�|:q}��|p�Zfs�0@V�G�X��?��W1A�i�a�H�Γ\&���-��iL�G�ދ��n:���y�h�b]�RR�A�c$F�1����}o�7��sn�8����ù�����p���/5������^U*t�Sks���!(����O�m)l�(�
Z8�!<�"T�J7"����fFx�&�}FN�;��G�t��`ߊ`P�V�ߡ_�w�f��
�0TcW>c��8雎KWS0�vh�K' ��������xI*���ᵊJ�
^$Z|/59� ���`�����ۓ���][73-��Y �:xW��#hu,[��$�\q���"�?�@ށ��rH:ٯ�h>�<+�=����aҮ�ꝱ����R��p��<���U3 j�����P��o~��c
��]
���w�p:��ٙ��A����<����r��#R���}��B�z$��-���P�do�I�Ғ��c����s�G�פ���z���2�y���:H�Sr���B�����L�m�g������h��`^�j��{�M0�����] �i�x ��vy�L�}��R�x�I��
��.���@���$u���4wq��xu��&X�1�� �_d�!�y�-9u��ۛA���}5u��u�_�-/h�g&��E��=��osW\� ���} ��FI��D��>�#wT��s����v����L<t�Cq5�N5�l^N^�<��G��q�����c���~%e|H̽�@�_�V���V�럙�D�_��T[l�l̗H��HG6�O���ʦ�5��xQ�%֤����}\�{��(09$@��mI/���`��i�{��J-��J&),��c�8s�~��3h�ZR+�3�2�RM��{7��5��7��x-+9ȺG�֝�\%3�MZ�r1� �'_�!��(e��]�T�T�B�S���Z�M��47�Dh�)�^�w@T�lKjʋ��=j�n�T������qZg���O�d��[!�ҍx:*q���1�	�)���d�ل܍� Ѧ�����D
����A�O{,Ԣ�e��ø_-y �!DN�R�������@�Ʊ�Z�Lv#]<�2q�]���"�Ymf��	tR�#��7�ȩ�^z���l��NJ�+��1�e�����wgq��
�<�h^�m�Y���..i�q�t�����|���K�Ц���fН��C-���*�&Ϧ�;��$���ϥUF��?ϊX�'�@��V�����'�׽��a!F�@<���v���K������W燺���\�4����~���cοw<��T�ۋ�\� ����RH?(�!��:�YHf"F>�L֎�r��C��9`�HT
z�vf;|k6�����Y���1�(�yx#�d�jQ����E��4�[��s
�m8U=D��̓,�����І�N% i�dB/�$a��_��x�-{�5�3Wwdv�s��ܫ,�5��,�Z6����e�*�y5����dS�[pG�G�	��b����A��n//y����1�'V}ɡ���WIjyƖ:�ė����Q n&�|vL�R�v�$�Ǵ?�b�+���������B1)Z������C��f*7gݱw���-ے�^x�� ���M�5�'�n�,����-c�FA�2�U�Ě?�qe����	���I���Y��+q[�t��E#�t�+d3冗�>�:����6Y�Q �~#���f�K6=�&=R^�����Θ�Bd3j�/`�0-���"TUJ��ٻ޴��J<�m|d|/�����df�ӆ)橄���e˙�t@l�������@�y��p�t��f��4K!��׫��Y14*m~(A�켗 -]$��5H�?)����������gO$���&����ۈ�~\�����}�m<����[OA�HlM�q/!	��[/@cuG���`B�(4��Qq�г;r��o~mՅ���r���Z��k��&�Tb[F�^c;M����h��uM��岉@�C���
D��宋U�.:��.}�ă�>yl%���]ѳſ����7�љ�x̐���p��XpaD4�����|G�؉��?��,R�\��qG	�i����&�v<�K��VAnA��?\�Q����ǖ��u�e������$����,�X��/?"����}��t�(ܨ����CW"���#�^��=ت�/�4��ڷ���ԋ�Mt���	/Vq� �~\�SR��kZz���I�U{�Y���Ô}:���ث��Fl�ͼ��Â\>^f�.�(�(G��ɰ	J���76��Dd��n�����������k4vt|����l���m<[&�H\��O�؁��Z�V{����!����Zn������O����m2wuO;~=� �n��v/�a�Og%�{�z�f���PA���(#I�;Yl-�_D��F����HGI
<�5|����������9Zص��<_,T>�R"�d(�s�A��~^��j=�BM��r�숹��U�.�Upu-����-�vqs���X�<y�dy�g��iEؘ'��D���`�F ��`��D� ĐM[�X5��,xD�����4��~����C\\�(ݞ����֮��%����1����;���95�Q�8�-���;-�����C=���#JK'�%�����#ݫ��;$�O���F�4��f��A�E*����s$�<>C��������7�]�\Ϸ~�{�ϑ~��"M D؞<%����m�Rgba�G����"�Q��N�������q�?Y��_��Y�[�$���MC5�b�J�3��KR)�:�i�)��G �#U����x�m�hYk�\)tK���p���=�&��3��ϓG����EI i�"B��.oٰ�$W�{���?y�v��԰����0�o
��V�g����N��J*U���혤e�7Lhb�B� ,��c�:�w;�^��Dw��'���iBvDҾ���ə��H���'&��A��К�]E������ �8<�7�����٥Sၻ;5��3{ŭ�u�]#c,����J�re]�}˕�����i�`3z��=�a������3T�������`t�	]}Sә��Z�h9��
���e�
�_5�"���fD���S����k֓"n��:̥������1h1�=[� �V�z)��˭W�)���7&$m�i���y"����^�����C�b�7�H
����̘"m��7����m�u8�p��V����͠R��Z�3�Ylϐߕw�X���TG��{���}�����'���D���չΓ��Wƿ���d|I"���r�4���4LD}Tb�=>�b�L)Hxh,�)�F[D�
]4	r,���b~<��;0�F����"	���b�W
g��RZ�ғ��p��3*��
�H�e�QJ�EE�3ND�Y$|i��w�$�'���ٛ���ΰI��&Zt#=!㟜*��So���_*IUgo��ׯ�R����C�wV^K:�O!����[���^lB9p���	R/Z^p����+��|�����w{�$�������,�Q�fl����nw���	n��2��[��AT��t��z8/׈i���.B3�(\�"�_�x���Gyu��G�����[x�d[���`�#�� s!�/\~r����V�hZ|�}��[ҡ��l�'2e�:�J�� �c����c	�3��~Sl~�z�_�Za�/+������@��6V�&j��+�C�r�y.��"�I\���8l{�?,$ʃ�����LM�ć? d�2������Q���I��K��r�(s��b���|�ӹ����]�!�:�}$��'�h�n1��Z{U�x���}1�9��`�Pr���~Ƨ������ )R���(�$��[��6��cE��f[���w��`r�R��
��eZS'7��� ��:�ќ���U+Li��Ş/`\-�����鹊�]��E�p���ah�����[p�VQ�k`ݩ�I���ڙ��u�`EI��k9��!K�y��cW�S�s=�i�������nɬ�Zb��d��o�)j!�PSÇ����[ψ���JR��ɏ���Հ�(��?�c��Z#����Wϕ8�d���j���T/d�]�0G:o�Wc'���{�p���l$)^�/�Or��';
EU�*�\�t$MD�m�ܜ�V�  �5	;l�gI%.nTQ���k�Z�1y�V���ӗ�k9�gOO�w��N��e�"��z�#���4<09��E�!��-y1}��:��"�Ju'cHp��5����\���bF�� �]�\��1�p�XԪ�Է�N�m���.���]�~��M�j��Q�l�oPE-*w���"���p��	�c	��:n���#^6��JXs9X-��1$&,aߑ�T�u�E����Em1����: �Ŏ_�e��P��0D�h��H�h�(�t�"E���V���c&�߿�)������8�2�Y�>�7HV_�Q;�zx�<F�y���NI��r�t��Y���ѝ����[�\k�\CB�f�zE�uu'@�g����r�"�Z�:�z�:��z�n�x�8k����2��W �I���0�A �H
������'j�m��R-�]Ȑ��i�616�N��aeO�_7��7��	a�Ɗ3f���,䅆�j�	ʲ=�%M���<ۛ����P��l����F�_�y�Y<Vp!���.�
�z'/� Ȳ�u��TNw4=��I�r���#�������C���I�'���N�h�����Q݉\�&�zΡ�>Ay��74��
���J�#p@�p��`d$��X �� W�Mq2�c�r�wW�	��1�6۱7���sÅ���MT�a_������&�?d�/x%�ђfhj]|��J���t(��3P ,�1�Ӄ%F8ڇh_#���ݩq�xSU|E-D������ČW,�%9`�g�cF����%����B�'��J�Ĥ���?VDw��&#L�Ece�W��y�w:����8�ӤR�c�Yts�Tn��u�F�EŢv�VB��m���+	�O!�[*'��s���&��h�+6 �^�\���Mc���1�* ��;�&�W��n_��3�����*��U9���D�4[�~���/@�� ��F��	�݁YsF &���+��"�Ѓ��*������7�c �Y)��Z���=��C� �P
��G���K��Zb��\\d���X��(_�ou|�~�Z2
ۻ�&�\�֒�r��\�cl?[%)�`�Ѥ�o�(*���&�R'�Ơ[$�;r���0����n��쌙9p?�����������^�ԓ�3T��Q��V`���-��h��Ey�I���Qv��K@���(�y�b�5�}= _U5z�5�s$|SV��D��mό8)0�Twa�Ĳ��m}�{��� �>�U�!�)[�^] 8,Յy�������v2�Ig'l�ȴ����z}��Ћw�M*��bq�G2�/ӯ�z���{�^^���VT-�UX��x�Te�e͆��i@��V)u��i\g�B #R����{Ʈ3�m,A�bN1eh��l�k�iV� X_ZzW�G	�m�G���GٍI�|=��FT�xrK����}u��l��g�c���h%�_}���<?�\w��6x�13&?�Ҥ��Q�?#�Q=���j��+Wj�>'�OH\�^��xl�<�O:�9�=�cG)���,`�OQ��Ѓofv�����Ɇ�]���:l	�T�V��1�2�^ ��m#k�GC�@��No&�ʉ��:T�o��xj�_�D��{U�͵�*�\��A��������̦���}�,G��ȘrC�%��0��F�w��D���&�Vj"Bט}+�8-$N˩+-�.�D������.!���K	����ׯ��R�-����W���欿�1`��"�_�{�ǹlY�ڥ���R1 ��T��@c��d���oGw�n�W�Xn��]���a�6�q�R~��f��<��C�[�e���ꏳ%�ڧ}q�����`pP
wQȄ�8�Ս3�)'���\GY�
�J(WC4�����ZN��L��1޷v�Q!4D�C3
�ߟ~W�J�������)�v�O�lJ#iC~��O;�����x��[���ҩ��r5���.df �{�W-Lނ�d]��@� �+C� ���ARJ��_�Xc��`�Ba~t`���������uWr�����=7�%���J��f��MesYGҙ?���*|�?B[���2��ŭN��.�©K��>&��盪m9N4�P��+��@��Ti�aT���n�v�ab�I������r�)IK��g!��5b���F�Y�J
"�f��ȑ�	�e��S�f�tT���*�it9��֊��A�KJX�\�ùcI���.��t�LpJ&fe�a��}[������,�v��"05I=JD�?d(�"�|&����:�҆�Ѫ�� �O߽�JފX�;5O�� Ni���ެ���V��rߞ�E�B���钿��d��5�n���}KM�#��t��R�q�0QZSs�ï&�@��2C�+�	_Z'��P���[%2�}��0U{�����&��X�%_����"�� ���+���q�)�a���L�r+=��_ع��q�O0i�NNo=��f�\��R���y�V�H������}�45�S���Q��<�f̒�>a�1^�ۋ>�`4��P}hQֲ�Z���O�{8��#v���)� D��}M��A`C},.� f,��܄-�:�[`�V��It�Q�3F����%e�$r��)�k��n�l���Q�����me��OBU�����zX���R�d��f��V��)O�5�*�2�ƛ���(F+��
Juu�R���	�+}h����q�YY�s-����L��Ӊ�Iy���כ������'����c���MQ�̙���ve�е�g߻��o��? ����?@ۄa�>]��u#���i�%��{��j���bT�J�<α[썭��Nq�8�#�20G>�l0	���������SY�PSe��V2������r;
|��S2";:֨�|��.����3q����U���b��/F�[����RIU�vO-�It��Q� o��rؙ�xJ�9.�]d=l�e��"�A;�����l̐L����G�y3���Q�~����c�q�6�

�3'����]��!nZ��s�	;񥃤��,�ZhT��t��ZBO�G#.��y�̕kS[)��^�z�_��4L�+/y�ӣz�����I�*���{��:����Ej�����}���jplwx�����Y���,2.s��e��l��+�m����MR-�l�|3��D��_�0���o1⋿��8e���-�;S�˜�ZÈ�6����Q�*���
]�Mv|W��65D�g��g��,��6���tcȎ&�(v����sR�R���c���6�#m���H��.�������h�PMϘ�&��.��$|y���>
����ֵ12]L�VG��J���ė�I�s��ȏ�C6:i]�Nk� �����������(8^2L|�������	L3B�������ήM������u=��������R�]�ľi�={S��OA�4��96|ƺlԡ]�*h�T�a!�kJ����m��/�=D��t���t��UGD���h"r��E��}��A�1,y`WR��g�p�3S��¶VSKOU�?�e���9�Cʿ�Z�HCь�2���f����$T�����O1��.�j�O��J�	�S_��fJ��>Ŝ�Ć��������>�	1�j�x�p�"��g���\j�o�Z"��oqY*;���w�F:��V:*X���0�լB�UM���mu���XP��c\B%/dN7�{��,����׳j	�� E?@vَx"�&���lJ���_�?g�R���vbs3��0O��eO善��x�	~r<~@�k�J��.C�Onp����#C瑲?>�r<�i�̆���iǘ����hp���P�Z�����@OϾǝ�I�%�\��L5�ŵ��̐�%�Pd�1���	T��Āu�Z�{�r���H��M�|�XG��G���N�Gn�Wq�o�!�.jش���.t�Ks?��q�� K�| "�H�#��M�K��w�P����E8�n#I0�q�����Ǯ�,=9Ќm�.��>��h�٪�`�F��}lY�߆��V��țs�Dts��������g*A)�&֗�O�񘶱����:i_�D�����}w!�juf�g��<��à�[�'�&��tNM����sV�c���@�ő"��=��&��U��8��X{�k}c��\����r1��~�;��z�O�W��a��(P��5�H��+Z�Q2���W��!���ۗ�����Ą(2����H r�DaJ]*� �#�`րƫwI���q����W����Kڸ��3��<6�`b��-:,H�2��zp�{o��%��y�����Q� ���Z$Q����{���N��_2W�
��ߎ����ԋ7�4`P/��T¯����|a
N�t$�Nk_�Y�D���1 Ҩ�\X�h�?�~r�<����7n��L���P�x�C.1�" <��5 ަk��	�j���[�9�T���u������o |����Xd��_��^&�z� �����*��a�l�'��Ձl F�4�U�]��O�C'�Ո@I�54���h���4?���l���Bp�z,���,\��i
7��Zn8{�+6a�R_���H��9~@XubO��:m�)�	���N��m~�RHR���� n��s:���g��/� ��b��R�-�rm�Uy�#vVM{6Ӳp��'�dͦ���(˚U�.�v#�{�6o,7��/�f>HF$��1|��C�y�~�LU�E��.�C�^]ltˡ��>�Jp���h�[��.�!h�^z�[���$����rGj��乩�i wS >��������=�@�c9t�_b��o��3�?�j�[�P?�^jWb��+��kb��`��������V�
aNF8;�^ �r�nz��J"�F���	�'�܍>���[^��d��x|�A&̧�齟��:0xF�����c"����>����C�J�/(xc�d��¦��`
\N���0�u�@k�X>��d����-Ö�wXC����M�� �أ�bJگ�]SA��[}GP8).�dD^c�� k�_7�/8��IY_ƍ���g�����bY���"G:��A*��]m�ͯ��0�y�+3T���%�9�3�ԑE�3�5��U�3"񋐻�3�2	��*o8��}��Iz�n���9	�x=M<�z��H)��+H_��c�s��u�(S����3t����e��׿�4$<}	�4��u^ �j���g��X����?^��n�N��K����( �o���(}t�ٍ��\���5-JǱ�!�Q����9Uj� ��"-��p��]	v�'YCµ&b��F2����K@�bG}.����Ϳ\?�����6�2�D�����_��e�NN��0���� �H��;}��J���{��RXf�;U��S�=޶��H�4D���)�}F_�T�"k���d #{��Ox�eA��Sá3{(�&�t����Y�,B@/xޫ;�<D�)FKgT+ð!� ��w����Hq6$�Ed�([��/[|Z\d��6;L�ǝy���R:�y�fO&�V}���3�F�\�Xݺ�S��z-�M��¥Ku��˔A�)tzݕ�M��0�2}a>� R��zT��o���k>O�f����6%~~0�)���^�k�t���������?��/>V������1������kؑ��y���_9���2ͩ����oֹA����ĭ���~���{X��TTjKP�t�������
�\]��g�?Xk�&5#HV��FA=V9|z/'�Rmµ��Mg�a�z^�4  u�l�����0�����4�c	i���%W���i�����KV�T��g^�!=Qw�1�b�j>L%Q�	�����`�j���h>5�b1y0X��eBM,�b�s
V�5z~ƪ��ROHb�ļ�����\VH�-��jVi�&K/Q�ݤ�	�|�̱�?��=a7kݖ�D��Y�K08��	+["��#�ޭLD��Γ\s47���@���� 7
�U$8�NkYn�� =����!���r����`��W"
Sv�j�D�߁�<v�E/9)�SΌR����x�LA=��T�C�9�B�"�:�]�8{&���q��8ȗ�`�b5�|e����K�݉u���<Ryc����+�
H��Z�BI�(��B�!ǽk��Wb!��y�"t�Q�R��jZ�r�9���1s�W���ƌ���;��4������Z��9v%���Р��(qn��8���/w�	����7�Tc��!E������P$�p�����C	�ۿ9��ٸ�JPr����.�Lڙ.�,��Ԝ&%��	ar_4�l�1\P�����[����,GH����ɝ,^�k�R��fkR��Xj�)��z�%ݞ�E����.���\A����^�ݪ��Qa���6�^��HFd1WF�W��֐�ΰ���c����<�%�]����cA�~,a�/�_�ϣ6>�f[�n{H��3e�bf�"�+A#p���M.�"y���tU�>�綸��|Z�&��=8韗}9���ZU;Jb5����N�\��G�6Ź$�O㜎6<N�+ν���6|ѕ��s�!�ɚ�ة���$QJi��u����;��!܈q
�.��=�����g��g?V�7PBC;��
.�p�la��d�'q�vk��`4�nl���\|*���G6YVu��z�P֡�$=1�Θ��l�t�|ܸ�̱*��q?�<9��k��)�!�CI77���,J�#�+� &թ�P��>y/����S�q��'�:)���xNG'�YK6�:1���8��,�NM�2 �@*H�T���-�ԫ��P�Z߃���a�	���r�+Mf�Ş��X��c���x�ǘ%���Ep�R��7Ωz�Y�y>1R2��!΢@�Sç�#'�	vg���<�����`М�#��Ե�>l��*�a�,����_��R=�/AF�a��K6�*#�ZNЂ�i�Ӣ:V�u���i=�{ܔ@#���+�4����#E�*�p�PHo9�@��|'��v�)˒`����":]�Ē&p}�8��zR	���#�L3�����3��P��~J���Kx�U��D��"���~.��K��z؏s�#��N���j�MI�&�Y\���?;Vu�()��\��8�Ǳ<}��_����l��MlH[$�͙�	�D:��o�����U�H�?����R@2�@�{�a�
��GH7����y*�e��QmF�Z������Bs^�c+ێ��]t��Fs��!|~oa��!K���֘�@��S�j��� |*_��ECrV�Gl'Z��/W�]!�:6!I��wI���q(�ͷ;�;�,B��ꅛT@���'�u3O��<�T����~��_!.��ݧ�2�����k���z��Y�����)0e���.�X� Պ0��d}|�����79�d\Z�+T�]r���t!�(���S�l����2��n)G��g4K2�UݹJ���%pn�S���I�)*�g�� s�R�Q�tq1c��rd x��_�zXO3��~�#�;��C#������7�v����[t����m)\	c+V��A���:<��Vx�H�P�M#N������ߗ�lnK��
�B�<�ڔ�	���<b�JV)�8����i;� �&8����_Rg[�V(���p� �ő��I���*�ߨ;L�׺��'$p����p�[o��Z�,_��'A�U��/�(p�'?#R�l��4����Q�2�T��!na�_H�����U�.�Cy�~tgC�Ì���\��@yC~_L1Ū���vj�r u
��m��E8ۚ	�z×�7���o���g|�*����Q;��%ZA�`�)�k�槏���p�:K��R�A��Q�Ě�~�G8�X�H,]5rd���EEO<T��I6J��\����G:Y���i �J�F�ez�g���Dg�N����[������i8���R�i-�n�]_�-<�-������/���ަŐ��(�-lA��$w�Qs��RA���ug�+4Zɽж�h��bq� F��6�MŖ�T�csPE��u��_�B^����"��u���1�;�h̚�?�o[滻{��0hʓCAS�@J�;��\�[P3�6Z� ����Ƴ=�ϝ�q�>`H-��p&��ϴ��Y�d�U�nH~|"�m7k��F���Gb!�p�A���Q@,�t0S?a�BF�i�}�M�ϵhҫ�wg73�t=4x�°1F����J��������`O�����
Q�+�����U8�#�RF�I�đ��~�n��)���N3Bs����=p�T�����w�N;g��?���S���,K` ��uݑ�%�ܱb�P�Zޓ`X��/�s_�Q4�&|:�,dH`�
G�� ���%�çedpI�G��d®d�@�^j��p�We���K���\mC��n���WT�o���q��|w��N�2	��Z���gz��~���ga�����g/�_c��}���	
��g��v~�����5XJ1X�~���>D�<h����V���|�{P�r��3��~�gØ��6�Je�^��kAM��Hd^ ����o��b��΋�/X��q��Ak
gc3X筹�{�Ɠ�e� &R���`)xa�� f;�m�x)Q��c|�t3�H>7ҌGj���~i�8��a�G2�&���p��"�1�٫��)�����3���Z단��9W"n�㋄��`�F�d1 3�5���g�j�Vf=�	j��F���g�
Й|x�1v}�'-l�;Z�i�������ٚX���G���6����C�*���IR$��/�P5����k�$��a����*3��Nd�f
��s����	A8p$e[��D,�Z�v�2'�%���ams���+S��� ���@�����=	���۪Wj���C(�����V�c����S��C|���u�׭�;VpA�Ɔ���J$w����L9�Ր�`U1�v4>2���YUE�扙&0�?s4^�ζ}��������HL�"����a9��z�4X<��kGr@HXS�|�}+���t����ى��%�M��Q9L�A�P���)�t�[A�æ�.�Ep؎�H~%�ZdBBP�B	_�sk6'=@=����a��1���Q�ޜ@E�&�>_�sMQ�/��'�NԎ�`�$v�pgR2���#�9��*��!cO��,Wx��#{T�ꙛ�ڶu���T�R��t�����H�!d͊#}T�0�I�h��F=��i�;B���<i����
��m�d���fFg9��`�lg�:���W�Jma=1�����С�������� ��2�O��R:�p
[+� �qrc���s��KNV/�w��!��{�����t���КL�t�҄��'n�2(z��
q�Y�5߁t�,@ɛE������LQ|[���T������\��P�����=&�@]{��Cfckv�t�(n�_�{**�����뀠��p�w~C�io�Wozg5̥�u���n����-pAFv�+YIM��<�<�`�(�l��z%��L�
KC�Əh�hT�D�Z�N�K�A��/��E�uVyhQ!	[� ͱ���ZV��"�(��cie�B�5*im���˞���[�-L}��k&V��9��//ϕI�����=�	a�|
Zo~�}|]�6x�.�v��,�V���T0yS���'��������J��E ����\wNn|����8�:��a,���A�w��΀7�0���U�<P��aZ���A�*�:�#����8^��J#�����G�aޠ�/�T�6���"�քM�<�j�`��rXĴ�TR�����O~��\��-Q�'}���4RPd�^m}����ؕH�uA�)�sγSJ_�S}�)_0<;�7�����A��i��B�B�Tc��`�������8D�(�fK����	��ꗙ��.�].zRf��=�w�Q��JV7�f��t�i��A}A[S,G�ck*%+�c�Y�X�(e�0�=g���}���/��m���Ȑ$�i9�2>� >��'`䴛��I���j@U�vytqQ���ًcU�5]����K'�r۲���(j��5��{�~�ܥ ᵲ��*�\�B��R`��%?��M����B.�d��� c�TW�Z��X�� t���ՠwz䴊�d�D������+�M'mu�h��>WB;Z�
|��d��-Z����#��&���S����@8[Wb����j�������ہ��E��D���2;3���^�8�fQf�.�:��l��c]��f]�/���t�������L�h7Iӛ%]X�mZ����[���x��Y��tjm���t5M�ftL��,�y�ɠu�h���u/&����Xf��J�=�A'���u�C%�6e�����62�^�w3�0�&k;��f�p�>��G57\�nf^�C�ʛS�O(��
��LN3��3
��\�9�qN�#���l
{��/��=L�!�a�7 p��iP���o�5A��U��>A��ٌ6Y�r^˘vd��#�\f��C7�_l��N�Z��l.�g~��  �/��(S*��s���k�:�u������\�=����ruZ�"�
�V'��'h3��j0��_�C"È&Sĸ������!��ZU=�P�]����i�F��?�6�懠x�-^Ѿ�{��Lx@@*�Q�fH3�Q(p "��J}�*�-m#_�F�m�.�e>N�WlMZ�������w�גQ`v��&�EI:u*�y����ȭ�;ϓ��>�U;�Rv�~�ޒEl��*&]����߉O�JtTO�P�ɗ�Η���*Ѩ����|-�c��)�`��Kj���_s��EsjK?J��$����䔲2̆�h�bl��g�m�Ta�,�V��*4x^�΀��S���،��G��{�D��P�8�X���:\&��yn�%��5]Ϲ���q��z6�8Rܿ�u��/l�Hk�@Z
���L�?��P��>�R�	븫������T��N��f�T#^J�A��ڦ�����;��=�7/v��u2>���2���L�&��rQew�6Y�D=�,yc�%
"Q��X��U�^��bA�Z�6�g_�����'���U���x����	.6\
k�-�[���n�_�U��J�д=dd�F��K$�Tϊ�F�)r�i4N��z�C:�,��Zt��o��\Y��ϊ6n����`C,����io��V�>�+����I�*�=[��P�R�3����f�Mrp���w��Q_�;��E������p�!`�q����~��"�(�"����oH�`�.(֞�����8��X��k�@�u����#l�8�ו齇&Sx?�R׫)�U���9�I�A�����,m�H������f��]�F�FFr��s�u
���*���Ü��l-���~���en=�%>����>D���Gl?\)���g���-�-X�7j�nϑ�q�P� ��7K�"�ܲ�L��m��b�l�����e�MG�e�X���[Q��2���
*VC/���z�瓎l�����</�`!r]��]!��V��r7�:c�٬���v�
�w�12li�d�f7���A�hGD@+�L�/��8G�QQ�-ǥ	��3�ldp�S	����c��k�s��]nl�,�:�h�+��rp{zJx~�[�S^����?bUp<�]BV�<����rpiP85�Ds^�w����Ѝ6�z�7M�Y*�C���p!�N)ٛ�JW�4ݎ/�
1ԁ� ���7⾱ ���V�xq��Q��p!M����,�K��E��Z����DZ0"_����
n�k/Ycj��~b�i�a�ڈ�O#�PЀ�lF��<���.��qI⏜Bkܺh�H<�ċ��_uQ�Ӈ&������@��Y����X���=�xI!(�D�Q2J�:��Hm�lgTm�F��l������XG���]X	��چ���p��T��u�p��9�p��"	�2-P�-,�Ӹ�y;%-�M�*����{�?�=ز7�5Ca8D��҅��k��O����E�7�ef�?a��D�E��D�Y8��J:
���z��J��x�]fdB����4{�+e�{`�������V�Q7�4��J��3iUw�kc��*�&��/w��S�djhM3�}=�'�*zw����,����3rB��l��֝��=I�]�sb`�h!}�L�S@�n�]?�g�柏�r9 [�_��۞_Jf��Ȣe*,A�5�tb�d��R�'�[X�I)�]j܊`[�gp�O��(>/d5���'��v�Y�� 9����3�?ͨV���X�>kR	`1��+N:���H�B���:�]�wg�!Bgvc!��(��M�%�ܥVGo�*��9pt���	��q��(r���u�p�6��0�xMV�?�*�����b��C/�coG��%�E%�.����.dX�Cꜗjs�7����Pu��~3o�<.�d�'K��veyݥ+T�g�֐���Ca2��E��[v���YΥ��|Wj%��c��Fx1�I�o����2���e PSY)�̈��<�c��LP��Y��[�^J��*{��5�M�'�Hr�z�2��Φ��~Y�Y����c���y.�h��U��������Uqcφ�`�����v�c���fy: �]���5Ý�x�;�1��fqK�;ʨ���W�D�5��-s����7��n�,;7�#2���Z}hx����l�7�Z;�2>)���a�-�}�v�s��E�8����r�f s[�Pq�k~��_��[WjbY}�1���Ki�֯;��,�@0F��X�����,�c�G���7��L�]	s`!��M5
�}�N�M���U�ڳ��Ad��~�$��p5ͩ����/�bK$W�gh�J`6��[�sN�_кd�� �2���t,g�����xKC]�)���SF�Xq��p���3_��*��%�0�.�^�̜w~ڧ�zNEi/[.��VF�gHD��E%�8�G�Ǖ6��?Qɮn�678D��X����"��ߋeI��R�B��VVM#D�W�3���
Yfg��r��Zf�^p��CzEd���YQxNR�i_�]�z���
��nZΓ��=V��PwgL�&t&���I��SǬ���$�DY�%s�+��V�����A��� e��g(�,�g��7��{���q�{T�	d�uV�A���W1�!�`p�ߧ���7xܑ9�L��-i���Tk����
T�S⥬�r���D��Ym�
�� !(:�yѸ��}��p�%༌~�`�]���ɮ��(_m�%Ϣ��- sO�� �dI㖪0Ȓ�i%V��d�ɥcYN�֩KN�k���2��H���{=���Lz���H��٦d�4f��9�##o9�vZ#q ͕�JϘ�^'7���9c�[[!�(, (;���(��A#d�o�Y�d@�#λ=I�k&=���0`��m�=��i�|���6x����x�X+�l��8b�¬ׇG�xyg���÷n?#s���ŀ��ظ����z���]�E?!�W������p�.��N�yU��#+�5W���\�]�K���9ކ|uP�Ɨ��9�d��W�'h�s������� �(���F����~}��l�L5�N@�D�� �1ߎ.J��SpN�ɒ��`uW���5��z�����2��p2��
������Tey4M"���u!+;��q���w�|٫^��+�?���Eޤ�H�A�	7���/6x��5ޤ����`{���2�V�	�M�r�"Ѩ�+��r�Y��\�f�IY�{Kv�"�G}�@���w�%9�(�J�5�h���
+��A�I}6ͬ���;h!�Tޖ�bM�D����+X��bߪ�D=L
�Ώ^�.]�%��~H�J
o�����q~A�+�� ����_s���*������ĳN�v�� ��f���<����l� ��>�{��$�H'�b�5���?,�!P�8,[eG���I�D���������|f�e�H�=���Ix�/�Ü'��ZRe�HS�th�ht�\4cU� b:tt]ǈ*x�je�۾�+V1 \T*fM��Z7�3>�h�
���!����w\���<�:�z|$e�@�o�S��*B�-%M۾���E�!@�"vV=������=���p�5�G�1 ��''�Z�>ԩ{��Gno�ΫO��ǳV�تPѺ"�K�m�TUQ��7����m}�AG��x�{�����ӿnh��Ld����5O���D�%�BN�a�V�CW��u�EJ��$5,�9#�$"E�0���Gb��K�bWV?�N�(��P�Q�I�;�oa���T5*����pίZK�c�5�R�וŨ^V��N��$�bt��<X6c�d�;,��#:1	Ǿr�x�bG72�?f�[�1t�na�H�w}�%s�#S3�1��3�]��U#������ZY@xz�Ct�i��.�S�"Vi� ��>�#��7�J�����MQi�\j�ö�i�}�o������5B�+���q����1jX����m��{=U�SK���0
'��wW�k� ڋ3������QAFF��%�)��F����1��ʐ�T�6���Eg���|��l7��k�v_�/D��O-��YBL��lډ��m@�N��5Ӭ7g5:�-�rx�@%f��=_󕌮Qcͷ��qX)�K7�����;�\��:`[i1⨋���{I�'5J�m�=:8��}��	� ]����G�n^�{�)�*��|�T}E��y���ѫtC�jµ�ֻ ��"pT1������cVr6@�������Bu|�� �X&�� �0���E.��@�f�D.���Ь��$���Z�f�x��Oac����auFЦ9���xB1���x���٣0?�3��SJO=��d�B�r1d��k���l���Ak�;h��o;��1���y�S?i�N��䟍�S��q��0_CX.9���HGTt�e�d:�����!��>�ͩ��A]�|}�f3���Ya���/��~>h�����yBW�G�r3z��(��C ������ &�"�铜�4~�θ`�M��H`m=���O){*J�����P�-B�4�{C�rl�a����U�~� ����;��v��<��&����T)j�.�xf�^��
��L�&y=�iJ��1��\Jq�
��WS�iK�Ή�����=��p#tM>rtj�S!zo]����8� �e�(.,y,#��C����Y^!�Go�#x�a)S��6�CETCA-��ӛ�c.gC�s(��2�@U�ݓ!W)O-������P-M���BE ���?�$�˚����I���Y�� /�\�:>{��SGR�k>�*H��Ϊ����RLmR᭒�۩�>�8�5e��n��()ߣ�3�(��F���y����W��s��/� �Ɍ:*s�޲wũJ����9���V���7̹��=�k��w��L&�(X>�k�K�B��3�Sg���]� "!ގTP���95�����-�ȰeuI�����}W�J1vS2t�_]�R����-��CY1��@��	��7R2�/�F'�l��`k�����zվXHUI��n��0!$3�_�f3��-W/� �$�x����u�|��J|�k|uQ�5R)�6� R���yB�{�;f�����Muff�16�T�l=����p�-��i�1�9S%�*`�ts�1��$���3�S�
Z�m�;ƭQ<B�Yƣd��x~eT�R.����$�9td\FK6Cc[r$E�7X�\���1)	J�Wi��}J:�&�I�y���w'�5�$�Z�fy`ޮ�0�^��o9)B$d�S�g4Q�op�41�H������D]�`=�o��;Cוg-U�dLP\f6��E1��V���Q��2��
�b�Yx�	};�ir}E�Lh^4�L4z�
=+�#�,X�s�ц�W+��#�_�%�?�p�/�m1I#�����/��K�y��݂�ۤ[!�^�)����J�lVU�YSs�P��HVaƾ���t�4:V�U<�v�Z?��|3W�.	 �s��g������H}�Ѐ-;m${L�ɾu�ܢ�7�u	л)����,�N�[���J�
"�D2�	�"�1u߁'T���+�����JvV~ۇu��R ��jOM�?�M�V������C� ϷJMq�f�t��;���'���m�t���H����n���y�ԯ�S�5��KN=��Q��p,�y̝��2�Q��<�%����(�\�K��'M����i#V5����q0�j?3�����1@�?/���%�>�d�c] #9N.V�����a��x`�ێ'ظ���1ꂗO%fؓѱ	0�ft���깆&�lՁ�b`������nE���o��J� ��]⦇��p!6e��Xb��6nV�А vܞ �u�[�M�̀���Ն����������$���|�V!�����5�)�*���P�V�����	����Q���l\�.j��^[e�m�Yh�g����v�"/��qb�b5o�(~)�8`�*���O�>ف�^	d�ݑ�7�J[���dJ�� ړ�ԫ�ȅ�4��#��h�b3OF�����oL�DC����ؽ�q�ąs.zYB���7(`�m�I�4��w���kC�3F�k@��D�k���Jz�y����:i(�v�/r1�x��XG��%Μ3m �Y\l݉ѡ`��������b��cU��r��^�FY�l�$f���ٝvCb;��G��m��޵�"����}R)ծKCh�����q��5�e�Y���_����*��o�aQ
��i�L��dϱ8Ǯ�0���䮉�����C3`�&��K-(V�%�@b5�`(���h����KꪂTy�C�D�a�t��l�VS.�-$�|ꃻ�N
�9]�6_y�m��N|�F"m�����~��]��6tG�m��/��b�t"E�y�&u5_��~��z&��]�d����X�2�,N�4�=Ϡ볢\�ɀ�����+�Y��`92�Q{B�D�($f���dYwDD��QtՈ�(v@J]�X��������'F�n���,�'���i!�����p���J�5ѐ�i��ů��+`^3��5:u��~_lw8<p*z��s�ߒ����Zԣ+fzS	?��1������I�s���d������W�#T�]4DG���Z89�`�S2�6$����Y�����G��H�E�b�!�B����>�����Y��5��&���dw@2�Uܽ%��=�@���p�Ȣ&j�"���rD�;�B�j��?.L@�B!h����� �ЍSE���9��
DDYA��hyw&t�NO�YC5pB$�����!�=�!=hF���B�`*�'�;��f��>d&F1]ʄ)�5��\&�V�����k*�CFۿ��V��pْА�SҐ#�-Ħ�2��E�t�"��_��1�t�_)�������`�a�? e)VR�0{��)B�+��� �"���z���j���LSa
9�##�){D�B���㸚?��.�B�!LI)��:�Q�v�4�!{���E���qDU?g*�O9z�,W��jT���X��� �)mo���J�H�_���[�6~ϓ�a�y�#?R�ud�T��r{$�fk@U���|��xfi;��΢�[3����N�����=�q�bs�7���Vl�#�-�K�N�0:�x��i�l���coe�(���hÆ=�# 6��.�I#,���\k�')����o�Q�e ��R�k��hH�T�A��T�չ~H:�ر�O��~�/�<.��x�����?�#��'�|�ƫ�m��}�sp�	��?�C%k����J����&��Q8w�4i��̔߬���$�D�Z��� s�1[��/+�Iٽ�?y֠a�^d����P�GI�E*����O��I@�:������-GC��ɰ�y�`G�.�L��J�9��_M�����@V��Ӵ@3��/sr��܁]Q��5C���n�\'b���Mm��?������x�Tz'x���'0S�h���dT��N��N�9�g�E��&�)r
,�+�����SX%�����6V����xͳ��?c#������j{��X���ޕ��9���m}�1.w���J��4X"\��xY\h���-�����P�w��p��^t�@���A.��|]�|D�R����4�a ˠ�&���y��;v_��������ضV[�olk�ڱ1ydM����p��7�q�^�\�֓+5����hL��3x��O��b�~k��X�BT�1����l2XC69	�=�nx�h�'�X�*���L���C}Vjz�ar�8O���=������8���"�{�n�Z�S�K�&�;����|�m"A�5U��D~;���m�u LEs�!\{�@�:����im�T\Г����0a���Z�����1�nbV�v���D�0�
��^���ʆ���ۊ5i3Ҝ*�!���Aw�a8w�U���"Μ��QR��YO'ݏ�f���k$�m��w}�B��>�U�z5�P���f<�Ђ��JR�֔m�wfzV�X���y�]a�+�mm���x;���	~�6�3�L,������;f`JV��%�C�W}�-�k����4��̎*%�N����*m���|�G�i߾*�孁<\y�Z��No�QJ��r1��X�x#��H��C@�r8ayб���p�4��@5�X��zVRM#@�pԾ�icc�'�E?��J"��L��~�BvR���Þ$6X��s��!��m/�.��C$����%��f��>�i|�:`Zr�[`i|M�%y�@}�əR��[\dq�ހr��. ��)�˫�>��+e�۷�<� qDM�4���S�x�.k��>9�H���+�p��x�����-�ʰ=�8�f2I/��6��ͼ4�� lV��Ã���y��Я�A31�<���b+F`y��lO#o�[Z���O�EJa�i�l��[��ZL���Y���뜖� TFA���5����j�~B/��*rB/�E��Ԣo,KC�e�u�޵f11�Un`=SJ~U�+������9{�0rz7s����m���R�z/�ˏ�\�׋���d���!�!�󗅆r��߈+�Q��u0��b�K{ �n)"��|k<t��1A���$z�j��i�>��6d��,�RT�$sk��{ςf~�k�LoQ���H ���NҌ�l*nr�@���S'R͎�g���n`Z��!Oh��Z3k-�kQ�MS7�C5W�s���`-��=�]��`z�j���Na�,� ���t�nez��M�ȝʳ3�iy^��Ϡ+.i�N	1�-��F�$����o�v4��{c�1f�����}�&�}�m��^NpG�;i�`�ҵ�п>.��@�C�Yz�<GLm�3��OD��������k���� #����pA��}��.V���w`�s�4o׋�iҋxz!��f�"�¾��ܙh����Ƥa�9�,1	
�,hel|y��L��4�j�S�M��)���}��s�ؗ��۔Hs���W
��}��/�R��-�k�#�M6r=�W���h��nuû?ź��[pL�i�Z���Ąߌ
#���&�շ)��f�s���Pv��@p$�ea���Ü�/���#���1��˹���;��@@*d�MO��)��4�d�
����������}xjH��"��r8�,�[©?����ן��f^�l��⾊�f!��uoL���\�bqsd�>�r3��;���茁��6z��,"��mp_�� #� ���E�wF#w��[�F��W�/������=r%�S���;ߨ�C�U p�$z���Ҍ���Įi�8��A+�`�Ϛo��󊝇a�D�E/;[l��7b.���w�6���<��0�=M�z,�
��R�B���o��/.�Z�S����Clz��m3����z~�X�c�e��V��K?��H�~$�����3��>���6�cc:�#�vdA��'7ҽ�O���h�٠4ԛ,��UU����.*�m�P�d�h�=�����8���YS�a�o��f1��ty�j1�My�D"��]ń�,0��&dPk|xd!��^���<a����Q��aZ����uV���G��^\A;�>�I^�#-�	���S�ω᾽��m`�`Y{�v��A@t���>�Mݨ8��������7��i�.i�_��p�߷v����M��Ko��8K�4�<Y�3K@*�o��q�f^IP�( 
���Ng��(�\����Al]�@+m��
:/���R:iP0�N�9�p��VwQt!�~O��$v\9���P�i;�&�kC"@#��牄���I?�i^�Sv�I���5<ܴ�1��uD�o HjP%���x`�x�kNW���:mj��\Q��l�
�&�:��ɖ��5�� �b��R^�L�B��25Jk��Z���)[�_O١dKN�y�^����tZ�2����-���[�����<�T��������x�ܮ�L.�����/@�<��	G0��ɀ� 9s��*��J/�Fq���L^�/9��l��Յ��"&^z\�[�ųQ�F��&�ُ���
����y��CH��JN/������e�*��Ρ�����J ����B�m��uh�G9c�l�7����-�?娔퇥;��O��$Y֡���Y{U���a11W�Z^��Ҳ�ښ��`�G��E,&����毆���g�=Z��P��$��¾?�x˩�I�d���=Z�-)$D]&ʐV9�R?뜥5�Zy���_x�qɅ�(���%��\���Aπc���Ω����J�
-|r��[s��2�?��]���rQ��;�_+��ե�^D-,am���x� ��i��]Z�u��J�\��˱������m�����s�ؙ$ե����iw�W]�>�}�9̔�l�lF�@S��֓>ؙ��[M��鵊u�P�\t����t�V�2Ja�F�d���Q�M�;)�t��嶦�ա�}w�5$3��t�Rj0�<?�&�VǼ>l��N �8�)s����T`����eyp�	��
8P��qv�&��UhSC�'����{i�O�������7�1'}�c�Xsx�_��&��R(�8A�;����Ed�e9U����d��l9"H�Zp�b>@[�k�Qrx�,������Ec�TwT_���P����k���#�)�:�!��څra!�1T~��
�m*��c{0;_ �<W���2�v?/T3�1���S�FK^�a5��)m��U-����X���:�8M��q!A����sƒ�%27��a�"�w���w��������	�ʁux���d����-1�Z��`�D]� ~�;H���\��(��� B��K�]~.(��F<����9����҅ �	�h��ýx� ��:��OA;A��R��9��UHc���ʷ%�S.AܹM�*j��T��}=j���u�"q���|k����Z�(ehp����¢f��ɂ�L�p~֪�\M"�V�@bx��4PW�s;:��~b�v�k���ȳ�՞�O�h�Y��+*M���������8y]�����a�Hʰ���>�Hׅ�
.N\�2��̖����	��Hn%WQ�H܄�}��|���@��ڇc�>CN;��.��y������j��\J�:2h{Q�a��ǰ�l�eփ�ڥye�����l��!۸g3¤}��~,���U~�֑u2��Ì5�Q{��fK�`'�K�����(�{wߛׄ;��8(-�i�l����6�^��Cς�+'��F,;[�C~kT�L�7�p�����&�,}��K��M`�jW��V�(��Z�XH�g����7?��IE3!�u��!<�~1v����=�(�+��R!t��ٖ�R;��ZG����
|CCu�����#+ � ��"!`{�1x���>��ٚ����*-s�1"e�}���:ܢ�hkܮ���0����Ѐ�
;n~1�
/m��]V�����-�<�$A���P�Ms��%p��"�o�e��J�G�Mf�O�ܐ6q��3�����#� �%��l�h[Q�[q&�F9j�@�\o�~��x��'�����Q���=�Lv�&��u���J����+�\Z�U�"�)2�
+A�T��(k��U]����$����x�v��&��w����x���fgڳ)]�(h�{`O\�����s;,�� 7-np՝����O�sT�__]�֫ړ�yn&���7�ͽQ���rk�5��ę2&"����'G8��k�j̡�v�GvPf�۟龒�Rp��NE�z	�Oy�� EN�C�&�8&j�S3k�j}y�o����ÿX�T�O�C�&ZY�@�������{�Ͼe��zV	�!0�&���\q�՘�U!����YGy$�
���J��3V���v"�%��3��Úuj�c%
�%K�G��Ã�`ϡ3ō7��'4��ze:&Ձ�G[��^��bN�ta9@�*G���L�Y�%J����  L�,�?�J����F��b�*(0��i��/�Y�k)5�.��IG(cV1Z�/��ĵ���/��*u���[�U1��0�9��cQ8�$;7���ҍί����ɓ����Q��5S��I׃�� T��/�% *�.,�����u�a�x�����R�2�V�H��#;T\V��4�:?�
y�"�s{�]/z7F_D?�VA�j�j��/��	��\�`�j��tM.�LӀ�y��"�5{�v�_���@�!�FO�=(Cqp��!�� b��b��%ͼAZ�<Bj���)SV��s/�eí��^`��@u��Kj��M�%pĂ�	>m��2��.#��mj��8�hS62{���o��wɻ�~/5�֠`��ރM6 �y� Q/ރ	AjJem��*ʂ�0�E�r ��m{ݦ��!�i�bOlo鲿,`*�ϸs4��sTQ��r�G�htA9�i!: �밁�a�˧n�
^�ܴg�$QD�ZA��ʙЌ�9��|
�����b
�}�͒���"�	��8l��\O&^mܶ>�8Qak�gr��BsY4"Ux�w�^�J�w�>.+��|S�z�Ό�D|sX���������ac�(�!a*h��7.���ܠ�֓;2�@
�b:@�T𰓻�����]��Z����q�R[�$���جQ��!��qIԞ����5���P[�f��w��$�+�+>6��z��L�^lwzʤ���`5�$�?U`n�u�4?�^8�I;eF���}|��0x n�ѫ/`L��5��Y���%� -r�گ�f¦���%��ɈR�]Ł�ǉ2�z??��Pkj.�: �t���>�ҥ�KL8BѪ#�t��Cޜ<YQ�����ɛ1�۲�R��.&(�V�����m��%�Q��J�I�%�<��4�`�㖲5P����/���q�d�D��PI)��G�&[Pj�}_&sa��Y��b;�X��PrTP.V��I{�h����E�{�1����ݰ�$����-��s�-�i��$Hf��na��$�0���fF�4\pD4%���Kv�n��,s��s�Y�|cZ:��dUnSv/&Q��R�4�	d�HK������p���e>�Xe%�P����\�6d�5�U��HN�9���N5	/ҵnAX��ڭ�"K�W�EͫWX
Bbu*���O9�՞���>�����ՠQ\$�:r9�W�ek�Q�~�q�آDv+d��0\�	�c_�M���#�L]A'��N12��W`b@�������%�"�E3i�"W�^����>#�����B$.� נ��/Id�;gF�D���wKĴ�k1�C�q{kӥ����z�q�\�=�����f8�g��??����oK��5J�j���o���F���r�:X�����3:�����P��5�.�@��]��ԇ!	���`(Vo��AuǱn�8I��L�ė�0�s!u�J�W��g���հ����
� ����x�kĞ�:����<J�.j+@�z�jf�D�:�`��7���Q�U�{�\�DD���
���G�sj�NaV�&�#��.�U|W⾷<���*r��!����ܔ}�~�3nQ���8:��<�@vr��vhZc�k��̮͎[Ӗ?6{��h�nZ\h�L&�� ��%��Q���jKj������a�I��A|�wW��A�t� ����SK�����Y)���p$;~�mJ��{����'�������/�&m󸰃
�N~%x��F4Y�8D�3���;T7�̄��T7�藖i�~Ayu�*p��=�~�hi6�w��_�D.�8}4~��h�w��BM�q�	�T:�I�:����gL���S�^$�}GM�R.s��XP��8��CCR#���A�&ZM��d$�$�c3�Ɩ%]@�٪6���b���XEi��,�?BDa]�0�Djq7���T�e,^J�0��Y��{��{��T��~��Y�Rv~�=���`��s�%��
��+3�	f�pD*y䒑�Q��\A��^tq�<sv_��0B�m��8�q�,΀�R�K�h꜑1JG��ū��o_������:�h�f^�mƝ{��	����F�GYK��4�ղ�	�#`ν����o�>�;�<�:h��2V?���tW��_�;���JIb��%��ޏq�TI�t[.;�˙Sv.�)J
qa���F�bp�����3t	u$�p�H��Y���]�#��ިڃkF
����ܮi(o���\(r`�7�}��jT�L\���Ah)ۡ��pF��=�P�M߷U5k����DN��W̐�K0�G/E�`҆n��{(��܏��I���#k���[8�<`��_@���fr���m6
^��Da���2!�+�DCt�����od���n������fOk8
�N��K�Ix 9I25y��Edt��'�~c��	�����x�ݰ'tG֠=a�L�ZRЏ84�8�����_8�N�ꙸO��~0�+�KŖ���|���A�#]ubN��>X��l����mn4´�
-%�;<4���%�yd��mxܒ�vCM g�pp�����@?�]W�1�7C˷��gE��k}�>Ϻ��[:?��-�\}��*b��y��,�P�ݨ�a�@�D_1����,��r��>)�{�ג���l��G�,saWؘM�∝Y��g� ��6dG~��q�iզhL�|=>�̉��'��&YJ_��+�>k@\7�$O8�\����Q9��=h��]L��=p��j\%�I�%�8p,`E�I��N��}Y֍$��Ʃ���ah�N���b�4�|�tr|7�Ew&�=�����JM�lV�p"E��,���Zގ���S/�'���Y�@����k�?�[^�l� ���15��Pݦ��r#��.
�$%#2{Ɖ�E�U
e��I��I�Y�1��T=t�� k�)�GZ%(����8`���7Xj֣Y���fm�@�x�����,~6��ӫΡ���ŏe�7#[Q*b�[�O����x�e�/�"(����,�������Nz�%�κD��:^��Y�A%����x'�R�$ϣ�BiM��n��EY�Nm����Vͥ��lhR��7��l_S��|��� x"�#>�9�]M�0���|1�X��DD��}�)��%��t=�D�Kqy+\$�ό$A\�f0d�z��F�y�>��-k�� p�σFAp ���Y[i1����k�H���6i{JFp���NY�W����Ӧ�L�-qe җ����	����9l�H�L�x��~�Ld��'3�୪�����<�̜4����HCR_�~x����=�@�cy���t�;c1D�5�\��u̝�ܯ{��~g�.	�,6��yV���:He�ÿi����I����6�@�'j�s�x�p@8W(��]���6�P�磸o�h�0ެtw+�j��雪���xZQ�Rg�F��?]�HFY�K ��u`�c'4a��%��q�U���Wй�8"Ֆ�����UXϱpmF�������Pa����E �K��%�
��@���r�(D�v�;z�Y)���&�9�MG�+2>/�n'f��xL,s�(�1tr�,�W����{���Bf�5��S��.����gPs�
�˾c-���󳤙�LPL���&�	��T�!%�+AI��J��l��m�`�ߠ��2�7�\}�=�N��1�(l��XT��:���h$6�d(}���:�{��R�55��Is�t+#گ;8}��?t'�j�	!..��b� ��M\<�\m]��l�`�Cm�	h���)t$��}�WY�)@���9.�[��8`�\ξuîϴ��b�8!��=T�v�G��S�X���wR�q�]��?]��!�����)7���}n��U�K�Dj
���w*E�]�Y���{q�
�F�	�몡�+Z���x.�E%�΍P�J-zV��dR�f�Q�_R��0p�p|V���
�r�"�K���ig���@��	�Bp>�]�.8V�������7h��v*�O���c�'͋$�+���';	z%��������"�cRG�(��z�h�rFz'�E֛�� ��y9�2'ei0�Ņ�`{# a�}wU2�&�>Y����gX��\?4g����� lgJ����k^�����L&BO��M>�j���m�S9�w�Up�h����숸2�D	ƞ��1����`���~����`"(S$�vW3�T'R��FU?rw����X�7Z|@Kc㓞�p�Ǜ�HF��c��)� ْ !4�NpX����q��e�پ����Ń���I�21����y�ऒ������y䅷�a�*2�cw~���	Y����^�z�[�	��M����f�V �(<.X�� �h"��Lm镖&�l6��ڟ�ܠ�8�XL�ꪧO�b^�r�d��J���=�Z6�_��,�4�Z��y;��<ǀ��u�x�1nR���l�r��$��4hȒU�
(���(��p���u�]Y}0�<��/&��0�dCM�r��Et� ���Q���\��J�>^��ӵݎ\���rZ-��^MC�!��L��nG(����
R��Ĕo=]��×��W�A���?�(Q�0�3�o��_e�Ib9;ɧ=�ֹ���w,��FUj�kɦ�(�;?/6�R����(�ɵ�Ϻ��H���X�������}�(�c}Nv�="�ęd�5͌�Q���A$I�ʈ��aac�: �3�4xF���$�E|7:�E������9��+��G�%(0Y�Vp+����ǡ����3B-��;.�7M�V��ʿ|�P^�"v�8��a��e�j.��L�r"��k�.�=�����'��ڬ�g56זp@�H���x��$a��w�;�&�h�%�i&s�t��N�H4� [Q��a��b%b�e��_�O���J'1*�����Ky�������e�k���2�Y馰&���d�.ｖ��I�/)�[B���eb�K��u�A��<+����&�K�"X�|Q�%�dR�O
E�K�q�1��
�y#��� ?@ʶ� ����ûA�I"h��>@���a�&	���j3��R�r\�Ϥ#��}z1{�)2�����?�3���n��<s,��gr��h+��_z͡�-o����Ŋu�Mh�=��f����Ph�7�q�Ӆs��d#E��ե,�Aiғ�I_}r������Й�.��*�o�2sEƑ�$����%��G4��I��3��s�^amZ��^:.�+1�c^�N�O�#�9+�z��Ld}�-z�[�&�@`��ϝ�)���/8��o6 �hl��&��j�Б�2�4��<R��:l[hp.���S8�?f�nΒ_H��ѳ��fr�~����.�Lh�O�%�MQ0Ǡ�z�(�U��c���OvO�g��7��E�	�k�m'�_�c5��Q�b�7���tc��y�;YG� d�20���N {��� ��5�~�g�BW��T<׻���|#��E?�����;N"Jm<\�
*����g�<��@��o��B@�<�=�ͥ�Er���}�����6�,��"��t�d��`7Ӌ-�>0Tt���-enEߋ������i&��I�nwq�S�Q��Kd��b�l
_D�^��S�������D��lO&A��@�}��$S>!+(��	��:T����y�T"�C��ހ	7x�-�Җ�m4��d�6z+΃��h����Y88��oD�9���@ݺ����v��W�1��Y �62;�ǧ��&L&�f�Ű�=����\X�D��>��%�����"}2�Xn���i�����i�����:4��� o�F��+V"/!�i|Y�|�h��_c�hK�a�QM��k�VN�hkO4�J�N�w��:�Q�_O�~J�?�d�;T���B��� �����Q��C��vz�i�I�ـ�ڏI�o�l�˒Ivu�n������j0WT������a�[:qO��LJ��H��ہ��	I�=%�}�#��ܜ�!���i0�8�5��}�wm�E����O3�u�"cX��֛?O�)q:4p���E�i�[��6�v-����D���f�M�6������D�2,3�?���|N�L� ����4�m�$�Լg^E���Ekn�Y}��� mFIF�x �'���U�E��}�mcΧK>�2�(��bv5������PRQ����6ڄQ=Uv�#ni�@����H]_�x{&�Sn�R�����;϶e�9uz��W�0;�Ld���H(�RF;�CF���9O�����y��g�V=ە�P�}���/�K�zp�b{��>�L�Oj$|{���5o���z����`�]rJ"�x��{��r&e(�|z�m��&�R������
�V�{���耡=s��$�!���Tu^k���iʓ�q�el��Ι��h�ɨ����=+��	�jw��'��v\���&k�i:��ҏ/!,O�O�-S.�`�Y�D���f���N��YS��J�e&���۫�c��ri5�ǡ�82���D(�������n���!��s��𤈷Sĩs7�'�XV��<�v�[���V��y��9q}�Tm�Ԑ����'�k�_�����gΔ��A��t',	?��T�8ɺ�X�9���'|�R�;�;1W͙�cw�axw��+t]��z-Aw6��8�^�� 9T_\KZ�4I�8]J�5�8K�5c�W_��p�Ӿ�8�~<�qmwj��&е|�N1��G�M��y��I^b�#N�cd�s������iU��_��a�3�1�!���6"#	��H��ɕ��-TG�8� ���Τp�x���y	`�0��w���\��%-M-�h�/FČ��L�ɤ�`@orl����b���J�I<`�z-I�M��������@�~6P@��7����:���h�p'��Т�%����_�B3G�C�]M�4��RV�X�lk`ũ�Nn�d�lJ�dr*u���Ǹ�gSS*i�*��3�\O�!��"���(ay�:��{�rW��B��״	��1"󗷔%Dr����7��#ܯf�X��h��7o�9`�48�H01�M"��֭�}��#N[����6D������6QG6�~1ĵ�50�br����Q;C��K��I��|2�k�ӢU���ҩ�`�
�l��o����𓅁n��bbK��,)�%T�'e�
&�[�d����:Ԗ�Q������������� �H��aBv�j�H�n���
�ǵ$�p��Lw<�����tC4L���T+9������L_�X��������7��d@%�W��&��e&oQg�	������e��$�����=��A��y6݅1	��E��[}7����A1ϧ��bEk�V��쵂��D�`�7,�̳�H��ZB�	�$�ձ=�Y�j~��/o�����0��\��x�>�x �rG*�����;��[���=��oŝ�~���P.��N�gB�y'[4�j6�0M������C���
�s�*S��L��QΒ�Z����.mK��ك�u\�}�^�֛�"�zLS�N\�q�e�Bm�-�&'9���Ks�k_m�2Z���ցTH�P>�KK�ԇ#���K�Y�����f��AF���� D���}��V�ϕ�آ�ZfG�}���s��O.@�쑜T:�UI��	O"i��ΆӅ���R-���[�5��*ة:x)-�N�����#b������W���ֹ�|3�LM�����sd�)�%5�s�b-֋a�xD1�e΀������� ��>z^�d�c����X|h�R,�4���ȴ��!�yE$����y��d}����:�M�J�B��2_�w`a���Z��&�#Z�#��	���,FG���8�Z
�jR��A��r�f�e�2�cu$e�?�nl����hӝ������#$����q+��{ޏ�F��Da?�� e/
1��i5�'S�ͅ����B�3�m����+��p�� �������G���b�wʇ�4X���e�MH�oR�ͩ��4�A�J����rA�)���[�lڧ-��rc�5�.�������c}�PQ=ǫ*��sh�D�~�Hr�E��5��XD���sk�#zXU��1�}x�^��8�wYN�,�����Zզ��c����:d8|˧
�g�������?�d���-�7ΎQ`>�C�;�
'��R0�������U���K@�l�a��jK,�<��/�&^�Q�+��u��y37w�9^R��@����(~� ��$�z8�!#�E_L���,be�%Ty%� �7k�e��>�G`N(����nj�9HM��G�-X��i[uIaO��v6���u�ڱ�i�c�XV�O?��2g{u+�E���~Z`B�K�u@��w�"@9"G���?"d��E����ݛ�f����ts9W~rX��c�d�Tm�"�����>��Flq���`��xF55tO3����V��]@	�=^E��ɔ�#RL�4�	~h0���P��߻��{-�~������sM�Ywu�Iw�;����1���'f�VQ༼]:� g��q��+7����2�ؑ6�`���F�K2¤�@I�8?��e7��/T�+�8Y��﷽�-*Z�'D0	��{*1�Xh�}͒���{2A�كYN�ą|�6����pyp��ٞ��2�(+I\��h��%b�[^6΁�;9é��]P�Ӂ����j���Q=�R�tk�
�8m|(^��|���d{rOۚ(y�@�,ِ�R��\N�\4�8b8���P�,��@B���2��l�LE':M�p�6��!uO����ъ�a�~aǿM*h���@���eӐ�v;wJ�Ͻ�
p7AHw������T/]R���`���bv\虯�XD%# Г�i����ϊ��'6!��~�I�
�"�ԓIщ^����-�Q�E~�psA7O�ml�����*�/	����U6���mw�ɛ ��Cf�C{�Q���c<8q�$gs��Y���gw�MF1�Z�a2Y|ĳes�ܭ�P��驽G���ƿ(�^�_ ���63n�d@S"�[�8���� �����pkq�s]�Q'62�짗��N3x���zɲPNI��8���T�Ԩ�v��IH���;4��_�=�����E\!/z�3�#q4��;��!UG�r��P�EOt|�f�(}ٛ �Ǭ �V�ri��Ptt �z	j����טX����l��B�^�{�@8�?�k0����JS���A⎻Cи6��4F���!�YBx��@4�����;`X@m�G��,W̦IL\�y}�HGQ��^��'
 Nډ$��	��X*-&�do�;��X��E]���f���n��rH�9�A� 9j�j~n�ڐ1�˿�I5X���O�K6��e[xV�z�4k@K!h?�۲�XP/�D �V�KҜ^5ע�C����m��Qs�J3�"_��o�+�����j���F�Y���/6�F����wDZ�W�:��h���po�@�b���ٙ���>:��C�&�@��g�ϩ�0��ؘM����2�}V�����'C���W�g���4��<'(H.R�B��8d�g�4rd�*����2��X�_@o�l�:=�K�w�ᤷw��C�:��V�~[P�D}�r�D���BE��s�����T&�;������c&��
w���$±�����Yf�
��ل��_��d&6�=`~Y�R m��,�jt�a4r8�ĭ���|k��.lt+�}��j�vH<@9y%3�d�CXX�x+Һ5�2�5MڨT��w�'H�쎳yВJ(��3`?[f)5�������I�k�.d�mOy�l�ɔ�ׇ+����ץg�ʖw��&�-��\�T����!՘>���Tb�R����$oa!^��8�(�o���pZ~Iu��k�-L�֦��8.*��?�?ugN^a?����6��Xؕ���Z��.���=�g#�nI}�=w�$�I���
*�S���	����`j���A�&��bT�}��]N�,��N�e;��f��Ka�)��L���W���4�C��rYf�V��m�x��"��Q�1����g-���No>�����	ב��fk,x;Nv���o�D��pEk�<�bP=�;��8��m��Uzl�_87�g$�];���λ�w#�%���da�s�8:-��tD�S�
����E�*�I�8��s�8qԼ�\�C]��"��-�ey~y|��N��/~��'e�=�Q>�\����$�B��DS�$WYq M�z ���wQ-�� P�2��	X��Z*�E#bn��k�K9�o����.�V͊�&�ig tD6���%\�uH�`cOu\�20?�C��M���@��y-@-T�u�mF�|I'9T�����p�s�կ�2��JS(=1�1�豵--j`�l�����is������N�BЃ�u'�J�b�����j]`J���MY3v�]�πB�+��Ma��68�q��m�|<���+Kv�����TAsB��r�'�
�br[@����W߶�dt{��ڸ�'�Ѐ� x�����ni�����\�Z�Cx 渜��0�4�@\����b���q����C�g#��\$�RE3��}�r��L���w�-h¤���8��`��oƏ` 	;{S�T�G��7��5��7�Q#J:}�g��V/�p6�H��%�8|�<�E��ћ�|��D�$�fѱ7�U8� fU}D�k�k���h���H��g�hX���	 ?�>�lז� xR�FnÉ
Rz�ؙ�L�I����@�_4<E�W�F �#����� h�'"�.���5��9	��]5�I�±�y5�"�����?��{��XՑ�yp*���d�Sc�7���]�(��Z
��u����i�C�dvh2���(1 i���]��H�3br"�)'�BB�F��Q|�]�j�lXv�z+
�Tۙ�&�
[#0y�!��k�蝧\M� �ٺ��<�����%�6)����P�G����Tf��
2����b@�s��_'�-8�i�B�9���餴���ex�$��ݚVhECg�@�xA�|C(���}oQ���t苌:��gY��,�$'�l�y=j�� �u�#,���(���⎎q�FR��\��e�oRg��K-CӳՀ�)��Z�^;`g�����T�.vIJ�I��-н��E�x>��3t����v�h���Ӛ6���Y�̧*.��&����5�o���k֦�m	��v]X�:��Ld
\;6�LE��TB�����oQ�~QǮ)�eM`�F�DXx0K--����v`�^oc�����k8��ۏ~T6n��h~��z�#����IzF��\2�g?E=9�o��@s����/_A����O��#u�5LۏF/�4VK��=�j�8.��SK�->�K3b�L�:�KH!�_ULg"�o��k~��������^\�����o�����[>ӈ���:�JpO��H�����kQu�k�(�'6ji������6�HV�t����/*O�y�9'z3��p��B�a�Z��z��}�nkC��d�\��(Hf�ɝ���	N�ޙ�m�1����'CR��-c�#��	?����ͧ�k�d�s�\O����c�-����L4�-�D�E@G�6��ܽϢ�(~��#1Uc}6�������F��1���b����r�B>I%��|�]���7���=�v<\#"ߋI��ʒ�Ղe�
�_� 8/��I�EV��6栗�L�&.��'wz�54TV~p�N�Z����J����&4����>�F�ud�I����E�c��Ү��dvϧ�[�eF��0��K�m��4ѺSÂ��'x}1�<�C����v2� @�|�q�d�V!�$��*�!,��4�Dƒ�_Z��*�1�G���L�C6�@*UyT$2�ґ��aC�p��t�i!_d���۟�n�5 l�|Wf������8ERGcd�����t@�^�<�4��,|œ�bRP��V�lg1%|��k��I~_"z�m�b[��Զ��.1��#�6��W��U.�s$ 6QV���76H�P��0,��Mq�+��p��
�
��Q�g|�P���3x����~U�w�nɧc1�w��~��s�b܃u�}SǞ��{�X�>�<WL:F^ԋo��{Ï�y�-���z�{�1���%�I%�E�����|j���u�ԏu�'W�'���.�Dd.��:\��Iu��jgx�6ʈ3T1=c�ޫ��h�s��g��T�������0�_��y�T�j����@�r����s#���Y����]qCF�vsX�@��2ۭ��žׄ���U��؅�R��v��+����g�����kD���H6G;�U�� �90_��7����w6�/w�FR���\����٢}s��}��Se�r��em&�mF�dݟ!�B�|�'WV;(�,�`gOX�{I#�dܝS��e����좵�y(��̃�Q���y�J/��M-�b#��2��J�����V2�r��B�a[
`�(H�P��5CFH�7��O�^�Q��A�`��˯s�"Kb���a����'	��g)ɶ�U"}�᪴:�'���.!�M�%�JI�0�2<a�|�b&K����ng
�sIB�X���}ˀ'�N�y�������.��MO�2�S�k��P(�wj�u�.�9t`�9@���S��b��� $���������U���TuD6������Y o�	A���4��!\;�M&��4�%��46a!<vy�U�@�r��ɈuIQ_6l�\ф��wz�2�\cW��1��ʯ>ң�	WC
^�ǰ�����l��y*�J2�A�����u��>�����͹�tw�ɩa�2�n�(�%�+�ຳ�ׂY��*���r���q����՘�?��=��uU�4��D�B����Yr�'��]+��뢐�X����M���Sզ�/�f�w(��ϼ��$��q@Q�٧���kX�39��d3��&1:�L�W�S����GJ�N�d$m�+��&|LM������	-\��i�q����H-���%WơHRC�^iƌ�Q�{T)��OL�<�|��;Qn\F4#��ߗ�byAM�E݅�OW�R	B�![����g�-�>��yE���:<:;�m�x��ז�W�+��>VI�w[�Ϗ�>�$����}�k�T�V��d�rU��U_���$_zתʣa�L�i꺾$���>c���z!�h���Z!�9�}���������51Stt�䵧��S؜%��	jH2k���U��q;RH�F�v%t/�W�uG�D5��B� �Sـd:9�=�C���;��-�b6
�����fM_N�IT�0U�ެ����B<#�ї@,%��.��90J�F�������y��JeD����y�g�=Z7KzY�yr�0�@8����_�28x>����/��q}�������eJ��8s�?Ą���U46�Ft?A�W��'�U������Gմ�4�	������gw���a���h��Z3G(�8G���:��U٩�v���XZgq��ƴ)�l:e^���.�kq	 ����UQ��[�avs��U!2(ot"Fw���`�1�v���=�K�i�L���ޑ�fRGJ�J�I��3�3P���J�f�-��&��Me>�z��E��E&���2��u���ɉ*�Eݾh��~�
����������G��(��Io�D0�8�y ��&���z~�06�<UA<�f�U��©?�����@��e	���a���BpR#����E<�5�;��a!^���J�"��#��@�
����j27ǩ�\#��ɡ�|������ҵֽ��aʐL	�m(:��	(٠l@F_K�f���o�s<	W5th��J���������m��Y����;��CUߚV-��>��r9<=��'�f�\����]ĸ�ڲ5\�����M����{�-�0Q���xW���Љ�nd�&�s�1��9�n(��़�"��r���PA�L>Г�,{�?�I�0u����� 	1B�r�e�ȩ5:E���I�&�ě�H������^��V��1�����%ž�1PN�lH����O�;��(��E�]�>*֣�߫c��7_�.��όV�`���|��Q��D�1h�D���q� ��H�NPo�������8��;�14�a��
�g)�H�f�cF�آ�K9YW�N΀�2m;�ht٥�K�ʼ '�S�G�c�g���⭞bM�o�.����轋���k������ɲ^��:жX�X��t}z�^��ӱ�Ū�#(R3aw��Ч�Ռ�b[��z�6������b+�Q��ٻ�FK�>c���}2�ɝݎ�����c�K��Y��(l	[\�����+�����0�Δr��`,5�!�P	����g����eFD��q���{�_�&����@��.F��ye�P�l���s�u�0��{ÑaZ	O��`����"��خZ�ܰ�;rT�Y9��x��ض��ܤ��预�V��M�u�䚴G��AIL��F2"%��Vl�/����I�:=��0��r	��Z��D�Z��u#����I�Ȍ�Xv!�s��[����"�C���&���8<�K�6)�D=h��4�!��l-��J�e��%���k^�����}3m�4 �ȳ��ôF3Z��}$������p�w�Z8xM�s�z���@���[� =�a��KSBRem3$t�~Ȇ�D1T��\h�'��DJ��C����j��=2����J�Pu��t��wM�Dw%��ȫ"��-�C"�aB{y�#T��2�2��w�MMh�8�(r[Fu�'� NG�Q�a��&��i��O��b�)�Q+��whb����3���L��ƕ:Z�WRd���X͑�AO��/���6�BP�v���Ȋ�F�2�W^ͤz����56�S�E�Yd�:�!�0�����U���z��/����f�I�jx/�yx�0�U�8�������Ap[i�)W�t�w���1��#ڼ��&6�4r����}�a퍼Xp��oS4�?y)�n������1� �K�IA��8�������t%f{v��̙�r����ej+CY"���S�O��P�-c�B�J�?���Ĉtg�<l�;�Bz2���@D�n�s.v���-PAy/8
�3���F�&8��J��G��� Y���^����t����]m�����o%QD�m��2���@�	�J�9vTW�f��)j+� �M� 7��Ç6��"����&�������=�"�iS�l�3Q9cDd�"�h��۔I��f=�����P���Q�X�4O"�`���m��A���Jykx��ωܜ�R����JKd�Cܧ?^}ق@�T���=��t��%Z G��ӝ`�-#ত��+Sq2��ӨP���J*��x&��Ǚo��M�vI!�W��Ć�=S[2+;�(��T�D�BV����T#���6���0����m'�����ۓlwUiȑ�����G0	�qr��zgYy��S��mW�Ok$��,9Y&�#��9���^�����8��	a��Z��!����><U<f�p�����6����B���΁�C%�RR��w���W	�}��=�M7
��D�Gb�6VM�|�Z��*�H7�H�8�Y����@[���у$�"�UZ��[�{2.ϸy��|cL L��lҮ�N�z�f��߂�X�3[��	�� �S#����=�P��]�@8�����A��:��q�`�ϐh�,��xMs�Oy�����((�>�b�|��B@��w�j����6�|��Zfl��6{��'�?��q	٦�˶ך�`�>632$�r,si<vp��ӂ�Pb8�dh�V'\q�%Ji���p��bСˈ�*(����R��z�b��?��) �B���1e�ع��rP��B_PK4;��vo�z�s��H�p���b4�3'P���'���.����hX׭�?9n��,�`�䍢����ݑ�������-�i�8��q*�}�bɽ��l���v�n�p��Bx6_Z�.��wдBd���Sos�-@��c��3j/zٙ[{��p�5�M5D� �a�g�Z	l#��(��-���¬!�m���b.¡|X=pǰXn�~Ws���g1�3�»0�B���8H0��ݍ���p�0e3(�u8ĸ�'q�͟��H���Q��t��l���c8WA�5f�18	H�p����=�������X���Zr:qqx�: �_�8L�����i5���R�e��F6��o�#�p�ky�f��/�V�'�j���C|E�okg���?"d��̯5D�!n���5�(2hh
��܅ ���t���#��)�uU�sF����%@=�#Xp��v�9����"�