��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#���������l��U�~�׏O����j9�PY���`T���x���s����uí������P��"��b%>�1eτy�<�gܰ�N�Y�	� {��I�ɍL�ݫ�G�R�k��Q�!E	�5E��.��:�͂2��y�m�-�.E��i�����YS�
��@�H�ۼ��nD��Y�l"BU�.TԊ�=�-�����q���Ǹ��j��ԋ����tr�a�ٵ�]�b	��%�ɔe�)rYOjX5;V��R�������M\�	D��ҏ����9c=�Vͼu��Ro�P�Jf�tRvsY��c�"n�XO��	3g���Q���^�Bʹ�7gQ+Г���$�-��t�8�����A���<����l-��*�|d���V��*<�G7.�cm��YX�*_/���-��e?5��>HD����O�z��`���;$����:�}�wz��y G!r6�sǬ���8��b�����<�uh�:����T���S��?�[��/X����F��*�� +�#��,S�+�Y�]L(�u+*���$�a�)o�x����zo��9f���5cE�ѿ�C�N��V/�|��*~�^Gt�'� P�_:41�t�?w��P�)m*�n*�L���\��_�8d������U�����o�~��'ۘM�wH���4]�+�ބ���?��ҐƦ@�4�pӿ���sX�����X#��a�3	�^VF �O2��ƙ��]�1�Wy� �l�cwm�g}Na\ ���ɛ�q�z�0a�v(�>U��)c��^�[$�����Y�:�Ԕ]ع�Iv�G1�����+
���^�Y$�b�ڢ�4��X�i���b�#��m�����}�w�@��憎&7�M�x̎�?S�`ߓ����D��q��`{f�2���3�k+��'���1�'��I�9�nc���._�A�?�#�Z�M$Ƞ`�V.$���z�*��A�E+ZZ�J�̜8�}�_�T��Uӷ9D�]�X����� >�94l����R��3KP��I�{&`K���X-�<�-�(n�,`<���2`>`�@3��X��ZD8/',������t͓����i�(��}x��L���pg�*��&�6
}�Ү�O���%�6���n��^����34w�c�:��ua�L���-p}���f㢧�q���ۅ�4z$���d�g�&u��� h(�]�t����!0� _
��J:��p*8�ѻʊB�"�SV�T�6���M����R��Lb!��D���D���X1��/��/��s*�+wz�5�8,k����V���5�G#���(a�����0E;��{S��O&� }���	!ꎍOP�lZj~���tk����3��vq�2�N���:�h ���u��+f��k`Q���`$��~fct!��������7m#��U�TZ���/�P#��ݼMsvZ(���.bެuQ�O*ݮO�H���x����%��A:w��m�>��^2͇���N��ZDʯ���M}�?�s��p2t�|�Bu���1��W�Jo-hS�$SwY:�aް���?[;�t^��wJ8���R�x�)�����P���@�n�!Cd��Kt���=E1u��ۨ�Aũ��S�K����t@<{��]\�Tۂ5�t���Ϫm�J�B5��/]&�T��`Î\�br�vv�pO���H`
�z���A$�z�fUp%�
�����A�n������2��� ]˕d������b�a��μ�2�cR��hb��7����U�)#�µ���-F�c]k���-� ��ۇ��`���ڰ��t*z�M�!y&9�C��B�zP]Jrv�.J�]��
�V�A��3��b�0�=yR_6��mB�2(q��!�c�p��}�Ǥv;�K ��d<����YoR�H3I��r�.�scq\Q9,e�B�M�۪'�}��i��3�u�7�|�)�c-�m)�����h����J�+�U����c��$�_~P�u����'�g���	O��s���v�]�����+���rm'�%�"���&�);l�9� ��Ϡ�[�V��x����C�%�&�ߜ
���̧k�Ne���������	�W��
O_i�Õ���b:'��U	2q�������u��N�H�1O�.��%Q�ֳ4�7��;HӋ�4-瞧�v;����/<�3���$��Χ���G�=���To�gf4ds�9��y^��u��Ы�a��S����R�%���-��<��3=׍���y[,7�1̹kvn�����h	��h����u4�T�������B���R�-bE��ڜ�[m�DbBV��6}����ý��	���c���Kr���\E���j}�J�z!�Z��ïh ��7e�b%�hi��a}Oh�h��z��1`#�)
�Yw��������x�i�;���d�\ f��	�wo�FlLu#&�!,d~nFօ6t��v��6�+HJ��WUg%7o|w0�@��0U=Р�(�"��n4��L����^j&p��e�m'ȓV���i'�M{�$��"߯��TO��;�9�N��8�	P! ��� ֗�}�ϵ|QZ4V�r������F��+Y ��[�J ���`5���0���v���,Emg!x˘-��Q�Ul>
"#xRp=��¤)؄���zP�ф� �t]������j�����]g��$=)�Ɂ�vF!ս�f�lc��>���x u�-8�G:M���?^r�\�q9W�j��}�n�2:�IU��.鶓Ü}8]���zļ&&Q���C�^���jȓ�/�ǻ���r�]~�FQ~�h��;[Z����J+R���b\�����=�F���d�%���|i�>��#府uo�jd8#������=�2I6�ٵ��>}�5G�h��e{vHVN`q�W.�ͻ�kz[(�C%�u@L4�>��o��.���]>Y��N��w�|���}b� v»w�֛��_��H�x��/�/GC��#��ĥ |�\���Q��{�>�r:)*�����M\�:��-˝�L�ޙ�F	/�ƽ�����lM�������
�$��������U{��I�A�<n���1_7Al�,"��a��f��݂(}������ ���C���0��k��E�*���`�7��(J�Mm:�f`�:$��B{��E9"�极�kd \�z�R��CNL͓��Y"&�|k{���uJX�}�H��,m�̣��hڃ8 ~Z"M�z����D�JBo������x�Ya���#97�U˻���!�V����-�����aZ��R�H���O�����y#���7�c%3�D�\$������iS�l>��c��"[�%��nGJ����C���?���c��o��Q���b\�}��dl����$�ŖӔE�V�iNNp �h���⽐l��ӅRseڲ�E��J��ю�&�ӫliЏA�0-���-s��X؅)���oj����-P��^���ۭ�7,�K�*��+i����#'�y K˜r�Q�bE��A��0#��H���snTx�ڠr/����E�ɃQ�nH��ɍ�cy�lP���OA�ϥ�v{�`}tO��v�ܸ� ��x�0|SA�簪BL�C���C�[s9W,2�#H�I�s��mk�=��[X%5b�iQ�/e�~�z��M�lה~��ep��c�׆������e��G��{68A�cPU��nJ���h;c�q�)���_�+��Q.Dj�9�.��Q����Qwr3�.�Nu]�	���(�،zKU�1j.xϮ9����Y���eY�7�~���zY�{�k�ᬳn�����e�J���D+O)%��s��UT�N�؟�큅7L
t�*��o�U�nd3� b+S�|�d�^tv��>y�����w�6�|@ޠ��X�D���R�E��L��v� �O ��Q���&^Sj+M@0k��J�[ �_u��U�n�C��39 jcZ7�u�mQVPОH��8����K!�;�7^�@;^I�������7
W�W��!"����B�\#}�)O�%3�j>����rY����9	�@�4S<�+,���Y'�(^y�T������)��s�~j�RW��:d��TZ%>�Z���K��&#^n�P`�9fb����_X8�?�9� �]�o��_�����s�������ˇ��<ys������Ñau>x����C�������n+�c�(�kKw����5��zzm����+j��ъ2D�h�O�	�8�DԔPh�Ib^�3�ǵ�3�\]�:�h4\͸�����	�f�'���W,��j�WS�Ǽ7�xٻD|#��)����-q�I��w�ʵ*^ğ�*]��,QW���<�sy��w̕���;��J�?�#�u@���^�$Iĝ,T�Q��9��۫�sǾk������wD'}��_2��W��[̻�e����P�n�zv	j���C�U�.N�"O�Z[��Gͱ��J��A�G9\>�o���zB%]��h�\��$C�}�T�T��G�k̬Íd�\�-�R.OY���mm�O}���T)m�<��sO���%�����{����-��4Ƀ����\��-q�s�\�dH<R)*�w��h����K��0�U�[-}�Ϟ�a�v(!l℉���k�}#7��!D�D�͉9���D�����>4M���J�#�2{t��~���4�2Kc&h�����FUP��m�	Ģ5��lI��]iv�ų �����h����K4��U^jc3�EBuw����J���E�4"���l�AhrA8���H2�]��v�Q����,�;1�dH�m��
�h|T�GU��X!3�]�e�h�����$yY��ս�ݑ�a8H4�
�l��oEG�_��$iُs�j�=�?c�7\hD�zbxk_4Q�rd�=��g"��;�������=�)
D���	)��Jw�)Ɨ6����JS�G�2/��ST���T��7��xJ�1�<󣬍q�T�9�(,���s�1�'�Q6g��E�M�����Q�`yn����rO3��+�N\��[����P��>�+8��6���1q&��v|�f�(��NMg�I��@���s5�ƞ�</�+�X��&6Ƽ1�i~�}Sf&;�ǶA���)�R]w���.�p L��R�ƺJ�N�۫j�OLnַ� =tD�,�`ǈ�Z�`��6d�����¿��6V��
�?�Yl�%��:� �OF3�!3Za�5t�"a%�����>Y�1��
�=Ȇ�b|*�7,<��%6c}��>-QcsQ�낮��F�'��&��t�nT���Iy��`�i�iX�[h�s�#? �U�)v�m��p���[e{�W�5vш#g���\4�v�~;��I�v�@7C�D�H0�>n�!(��������An'��ǟ.Q Q���V�<��7
��:۰˜��d�&�H��^ SnS �5�����-̀������-�,�6;qm�V�5|��p����{\��P%3�^Q-3_=�]3�d�u�1	e=�},$�og�GƤ$0�P3q~=�����g�P ��L<x�5.�)�!�C� �v*YR�ד}N��\9`�x�-13�I�g�&�w��SmH� e_5:f�� �o�l&0U��.B5�j�+�H$,ʲ���Ѧ�5�6�Qa!5��p(�c�?�j��P�>nM��]i�����%��N��~3��P���w��N2�#瘰���Pw�,��k�
�L#gC�Ix�"��Պ:䪶�+��t�pD�p��@�:?"Z
��<�m�\}�:C���g6�����U�:;�gw&޳�O�[d�������x-���X��U�z���Y�c��0���k�;.C]�����v���,���f �sn>)��B۵�5@hIC����%��%����0���5bT�`l9h�
�.]MY��$y����Yց��+�����Bm���m�q`$Vֹ�9' n�e��<��>��Q#p��.��;_a)����Yb�턙�څ�m'�拗�~O���n��B(+���%�g�x%?yȦ������3��n^La�?�	P���=��a��Rod�o�v��%Հr1�I��k̫�L��jC�ٿ֋I�0����t='�7�p�7�X��Z��5�0/t��)��-�X�}Q�����M,x�~�ϡA:�:�Vފ��b4J5]��73����g������kwm���Q����cxp��?8���5��g�(�r���?�y�S��.��~�&�X������Z��O''l[Us҆h@8�����á���	3�;xT�Q���nc��Zd���ٞ�ȍ�q�B�^�Ћ�!��Њ58���܏���K&|k�f��ʤHA�[q#�#�T��r=��GB����yT�J�����B"s�7+��ԟ�ek�sk���@�q��w׍ʙ.@AD��2�@db�E�r�6LSo���.�K�$��*|�Fr��_����c�%e�b1!�>%��m4�Z�����B�@�/�w��&��yR���~j��Iz�I����s�l	��bH��Mq�S����ߌ��z���,�ӊ+QS�`�~�I(V�j$e�����G-�t����w�Y��1�m�:�0������2!�ڮ���K���[�:Q�7�T=[�W�dw�x�U�A�N'$D�,�+pc{0S��A�������?^%w�d`��[�l�ʒ�⧀�{.1$EKcn���|����L__��{���*����cܫ�F�h1�d��R��L�`²I@)��z������i �47��"HD�I�\��޼��[�F�
�~�X�U͍��B6���Y�n�����I�-O�k��5Ktw�6��G0�4�O��V����s<�r~��q�a�Ha�6�èn}u�����p����b�O�"f�(-i��Z�%�{ �qZo���N�M���g!��D�? g����o'��.B� ���3��H�Pf�\W>��9��kӉS͐�n�(	�``�4�8�~�nA�G?�2s�n��H\�Hљ��������WR��R��"]��a,��΅1�	Y�}��L�TŅ�F�4n3�����_H*'/�5CS� a�	������B�wl����3�K�G�����]␦�.�3 
���Y�z6��݊�` ��N�����m�Z��Z"f;��`}eeu�.*��BW9�俒�������z0ր� ��*;��)ivz���\��Hg&���|�3f�$.��a�k�YY���
����a)X���= :���f�?o�XI�{�Z��b�p�G7�a�$.#lQ�#��Ӽhb��ҏwCD�����U��K��U�]���s���08�֨on7�]Ĭww�촀��"�����e��tzĈ�	����eR��F�Ƞ��!��B|�=TRRz��=5�����Nu��s/{�3+�ԓEϷ�tvT���g���d�t͜g;�lĻL=-��eFR�]�W�H�~�2H���E��<p?�E8tX���L�6뤠��C ��BZ�x(h���F���f��N~O��ݸ��M{�F�6'3wp�s��'���sy�G��m����t�$
D��K8�������<�+r9�7%���ˋf�}�TzT���*������Kqf��77�hb�:��D��d��՛�[�H�(�-�*�pŶ����4�#�2�	��� ��Ay�P�t�2��& ��n�i���LSO�utg�D⨪�F�h2n3.ַ��_X���=�ܺ�bB9�D)5�:+�㛉�_
�}c��1v��;�Ѫp6>�f��]g�ZC�4��H���'�["j
�a{QF��+�O��章��R��+�$)q���l�U����||���Wǐ�<X��*'�ߊg�1{;B+C��8G��"�W�tް��/��z&d����ϙ�7��5���Q&<߻��vH�Z����I=�4�8ϛ�Zۣh��f(������f˳�2�ϲ� [ۖ[dT�Zz7*q����Sӓ���v�>�V'���x)�JꨒMS+n�V��`�{��W�51ZQYN,e����x�H�N�yA�>h1k���QE�h%�¤zD�X���N:헾�=�os�-5��b�,��F�$O����SEd �Y?*K�F�}�0ak�������?�97�����'���0��7�8�w�m�SiZ,Ĵ�.�y�����9�Ϯ��&����E�׈�Gj����n�v�s'�v�����vy��`M���ޅJ���S/��X�o�
���V#.؇S+Jx~�_�&�:cJ� K�o p�����v{;o�R����o��bG8���意ؑ�{r�ɭd?�ֈ=���l�hP.z��s�	��eEe>�M�L� ���r ޣ�V#�� ���
��4���o��^ï��94Oa��igs�kS��K�N��~�C���	M��2�]2]�jv�e�`vd��D+uJh��/����'��E"�hP�N]ֺ�����W�"���/h�Y��E�i�]���pJ�s�9�0��¡��SK5��@��o�݊|y��ZA�)��:h��GV�N�ws���u�qeJ��v��y�`��Lh�4Z�a�p��y����Η�C��������xR����ȣa��7�_�����f,��}����FD{�(�e�?4�9�πP���5�e��\��W�¹����`u͹��0F�
'˹����ה1��S����g�y��?���)uƧύ&gc9pg�����q{�����y�z�Ěy�|tr���Yc�^-�i���Ka]������2��0��,�gw�����������S*C�/>B�_*��%x����S��q_�
�sL'D�۰��c=�Z�hWX��ή��?�1j�;k���.:K4+�Y �arX��a������L��kD�E����4\G�h��q�U-d�+Z̽�! b��/�{�
���Sm��]A<}�C��ԤHʹ��juX�䂢\�u�� ��RN{l咞O8iD��"��XYt�I��qş�4� ��N�cu��s�o#G�,��T�z��eq���`t>}+��6��3j���֙����۬,U{:/�SXхk�k��@ks��eꎆf'a�H��v}f���
f��p`ϰcXj�)�r�ks��r�`˝F��ʐ-���Hp��VB���5WV�F���r��Ef�^���rH�Q�=��t��1��A.�l�]I�Y�z�GR�O,ǝ(��3&8��OP���k��| �a�!�&�U��q����m�%�dBF�Yh�#��2���f����u\�h|k��z>z��]+#���X9-�����x�u�|hnOa8���e��ƫ�?�N�`l6����7^w_9���J��Aթ�V?���%�V�&8 30~�;�s��,x�}�a��p��5���=��827'Qi�/�b������Yi*�gB�~ޕr�]~�����+�[�Kt�jN���|���O5�A�1P��`�Mޠ���F���x�r�&w��ԕ5���O�4�c��������	݈�@1��&���dqLyxr� 9��N0�����m5�^���M�#���4|��1�!�[����
�6L�W����pJ#��w#�W�B ���[Q�b+��WB~5��feVއ�i7��ڪ�i��hȻV���{�������u�6d�]�u[j�ث�j�>������?D:�?"��]]d/˦�E�Z��ɛ��"#f��!#��&������K�v���ά�|�>��y[�O�������`*�Z�\�:%VH���� ;�Gxu`)� ��)%�E�d�`��y����;Έ�vn}���#x@w��󇶞�h���ֶ;x<	�W��$�����J�C)�j�m��Ōt�XC���Ͻ�>#������D8�LG&Ңy��#9e�#�5r�g/�
�T��eJUî��|u��}$Z�.L�4�$gWh�Ǚyw��53��M���â�n�R�H�u<���)r�9���э�n|��qR�ɲ�ɐy�v�b[�;�܁�Ö���ǜ�I�A�0�'�����|�}�y�'�Qlo���*���W�p��`��Q���:C�#])��!�;�a��$�������`�'��Ɓ���j�[~.f+|���Ϫ�C���t��y���qGK�.����lf>��쎥h���L�L���J<�2n�!֨p2��L��5�r�O�A�VI�Fd��D	���o*� ���!j7����q(oNM��9�7]\��z��@�r^4�ѻ�����$HJ)���y��ڎC:��)�)����L-�N�J��n�J��x��ZJ��^��@Р')&򔝩��S0�;��Ry�h�Q��Z����L��V�;�=�~���G ��,~&��?����Y_����L&!>�]bWH����EX�۔���@��Ս�Ƥ!e?��}�V��C��kZ�#2��㗊QX���t�
�T:�q\5W6Ө��֕b�l���G�O�>i<�CP:q-3�
K����r*����/7�N�HH�� ���jJF������x����X�|��T�[����~�1���\2�����м���gj����N�ǈ��f0'�׵5���]�)�hfQ:��j�?���dm�cY�g�����$�'��PQ6x��y��\S����� �R *
큪g��"��d��/��(��y[*7#��£�_��|��z��+�����j���޿{��8��5̣������Ȋ�\�0���������Jxy@Fu����LV�ǹ\��C����l���K^�O�Hm�4C�M5�Lk�ȍ/${���Cx��5 ���eK�U���Rl@:�L9(/S�ק��]�Lz��[K��M�
r��O��&(��+Q�p`�����Nڭ2��_*f�(Bv���؉�U�Z�gަ�G['�e�"m9�g�.��9m��+lR�
��S�E��¯�&�ީ��K�����/Dl_��SZ�ޙ9�H�K~��\�(ӫ֧(���d�'It���)�Tw[~��`�<1�+���V��y�Q/.�&�$R��?2y(����$�(����n���F��s�s{��qw��C�`�4��G��M�_ZI�E����f7-j�塅 _�B�d��fL�iÄ��'YR����xtC����OZo���U�C�'dBg�P;�H
����C�ڠ����A
��K��D�55�d�n��R�א�az���7�?/���k�������'<�)ʩ�ފ�ƺ��-
��	��v����+�ꏠ��X>�����D������;�Bo\�^�_��A�5�,�&]���"�6���1������L�yW��E@�-	�¨2%v��i��\-'�"/m��B�$1����ϱ���qI�ﰉN�����ɡ"�1.*��m�-3�_a�ٺ� ̏�ū<�LR���p����R���3P{�hum����.��:9�&����$��#ݰ�"]�������-U�{;�t($Q�Do�.Hb?n��p���/� �3&VEKv�t���B�#�*w|� @��#
U�vnZ2|/�C�I4��x��L�v!P#f�������M֯�#����W;�es�4��tl�,1��(���;��"�5�0׹?��a	`�$V�Mڹl\�r��g�MV�@�u��1ֲ��g)-)3�O�N�rL|#�Y�(���ξ��-~a���Q��`_t>��ʺ��B���ْ�Gj��O�x�7�p�N��oˡW��/�1����F��7����s�
GFn��V��y�:V+���>��:>�m���B�Bj��
�= )����ԶڨE��[�[������A'WR�X�S���h�bC��r��ξ3{ͧ�⺳���Wd�yId��*_�
7��]�$�����J�c�O���������LDG��MT�iC������\pbd�h���ݏC_��������݁c�x#LA��ĥ�ȫt��"C�s��7�?�����:�����=��fX��#�k�\��f�!�={�,��1P[��?����?�z���?hu��v��Za`.ޡ|�uQ׳��	i'�9��6U�DY�v�"�f������;��"�tZK]~�0
�O�A�i��ӥ�Mjt5q�B�cnmst��&����JNm�l�=/l+̿�zf� ��@�!?d釆�[����(B<L�M���������*��ߧ�)/Qq�
���@��Ǯ͒�����ϟ§K�m?eg�s3��M�%A4��d�N�l*|���3��>�e��z�^T���/!P+���1'�m����	� �+��UA�� Hr�=o��{��`{>�욯�K�`ݪj-�♡��<�oH
B1�t�E����P}p�L��b�
��go��f�ēPL����?ZEab�kȥ&���|��_v��e�X�f�Sϳ\����D�pޭ`�έ/�$z_��R� *A���A6L�a��[��L���(�Sѩ�jӘ\�
�	����O�'_��Ņ�x锏���^�(�M��ɸ9�[���r�h��4�}Ӑ�vB�0�v-#�� ^*�/P-y�3�wG���`'Zd���RF� � y�)h#���?����<oY�a�B;#�\>�\r顬#nA]2_K�nVe��N�Ԥ���a3�`L��ck~/i��/	��dO]�2�A/=m�:M6k�XF z�զA�����}���b�h�~g,��ed�4�]��{L������)X>�9����q�d�W �M-�������g��>��]z�h��{��n>��/6M�����SH�|�k�3��W��ւ�X��O_�s���B��ꊙ�ZD7������z�*�4��d���MO��h��fлK��Έ㜠x,�W�	,J���J�Pf�&�qǉ�hD���	����8!pc6��˰k5��Ɂ���u��-X_�;c՟��DM��S8ا
{�j G��':Hw�5��}$`֕�D�BR��qv n݂�n�g�+�8a�0*���{��c7�`�U@�u�Ά�"�{<&R�PZ�2�(Ӟ}-�a2"���Fj�-��D`.I��n��` ��R��.ұ*�i�R�
7܆'zj�>m��d�.aY_N}�Y�"㸐�$��5�]L�I�a���5�bl�)csӝ�s#�*g?;Cw������4Z���;�5]"d�ԍ���P�W:2��1�a��ۈ��ʢZ�Ma�M]�}9�Q�m�!.�qh�� :�L���W¯�Qh�2�r'����W�6_,�P��(�O�X��.�ag��L�﫻|6f�d{5(,y��>���yx�\��Ы�?ҋ�؞Е����T�H l46k0a�~[�,��X���Ov���*3���+�WlH���������	�Χ��^-�ǖ��!�C�w���b��3v�r,�8�_MG�8}]�7c�����}�8�5W�:����8�h,����9\n��µ礗�@�ƭp�i�O��IcX�i��-���Z��-�������o��z{��0ϡ#	|�kӅH�����
���@v����J������~M4�oR�bi:�*�V�՛�K�<��Y}+,U���ɓ�[����$�Gɳ���ui�YRM&��qRD���O-3P)����6A/��d0O��W)�bj�����A��uڦ�����[�o{̅HZaC��$�-�G��)#Ň=��ϻ����@��a="@�[Er����+EUgض=�ZH<�9E�%��;����Z���i��O�=C��sFO�:�¢F9��Y�AN`�-#�KQ��gNi}�"�4zӀ�[��6��D�K�'�T���cR�R!NC���]�#y�u�35�,���UW�3$�M�h�����者�oj��0u������GkL��?�ѐ��M2�P��n ]���Jc"�M�6�Q��f�	�h�9�{�_5����P�!q�N���o�����,|��d��+�G������|���k����f�W�D>�`}{2ć�B��?�����k���ZG/�n`)TVC��&����x!�Q��W�:>`ބ�	��kz/��p�c��U�_�u�vT��9�|�F�N�b���fJ%k'	n#>O�3�D��_���z>��g���i�)�81� �>\32�?0;R�-���h�K���V�j�q�Q}+��|�b�啙���>Iʡ�U�s��a� ��3b^�U�<�&~����+O�{�dN�R*�M���>@+ac��·��(��'���z��?Tk�Y,��� ���g�&.ȪBF�1��i��������"��ܝ���y7�N��=�]�W��^&�8s�tk�-!$����ss�*n�������|�m�p�2�zl��ɫn&�F��I�6��(ظ�2g������e��0�3�-�eh�G�������p��s6�&��~���bp�j��[_�
��%���3D���l5o�}:$��57��$T�)v��iO��������}U�_B�0A�r�����&�g1�6Q�Ճ�,��j���Ů��X-�*�A+���G�m�4���U����e�l�bϓp(*~/k]g���z�ǻ`\�%ӟ6�Y_e�7�V�f}3�o�!�2� �j��5X���RP�G�v-&&��pT<6��q.�Ww�
� \f��┺���P*�p�ɮ��W�G�q��$�цc-&Q���+��+��|�:�����{EZe�(�����o�^Ƶ?t7��M�̩��	�[�=!�`��翐a�K��������J�7|����Z��ſs����6	�쵮I����HѰ��{Y�1�V�!a��<���֞\1��E� Û~�U12��9��Kg�9� *�8_��M��%��9q�àn �a���mR�&!*���l�"��o�����L+/��7:�Ր�:���!O_���nN�/0"@^���x]鞠;�C�[�(�u�!t<c��Ƃ��.J5	���aP�����\AJ��p�x~UtjH D���^�����Ҧ#�|p4��L���v���q��R���E�<��?֪�ύ�D�����|��H�O�7�jG
���} ����gB��Q�Y�d�3m��.7��2]�Y�z5�	w|��;�c����ň�mj����������)�"P�׬E�E?C�ܨ�Ѐ���2��y��z!�;c�̖��|�棊TP�MZ�E�o�G�"�t�*���x�ǻ�	О��������S���B�����I���أ9tFJyi��V���U���x���+Z0b�˚��j��O��^k됙�=K
ȗ}�e�&	Iap����{��Αg;s]��j�z�����<���)n�����m��p��q*��$]�Y��s�q� B��N�I�s\sE_o�|'��W�ћ��7Y5M�	Pxz������|�lS������^{J㭼�'n4Qc��H��BSt+9��P��a�x̈́}Vؔ�xn;���Mm �A�h��YNR�C�u^��磼���5�����[^���
�01]��.nC�o�Pu����4rw���pǄW(�s�ō,6( �ɨ�N8�<��Wg�u72��o�gFLd��($���[3;ee\ �O���T���n�fךW%�}@T�r ��` ��r��J�����@��Vx���Zs8��FL
�t�l�k��s&-ǻS�~�<���(� �7��̼�:���m�Ч��
��_��QA����K�i��VN��n����Y�8��|ԾHԘ��d�@�]m����M*���ޛN�%�����ӌ4 #G�0�C,���<�]$��e8��>��ϣ�=;�e6��Ɂ�@6�V��l��3.�-F휉�iv�~l�ܽ
`H�f�m{Sl�w����k+���)�"�c��wH����L]��EZ���׽g-�8H��	�۽������̈��\g�cb#��3g��P[�т�N��w�'#uЇ�6����@C3��֨d�?N�]��-T��yL�R[�����[�i��&������Ю���n@@"\Z	 �y3�����Z���RFW���#��CFBJ0N{���T�y3��־������#�����k�@U&��蓞njt^®������|z38@m�Z��!v��sg1���D��"B:r��#x���~�L��f��ꌓ�jhV
Q�GP��m}J9߲�з=��X��f���p<�&�Z�!�o�������k����и�����E�Hb�{����d��ɓG��D2�Gc��#*���3O�]����!l��K��_(Z�1�k���u:���|U��'S����ƳC����H�׆�Ħ�.6Ɂ9��� ,/���jd�q�␮;��D,�!��5��T���kG����?CT	=�
E$F����X�T�*7�Z@�ݥ�(�p��pR{�|e+�r9�e���w9Z4;W�h�X Q=�`#�-lQ�ui0��1�}�OgRb*]���i���ٚ������KO�>�E�oԖ�J"@�����a�\���k���ԅ�~|n�˻�cJG���c��*���#��8L+���&��9��@�t3�e3�r^��S�M�1o~��
z��o�=_r�Z�ٗ��I�s{��럙�4iٳ��{Q��ψ[��M�g�gJ��m�����H'��5ɺ�Έ٦L�֡��lr��v`��:�=4����)��{�R͋/�:�~�O��\$���	6$�R�n��i*�@o�S���Sd�a.p�#w�@����{gcCY�/Y��vϡj��J��]D���tLե
���4�(���}C����fr��Í&6)6�n�"��4��2 �sL�R�i���#���͐�#�RP�,�9����d��J_�6�N�8���M?��R�,�@-�l�S�8�Blz�bl��;Z�Ã�cH���P�0t6:ais�J��CZ*�m@ue�R���lV]��}Җ}�<ۣ�S��� �)��[����y�p@��<)�Ȟڇc���5�:�6�����D�p{/���F�p��u��tfR���b �*1� vI�p��H��b֟�ѡs}���/P,��l�`�h=�ʿb"���n�n��X�]ʆ��H�{~蔧�w�� )�����0�����t̊�zK�����o��bHx9`�c+���$_���}�ܡ�&�J%����>ikti�x0�q.b�w�1�
��U���ʊ+.��p>B�O�C&CE�(��>�����K�[��ߕC����}/sPP���-&�%B�;��p�8d9!�Ťuz�c�kQ��_.����*�f�d�d|�cIJ������bI����~�)��!ZA�c��Qɘv3ՄgK�0�6���
^����ȵ<Ѥr��z~�4y<0��c*7�{�X�u5Ft�9)H%斶��.�q�KC����H��5��AY�X?V�a�mڷ�70�@���n~h1��FPV�{� �!���hF�=�Z6�<x+tN�7�0�>'x9v^�at��1�����Wؼ~��9����(?K@n�*��s���lD�Ec��Wa��C��gCA��c�[_�v��F�1Q�����zã���i��*X�d�P�F�i'�����Z�-)Wy�"�������ܮEL��Y�k��v�!��(�j�i�e:��k"yh���2v�Q�f���z�;��o�n�d�񥉱��;�����9B����/��`�:"�Z=�	+�Ns���."��^ި0W���pX�	SK;���-�� �)>�]E�M�"d�:��F�����2��!eZ oOyZ�W�Ar_9�(P��{#�󎳝6x
a��TN�G>ζ{��h'D��~^a��1���*�#���%0a�~�>��/��c��X����Y�ٖ�AK��B���/=H{��_×��Hs\�fA��~7���we��[�2b-�	^��V^t.��C�]�@�X"����Q�߸H�-5o�fއ:��;&�t��V嚻70 	��њ%9K��mf3i���;��a��Az���:ak�/��1��:M�fH�VSC�g�X�!��8�f���w�R�7�z�𧴏?�����W�01����|�' �`���K������O"{���H��������>�	�.��2��Ku3��Ay�i�2+24ۘ�W=��{�A�� ���%�o/[IYA陶k)k�,�Zv��0�,� }�~���4�1[M�l�4��Y�YP�� �3I��ס�gY��O�?Y_f���-��z�����4|-n��B`>��}�T%i-���-�g>VF�%��"��+��?9��(�ZS�sDs�Y�w�v�03Ѣ`���p�t��Ӫ��R�m�.^pGqF�!U��abӟ{_XH�c�*��/���N�'�D���[���a�]4ci̤���Of?*�㭾���i�����{��ɛh�4x�T*ӑ	ܴ�)N�h[��@7�w��gQ_���9�l2h�R�3 x�7f��v�I�:�FW$��.@'d�����5!'I�3�����{�}{)�_Vn����g��m!,P�QD]V��"v�S�)���O��7Ԓ�t����}�l�WY�_8g8]��l��'�(v��&��E�=G1\Z�L����3`�0��n�LQ�cf�fVR��q�B���L�Z&#���Ab��9v��f��cX���=�s�u�iP�V��o�a��[d��~A����s�ׯ�H�}g��l9lG��l��L��2{.?��9 ��Op�	���������i,�~�2��v�3
�rЯ^Q��3� @�|b&�x 2����2�$�q���F&�!� ҅�����p���KèC�U���o9 \ ���Κ��[�@MHI҇�V��5�BOW^�N=_