��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�/Fw��x��b ayk��]���
t����jw-V��k�d<a�f��xx�Zs��t=ߪk���M��N��J]Hd3؀ADw�`��搥�q��mb����/��7��b���]A�=�!VhtJ���`���2�Pf��i�3�b�Gs��̰�O�%^���rH�+:$���U����88s�ډ��!|�Q��*���bUæE���<F�H}]�1�Ǚ�ծ�:@�[�҈�4� ���W���5|��W�;�h���]C0����0p �Bq1�r��zC�>ּ;g���	%�;g�bo�F�E��9H,�qY�Z�v ��������LӢ��1"?B[E�4�Z���e e�
�U`1"i�qC-ÓԞ�h�d���3Jx����vz��y_p��=z���������tc��dWD����.(�]�T��ͪ�	%��4�>_��L&�#7����L��3úC��0х��0RޝI�&�ܿ)���0���)ק���LU)������0Ɛ3�;�kR� >܁a��HJ9;Fi`�P�h�ʿb�1"�'��I֦M��@JyԎ1߭؎�����O���Rۙ$�_�6�����'�C��@�͚��b̖ w:�[��/���1�+3� ur���@��0G�¶��	j�,	h��%���o�d���)��L�.��i5�2ڳF�Z�Ȣ�[��U0������So�{�?���?�z�K�"O�낇�Lh��}�zR�}�\�s@+4�Ǎӧ����,h]	r���o�m+��]e#}e��pz��S�<��K!ά¨�U���;��qG�-��?-&i�Ӳ���#��կ�jѾʰ���WP>�f</ʲ�4�q��o!� 3v{e����p8�& v�Yb�;#z5߈�*�5�?��Ftr���F��4�ؙ:��U�����^\��E6�f���-3��G�F �y�&��ߕ~�?���]H9c.� �I�s��ӱ������@ę*��t�%��Q1��4���+���2;/<]�4�����ݻm��r�o�t���~r.�V5���y���"��\��_(���0�C�7V�-Rn3��P�+S�ˤ�P��pXP?�D:�px�{6#B�x?���;���tW�+ `)H�P���?D@�&�ǃ<���GdH&q�s��{s��:���XØ�W�+8��8� Ncΐr�PO�m��h(H'��A@_��G.`ƙNZ%Ț��c"���b�����{z��O`��Ez�5%S&�6�Rm���pc�/�I��#Z�R��n<)����=�����+�a�����^��Ǩ��'�	9j`���Ԇ�ʏq���nCe����A��w+���f��o�u~�Q�5���,]?��wnd8�Y�y��,�JH��o�/�pZ�zR5e:C�4��?�̶x����:;�vp{v��}�˝$u�ʰ��/�<P©�aq�=Đ��^O>��Y�;��>�)(U�\���{ϗM�Q�v"	Ͽ����h��t�.�W$�\|9pWѻ�von�ќ�V(�KwfRʥ����e�4�/Ld������������XE_48J����O�_��r�M|�<��kK��5�p�%�k��|��K��S�y�Z�dG�R��~c�����z�����d�����Ȼ!a��c�\M4Rj]�N�,��n���zȃ��mw5�BEe�@���@o��U�ȷ���0)����i�D�t��B��K��<���K����p�SßA}�@y(!�k`r�%���px�p��6JZ��iZ���fWW�7ֈ��_Bi�CmA8v&h�ze¢,�Dz}1��-%Z,H.O5Nı+[:��h$Ŵ3DW&�����w;�gNK�C*\G� �x���L.�>��^U�+ٔ���ـ�V<�(�?"� x-;0~Q������9)���t��u9y�J��Ƈ�
e��{A��K�N<��7o�ۙ�`ts� ��7���i_���Ę�ȴ��-,���I�Gn�{�*<��Ą)d�
-�)zv�v�f̆�,�,X���H6�#��| �M��]R�&�*#�P�XrE�9�W�p-�V;����l2!p��P=X2�Q4��5�\������Ԍ7���8R!W�"��-�Sij�>z���*�ʻ<�;+C�b��-�._-�q��N���*�]%�ӑ�z���pp8��߅����!�|