��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ���������K5���|=��]�l&���,�Ѷ�Y̆P�dI�#*�S�ģ�Z$���<��\i�-�W@Q}��Š�ﰜw���f3�2��S��K��f>�"����▟9���RzV��[nQ���@eU�<����w���Nn�о|9K�S�M-���-˘ԝdT1��ި��3d��<@�Ɗ���V��ՐBw6�W*��� 8ڏ"&��}���$K��K\�y�P�ÞIW�v��{�y������E���>:O��L'L�P���aT?ݑ�T�6-A��X���& C���V���*M?��Ǻo�������^�Ӟ=3�􃾾���^1�6�[{÷����pBA��c@8<#����妭���K�p���^�KY1}����O3�ce���$����v�1W@R@^�k��XbOD���~qv�
���Tn�d�wB��`���Aᣆ��� !x�v��Z�M��h�Tvl�q���g��$/�#ܺa咪�j���w�ݟ(s�%��5(줓P����S�ܡ6�,�d:��B�d�HD�Ѣ(E��<�����4�X�Q��u�P�1�#��J�Q;�Q���������X���딩GAT�����C6'"`{aعڌ�i���QN�;)k{#��.�?ڒ�_�7�.&1�$��r�-F�t�4��ч�%1Uy��P�n����<�l������~*FЎ�mn#������~u^���C3���T~f�A_�	�⼁X�5�j�D�M�C�X�I�~ �EN���+�k�po��	
JZ}��8֝��U"d<�jj�3��tB�8u�+ł5��H57q6+�+�\�����@O^�)ϥ6�"���W0�J��P���N��C�Da�N���Vh�  ���a�k��ɶ{+>Հ�ހwE�=a��&�"F"�0�qL�Lr��o@�~���)"s�B�]Rk�q���q�e� y醀k�U����{j:f���u0C�]#pk�l����(�"(�q��P6�dD%N�v��ʼև�vU����������`���P�U���k�o"շ�LH���_��g/l/c���I��ӥ��)�Y�+��
ζLRB���[���ǭ�Ř��BX�����<$��V�6/��v!�9�v��-[�kf��� ]0�]���y�'��`�I���J������'a�%}Tq�~N������e
q���4DI���~�
( 3t���O".춁s)[����uL%��E�l�{���#���B�(%�����~�����Q\�NQ��ED0mX�yH	L��Y��
ܳ�j��9�;���ǘ�`�ɔs�%�HpD��苸��&$�Z�u��z���+٠��%9����)��:&:hI�+Pq�sk�(�{d������ �Kw��h\�b��fBO���x����ٷՃ�r��ˁ�u�'d|O�M�F�L?���-��p���F�K}�m`�PR=*���w��س�,r�U��~v��a�t�[M�mԬ��U�;��\���H��8�`��/s�o��]�Qo�[c��{��Hgg�ݳ#�7�=�p�+�
�X�����Op������ߗS�q��"݁�kʵ���`��������z ��v�	����n[os$��"�a�q[����̀��0c��?H��U��w��!l�\�7�JC�:Z��݋cϲ ��S"	��9����}w�a���Vx_i��k!/�Q!W�o��fh�� ��е��?��[�Aq�\�sd]�߶����(�~�PF%s�& _�/�qA�{���d8c�fٴ.{3�E�x<K��uH�o�ōs9O_�DU�	�ٽ����t�|
�	OM �9���ܥ*�՞3�"	�K���#F�W)I�T�f& �:L�I��kL��2��J/\k�C��Ќ�y��ƒw"�ϖ���e����f���{�3���B��'���?��=�g��Q�0�J��3������w"'a�(�T�>��B�ӗ=�C�h�$NJ5�	TƠ X $jNq)Fq�8���_����viq5�aantW�̠���.�c���9v��>��ϼ���Y�}�����#8��* vE��]h�ks�x�!?K��GU�U�B��ح��Oi�d.;������]D�B��]_��i�	�1<�m��çTT���1	2M�,��Om����5:PCx|P����*�=�aM/�W_h�F\�[���wU��w��T�&�@��t�1X�c����$r���E�D��9�r.��W�
������I,|�M1F4Ր���-wQON����[�m	.o*�G���+%��s巷��G�	gp��4B)��@ @��%��͞'�V%w�-���h��^���%�pAd��
0��y&��W��
��w������C�s#����L�&7��5�ͯϘ�.��:>���ձ�6��_�����;J:~q��c2��^�����3��lKU����H���еZLXWcc��M�R�sk*��b��P���c��>�ʝ��4�W>����Ik��an��(�U�,�=)�Q�C
��h0@ӫI���Ɋ�(P7���	�:�k��)�����ĿPu�a��+/\�!H��3֦�c �9�Q� c��v�e"��VYl��:^U
��cJ�gz� )BũJ7���rΏ���L��9��z[��9v����U&�蠁!� 4�ʚ �Kgyl��$�ҿ0�p����@_�B�������&��&�{>�H�/m��`��31+�D������@��q7���4<
�����C�ʒ�(:�xVs1[U����B��j9��R�����40$o��ݣ�R���XBL��c�����8�m'~FТ���ryL>�R�5!�������מ$����+}�T�f(?��tp�2�^R5��b�t�EZ���p�h�+��W���I�!��0g��S=�����������DP/�f�9�s�b��;(ʍ�6))��;����1�8?w�_\1�\-���*੎���<�c�f��	rσxpr͉�W�Ǟ���j�$PL,�)h/�
��8�����K�����T>��P�����2�1����������J����ľ�ڐg1˟�j��׽;%���Oz��2ރ�N��4�gu��3a�s<m#�"��8��f�����[DeG�QK��?U�I�o�V^�|D�1�\]�jT��Q��/c����3I�|ePF��S��j��$���{�1�S������ǵ!7�
��ce4�(�~�8݄�e/p���� FAZI��!:]�+H�%�Ai����]9j_��
�?�p��=W	����az��ϐ��d�D��-�A�`�qZ�`�����࿴E ��Ԫ�5&F��c�y������~"}dje�-�R�f=��ҹl���}2F������UFV�i��l��}s,�u���@�2�����B�}1�0��C���'��챱d�kj�o���Fh�跞_���&��

��9p׎ʠ��a���X.�q�;�@���`t@:�/$.0�G����	�ؕ����9��$�#����5:���n��h����=���xFE!U�8��ʨ"y	fF�cJ��#'��g�j�p����c2��w�V��{,�^�f�?U!�!5����Hkm��m01<G%����o�L���7d0��G��_hƸ��Q�J�	�(TX:�	F\z;�Q-5���o�o�f9�)�;��� +�DE} ��C�z�ڭ2����N��䋐�]�zB�*lq�{d���[G�����Ƽ����q34^h�MlI�����1���>�0�h׿�t���-	@�y�� ���a��Ẹ�M%�F�H��������-b�V�
^heP��I����m��j4�/��Ɲ�#	8"��,���\�n����������(�e,����>�|���C�_>��S�|�&Q& $�-+=i��6���� ���?#m���7U��i�,�����E�QI����L��6���\��]�I�o��*�q��8u�t��ȭʭsವ^tb�/������Z�2�"�&��k���8I��:�c�ICùh�˪�`z�t��
/ȃ�p���y�I�@���o��J�V3�o��}���7�_7:�<U��$4��n����z�ĒG�C����@'B��q�m��K+��`�H#@*\\��z5�,o�%0�G?U�d	��q��n��0'#qCm���F�v`H�����k�@�?V�4 Zrӣ<z�D�e�8WK��}��3�w�ՇY�w�.�(�t�Ǧ�����@�CK��$.Lj�e'`>-��~�³�xW���`]��^!�`W_�s	�h��Ͳ�lý��	��?�!�#零́�N��S��	%B*����ڪB:�|�s �F1 �;c�7����.�@OR`k �˴������d����z:��;Z��'r����t�8�1d=rQ[!vf��.�2�\����H�ۚNx7�ȁU s�
iO��PT�DN��eY~�>�]���滊�ŷ�!��ŨDh� �T@x�[������	 ./��VFo����+�#���G���MY�\: �b��x���_�F-�����r ~�[u�Nt��M1w��m��`J���C�* �P�s��a�6�ز�Y��j�zm�}�lJr�N���q>�!�!K��չⳈ�K�C��SEa�:���8��L?z^�(��	�`�h�
�ȍ�خi���פ{]�����d��P�	71�[3�d� 3w���C��w���{��v=��x�֡	>xml�e�%�!�ܔ��#�-�<��DX��D�=
+��d���f�����B���m�Y kIe��~v��Q��x����' �F-0��vS���w��_��Kro�y��M�X��+;�w`�S��ʶ��i���M}��-�V5�u�(Dm��!FgX���Vg	v?Mjd��V�=�D���Y��]3� IPR~,jq���Mq���|������;Y&�ao�G=�C-GeSmM:�RQ	D��ť���3�?}��)�����&ぎh��Y�.��Ap����H�A�5E�(u��%ʠ�}4y'�?x^�6��r�<X��mop�x@]�0{n�G�\� �y�ᓘ��d��"σw/�� �;O��pܜx۰�O���X��}������f����f��@��vrW�-��\
߻�����? 〿���>� ʳVc��z���k�]8���Pd�6b��"�vY�1P�P���7���o[��b@�-�F�$&�#���q=*��''��kR��9t[G�5��\c)ڪ%QF�����_<&I*��Z����P�U��_��ʚ��4+ *3�3�u`hC#5�ee�J�^�)�Xn���U�@��q�kƶ|��/��X�Vmn���'|�?��2_���g9��$$�6&��xMl$����_�l�MUD�?;Ү��e(�P���N��i��I�
O�+K2򏮀| ך٩��&%c*��~e�6L_v<I[;t��Tѭ�g}�+�`UHM!?��u�m��q!��]j*�/�А�+L�j'��� �n�)���`�! h�����Y�cnMä������^Յ众��ڳ�X������c���6e$.�)�!����M��k:er�)B�Q�Fre�s0{u�ˇ��~5mw��Q"�r��^IQr���J�c�5g�b��3��O����ê��VW�.1�f?}�8�4�K:.�*_l���)�,����K}o�1�{���u��Nj:yf��.\����I(S�]p`@#	��a���q?K.5�wt >��&�����?7�v�5�V,�=�|�����r��b���7)���]��q����)��T��C����x7��H�澪EǞj+O�X'l�`��V�:��,�*�a!���`A��-�EO���Uai�&o��J�H "��MD��]\Mz����i�jcW���PB�J=��'.��e�V�l#���2]1V���*朰ȏ�o���*R����n	6#2�{X�&���|h҈ϫ>=�c����Q�('���<U���&]���X����W%[��Ճ�~��w����e�Z �I���FT�d��+� l�T��`n�dG���kL��!U 2eU�7�׵* ?.Epܗ�Z�H��iK��q7�C'\�� �!d���9]D�w����=`���n���'b)���^9�ޒNݭy=OB'̘L���Qn�4:�Rj*�M LX�6��y��q�B�v4�ȧ>O�B�,8���å��2,����D�?����41Bn> ��b��L`'^�~�􊻩'�DkE����3�{Y�l���ݫ	���x�%�~މ=�A2b?�U�w��5���Ե>�uEf�X�*���W�=`:�5+
�u:��v�c��+^:���#/MOc�Y�7��ä�:����*U��k��?pc��>�zrd�b:����i�Y�.�� ����������ްMj̃>���AZ%�������{n�ܿ�k&�3��Q����?f�ͣY��ݕD��S��ȴ8�����x��
�@��Qh��=!3
����D�a������|�Xp�0ڸ3�ʾ�l��Q�I�T��.F.LAv���<�y:)��] 瘚5C��z���}�(i�]!���{�bIM�	 �]/�G_��.��Y�#�U9&�A��.���{/8�CLT�9w�ozm_wg8��rJ����bro4��Z��e�X ���"��K0�s�S�؆���Q��5X �l��B���H��ئ'�er���Hg+k1D���Orה���v�q����1�4�(� ��(iT`PzѬ�H���fҤǼܐ8 ��[��\w��@���Z��^�dF���������s*Զ�@�5�%b�����l�[Fg�>��>*�g/b�.��v̽����fρ��bw�s�D/XK�%� QRH�Y����g���ƱPY|$q[�dP^ْį�,H�r�k\�7��p8�T2eq
I�8F��	�皸�n��ڙ��^����䱩�m[ݡ�B˪�!"*���NR�߯��G��iS=���Hլ?��>�ܮ*��>~#�l�*�<y��o؄)�)���$�ҰG�\���L����7�I�������.��K1�Z7���.KA�>\�ؐ�����!���u�_(�Ў��@���ݏ����4ʉ��y�	����)����n�j��zh��ыO 4��F�|����\���8t˼���+�V.��-�3�~M<Bf�$p_( ¥��#�K��-��4��Q~K��X�L�g$tm����IBoȔk�	hwѕ��%��i�fh/?ƤP=��(�Ցg�^�":�K��K��c��=;�m�g�����H�5���;BsٍNh�[`�9;m��\�9]ͣ�(<��0�Z�>�>.W}�mq='�I�a%����ݘ�NN�Vgm�t:i�	�4�H�Ǫ��#x�h�`Fo`:]�­�~j��B��� �����W1���$�{F�և!�R?~����0�J����'ky���P�@]��|����X�X�m�#׷����;�i��e��١�]̊3H߻#�{usj�uWl{0�qC�lǑ�)�o+���M0-bZ��^�Fʩұ���H��W�j�wR��$���2��t��#��5���G6��LS�Tnt���SP��1:!~�-�7fM�V����RG���zDRq"���#bp���r ֛�5��s�V���q���U�����Y&0�L��V̛�>7�1�9�����1��)�0}|�%0������^�6c��f�"O�"��[��o���MCDtǣO3�.M|!�_��;����.c���!]H�NT}��0j�8�O�V�.�"$������������G�/������!}�-6�A]Hv*�}���.Ֆ��������@m��-����G�$�K���7�%Q���Rp�B(H _Ph�CO+�U[Nȸ�o�wg&X�@�XI3�m�QִВ��}!�k� �� ��}5��~]��>Gs��"�U���l�gӝ���&��0+:x|΄���ءs7����,��yK�&�R��=��?�������5ߨK�e��~'���xV�,Q������*�HQ3�jf\/�;Yv�-_��6ņn7;���O20��`n�Vd���������~� �f��7���wK���e�"���b�k= \W�~,f�}��#K���L  ΎDq����JZ9;أ�#����1k���U|��2nkS�gMr�L:�E�9>�甜��XV�!^2�?n��@�k��I����Ό�As�ۥ:_����L��UyQ�	�6ֈ��s�����f�Vg9c��*���ʻ��+o3;����mw���"`*���e}�/��m3	�C���i ���[l7�{(�="��XVQ�&9���nF�ʱ��y�.�?��h1��A���e���:��/4��a�YfM�T�L|ɽ�p�
2��A=�'2��܍e�z���R���;>�Rvm�@��!�'0�%��g���h�|�J�`���u��UR��ѡ�Z9����w�d
�6{)�^�z)�}(p���KB/��mw�\�Z��<5�
x�SƳs���_��������!5�8<G�:C^�� ���4���!juWb��MzDL���B�K��M�C���BF
���Z�_R�Nb
�"�H�,1�G0�O�	�S�;@|�C�E;�6���m����H�άm>�Tڎ%��Ԏ��C�.�|�8�v1̐)��zZ�m�"�`��2	���)+�fp��\����<�Za��J�������FrZ��z�@�G�+3�
���uu��8b���_��w�����y��W>��yn8���#{t������h8�;W^��?9Jp���g��7�i�Kd�Y�׭r�%'s}ݰ��6&��C�k��O4��d��ӟ�?���%aي�t��}�l����q���*�]���ͷג���Mg�k�e�N���[rF���RK<*S�v�ޱ4��V�!�w��h=�ZI�y���l��9<`w�A���Q?{[���N���MS�,(���ǛI��������KWRm&�{����+x���4o��R��'PwP�p���)�AG5h9p^�έG�,-�N���L���R{��.�&4F�l��Kt:9p��ԅf��Rj3��  f�����auR�J�Ҩ#�Q���Z�I��Y���[�n4�(�+�����(�y�c����M+��%�&0��!��k������$�z�lF����@���'����ofz��2� �)�(���Rk������glх�����8"�4��ٟԌ�߹ �ѥ@���2��Ǵڊ���<���,Gp��������|z�t݄@�X?S�<��R��a����fr���6Ļ]��*�:1>Ӧ^Q.d똰�D��r)�	Dx�f�F��H�����m��[ �`1��~KAs����M�`��I�;p��ԭ� �,��s���]Hd�Ό�*h�V�] #�\d���b��Yac�myEK$���s&E�U�(�\&�G��G찍����	8��&2�F�����I��E��\덱��e����Wm+�Hm��*[������kVS���n6N+7��d0k,:�'bW�Ë���+��氄-�@�@M�!D��]�k`A���@�'�k+:�å�rZ��l[����H�F/"�\��~l��
�c�@y�=��J&*�M�� 4C�XC9�q�O��v���xy)t�ۨ����=5]���>������rY	��.��7N����8��Th�4��A��0so� xDW��a ��*����u�H��**���s�� (�Xy�p[MfJZ��
�'	��a���}�J�F�>�{r5@ɛ9!+�EOF���nu�/{ޔA *�Y�H�j� -tc�y{��'�OF�x%k��'�}+x���3��v`�~��ļ���G)