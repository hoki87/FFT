��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ���������\�'���KgJ����o��W��hne�ͳK�}�%�w���7�D��2�8�A/�b���
ǛUBͳ�������|n��<`9��|X�)'�E�^60.ct���8�
�*�ة8ᆸ����~_�x����/"b�Ԫ�hi�c�5kU�ל�)J�����&��Wp��?<�g݁�;Н���h�����Uz}q ������T�B,�Y,���F��G��ڞ�s����0#G��̂P=�CT{�TЉ!�Q��T��Aq�E�*y��,"�˷�36�H�p3U�D�����s���h\���@���G�朗i��o�K�wx��uŌ*���%�@��5�n��A�u�\�~ ���f��Ӭ�����̘��i�����r�����7VA<�:��v�e��G���V�3��6���9����s~�gU��^�c�w��qb���qA5A����[Bm+ܡ��"#�B�0�4AWZ��^ �� U�Ai�h��d]��R�����rwi2���j�+�q��e*9,7�:3�([&nL���hS;c�O�I�o3��j��&M&<������0hC���M����#zbӷxz�hd�C��j��s����f{ky�k*|��;��=��țp``I�'@պ�M�!�9�ω,��C.V=��,�ŇR%E;d&�(eG�Ӛ�<�rڟQnN8a�kѶ�1��0�TNm�-�+�]uq��^�ǡ�|�8�pk�殔��]��,��l�2'Z�l���]u7��d��6�T����o��]?�~-Zؽ��D���C�q���$0��k�{��M2x���M���!y6�G����j3a��!x9���ȷc4wxBZʹ��r@�ѩ�z��G2�V�B��b�$�w��fY�,ͻ�&U�eyтݕ�	���fd�b��Ut�[u2cj�a��_Y���{�ɝ�X �ۂ�:����e�Dn=/&�`�>��9&�n)�D��Dß��<�6Rﬖ8��,0P�~Ο�T�:�yQ�Y	���IW��	OϭevC#M�Jhjn�e_�Vh�%R3��^L�hd<�
��8�Dh�f)�R������u�(sS�#X�����K�Ix�A��OSb�*��?�Dπ�
��$�xf������*I#��D���F�!97��?8����7V/q���l,�a�C��{߭��{l�='� �nN�u��7�qve��]����s�������j8;��w|?b,�������;�=����}o�	�ԃ'��t�{5˨�bGϡ��A�E*�w~���71����I���ӘT��R��W2���5��t���G�N}�����A�3��T�˕�HZI�EHq���5ߖ��yG ��7�����u'�h��r�G	-f=z����ͺǿ��X�9�}�.=u[KZ����m��[ݙ)���x��?ſ-ɧM���Q&����P48�9�Kq<Z��݋da��.MXYg�ƻF[�S��"�vX	b( Z)�c���4���t)<5A2�7q��+�������,�i�C��@�`���$��1�(l�H+��*����B��|�C���O|��1N��a�؎%!գf��M�N�b��G����8C��]��J�,3X����9Jf� �^�3]q%��i3]�-o^jB0� �#��b� c�WScj?���% �yR�Ա�%
��#)ˣ��j��:	�u������6��=�y�v����.�|4O{�3�ɫ\-��MuQ�i�L�A"��!^�)���5��:P C��F/�Ԥ�����j�/��3E4�ݨ��ᴧ�;���������I�qn�~:�v�U�Y�Nџ��K?��s��9���D:[8�%���eH��i&���7f1e��!��qF�n��UE#"��^�w��I�im���u��B}�, ;	:�{06��he����� Q����o�f�����Ah��h�:c���~��wc��s�� ��ڙ��E+! �"�uKSh�ñ
���p�ߞ��/�H��;|���`��֭���O�ee_jN�\���I7�pC'�C�q�r��%y���5�~�h%�l���È+�U��_U���� _��aمv)h��i\(
~�I��/�Ym��ú^�����O��qc�5:2RD!Y�8=����IW���}(�P��4{7�T�r�|�%�f�p��MgB~�I�PA@�^SWY3���_ym���� �A�`������eT\a��SN�����U��u�J	��C^��q}j���K*�F�Μ[�����R�ok 6�v��;M4�g`2� �;TV��~=��t��~ϋL��楛)��!]z�0
&���L2�������}�A���>mIk{C=Y�m�xa'�1m�ΓRh�D�K�d�I��.�Ь%�\�>&�_֍J����i1���(�y��q8x�c�M�v!C�%Ѳr��G�8�t
�ct��e�|TX�Ѽ�f�����s�V�Es����~X�!Iƒ�����_!�+�8�.^<�6eS�+5�6�7�z]=��!�w�:��t��>`9����v�\���ŗ-��g|o8�"�)^o+��z�<ȓ��];�	�J9~k�Ɯk�>��}��)z������/��^��Y��M��O���W�Lҝ`�x�>�Zyq�E�(���m��h1F�a����$$�REUX��ҁN���ܡG�⃢!�Ax���K�hc��`�CT��h�Z��x����+���*�����t�����vִ�F�ۢN�b<��U�f]�m�-�#�l�i�@$����w�`�VjlRQ�0GQ��Bq���C1g�F:��k��q�w|���ʩqݓ:�H�L��f�h��� [�v���J��O�LRĽi օ��;C�f��H��G��4�n����|���x[��l��-��n�(~�du��[vd�)�S�Xܭ�6���n�V��#���O��q;�5�4O����ȫ�4I3%��L���O]�N�A�����>��/�m�'�DoSF,9�S?�!����8�
]�*�q��)s�&Gl���\�] �8�!�Ɏ�ڎ�_��B�i%�m����Eq��>lJR?|(�:bs�,��6.�ˆr��G�/�O(��~6���0ɓ��]xCD�Uɵ����a�P-��4}cr��~y�w:"]��q׿�1�l�&����	2��_F��{��Tz�+��LY[hw�:9��q]̈́��8�V���(��4Ž{Dv}J㡰�#�,��ޝmt_aR�q��`���(l;�}j,�	��\9�j(���qT��07����wMoW6L���%w�0ǗL�N�]���}���L1�J�T� G~���qokEyڦ>��$�I �s�Q�e%]y���k��N�;$���
R��IS���{��9���壂�c��D5��Ѣ��/�)RQB���w��o��M�n��Մ{��I��?�$��LTl�)��&oQ�e�1S=���5�l�S}�8�h��^�p;��q�s\��j[8�еA��,�RUO��C��w�\���̡�I�E~�׊�Cׅ�նT�k����0� �MG(�R~6�@�[�K�-�2�lQ������XUd������X�r� m�h�{!���q_���Ϫ[��
�苕1��:
82�SD��yŘ"#��0��H��kj�#)����i���� �eQ���D�d�v�wz�8�@W���.����sS��jQ^E���bCu�2�}G�盗��3x�&,Mͬb �YN��x�6�J5����d%��o�Sp��S�^B�s{�(���i�\!o��S��$Z��+\M?�
rNpU|
�t���6���!������$ ѷk�鎵�*=|XJ���UW��ꆝrI,��r]uF0ޖN:���{k���_��wֿ)�!�D�T�t�&z)	����Q�����_�7�z�D�d���vۗ�E�ּ߇�p(�����j��^��㑃�����ZzȀ�V�;����� S�7J�L~CW��UƁU�,�hIc�W޵Ȩ��d+{ykIzB���l��-���M��#�ds��TKX9	�<����j^~oW�����/r��AZy��S�Ѷ��̹/�%��U�O8c��OX4<�[�p�\�S�4rᠽ�̗����B
�Z�O�����W��[)�pÍ�x7��!������a�vì��Hsj=�H�jD<���iSx��I���]���Kw��X�hk0	�\�5�����L@���=ٮN$*<��1��'Y�}WqN�m��M���Ơ��CE�G��Wy]�*��l���G�ers{G�kv�� ]Rd�r�ًOx�3ޛh[HՋ��Sϖ��	鹄��n��	
���VJdpZ�{N��%��=�@��uo �����K�H؟���",���P�	�m���W֥o�*#Moc>j@����k�+����8�Ҷ8Q��IN���K�M�Y�_1��
��{y$;���b�O�YCi
��]�nXe��X�<臙_����-�*������f��M�}���Ұj�E3����;%DY+D��iJMK��5sb��d��2�#e8)�^�KH��$�`���8F�.a(o�l�#��c�(>�^�ey=��6@W�=:uLW�D����5Ʋӡ3��0eu�5|s�]4'ή��N�t��	 �h�Nq4O#�ӷh��Nm�G�Ԍ�%$]��,��wt?�F�ol����i�³�<��F=��f,�P!ŉ2`�*�h��k �2#O�v�A�!�A�(T�`k 2�Z��]p�9��pE
hi!m8�p73�hEĂ��1�z�R&Ac$"FA�M���A3��eK����z |mZU�e4�~y]sN�*�8&;�r�H��%$s �I���9��"�C[t=e/E�:�y��+L�C<;6���4p������럓gb�&G�Kg�
��vTz�G[CJ��Z�Y����ՁQ���a�Ra�Ƅ���y����=Ru����8���+V�J;<Gƽ�A��$d��=*2pf��E�Ǆ*�6��R�J��#�cQ�s�ߩAJ0�~����EB���]�
z#>9�_0��>Eh`�rv�4��^P�#�Kv���t���t�y`p�� w��i� ����y�ebB�h����l
dJQ�l	 
d���=m�~� ��&T�F(24���*|�����p�PNz�1�����]0Vӛ	��H����-�dG��;Ӂ�L�)��v-<%�5�}P�M���ɉ���3��)�^�)��t
j�+�2NM����S������D��{��\�N��q���_{a.����"p�і ������/�O�N�*!B� �)I�~]�_��|v{��5xK|����kiK���5�f*�J��p2~$I���8����7|Ȁ��mȞ�T��/�N����՛�l
�_W�[�B���y��Uݯ���6��_iY�A?�!�J��n�@Cl^�#e�'E�~�	�&?Ӹ>��y�Q�ߟh#���[��nM�@�A$S�����%��E��m�~���םA�j�C��6!&���_63ٜġv�౛0V���Q2���UV]Gdr��3�n�N&;��#R��+B/|yF���D�Ϲ(�G)��,n'|m����A�W�"�>��β��-Q�&�J���
�],eo�� /Ph�q��p��X��d�8���t�>��k�`f�9��g�G�z�zF���
�[�5��3A�u�z7�u�O�pDb{$���b�9'�Z���iNf���1;Vu���>gZ�����]�)��né��!?kYA�T��V�K�W=�J�#�qV7����Z�:at��