��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#�����~H�����pl�Um�v:��L��Q����;�~��?U�b����1�w���`� �2����:S���Bq��6w*��v����m��<�,E�H����,�b�M��1>k�^��&�SV%�n��b77� ��������m?��8��O�07�����v����-��Z�h�-"�f����v�Lk��em.������~A+@$���V�����z�K�Ex�;Q�2���Ij0�P~�ZR[�J�>��As6�a�!9�D0��c7�w�䔋G���ITwߦ�8k��i\˧�Ǚ��3|�İ^?��g!��
&�GCW��'W=+4�E!X�m���,0b�f"����h��D�z*�s;C�w ��j�4�������]eB�帠��!�,��h]��8�g��rͯ��MY��J �:�E���c�0=#n>N:���ޑP�S��U�>G���SQ8Bs�Nk��t%�O~`1	.�%��f(���R1~ZV2�^���dL�҃���1F��4��E�k��:'P 	~�Ny*0S���a�v`3ĥ�n�������@ʷKխ�ڂ��?�%\1�4�Í_�0���uT��k�{��w�2Xi~�6*Y�?"��L�3����L��r��݆Ej�L��.����r���1�b_V0���y�F>����Y���`�]&��G1v��OFO�;7����~�W[�C���X�\���ק6����`��G�E��V���yڢ��#S�t�^���1��>��d�+����@f��":ڮ2l�T������n��<�3_�}�`24l��֮��f�mY����-s=@�y*h��GDq*��*�f?:>�U� �u�N�����n��i8�ҩGD���Ѥ9������Bo@��Е�
ev�A�Y"@nV����#W	?Iu�[�c��no)WZ+:詪�sӈ";e����[�Cl��5'�1�'�r��+���Un۞i�m��X� �`P~T��{g>!���
j��ﰧ��v�N6(�x��2Pqce9mDy�8�Uj���1*[�7�����.�5�ꄘ�Wt��FIC��4P~�e�/�|3��G �M2jP�o���R^����A���ʍ�i����`YW���v#�{(M�	�U�lr�sY�nT^P���]K��O�1*k?R����|�<��Fh+.��w�W)2��b#8��?繃�ϳ��+`5Mɓ�Қ|��_����;�g����̻\�n8U�� ���/�G4l�K��Qm �AS14��m���a��Tf
�߅��qE�t�8���bt�R&ʭ"n�۟�t�HF�~�Ox������/�:���{Z&�4E���J� QI��\�M�Ԩ��z�����E+*0	f��%
���pVu�T�A}�B�c�A<ZT"���q����⡺��`�SytI��s�k�Zk?�c�����ā�.�Kj�#� ����J˦��3uYu�JJ��vc�ɥ&�����1�\�(������9��:G9v�\q�&.��;g �� i(��������N2����L���ή���4g�\� Pֈw����vsw��o�RGJ��2t�v�L���o�ѥT��"C��;f���܍��©5,�0udO��) �vz�19 ��~�Jʘ'��զ�d ^�a+۽r���qо1��.�j��+"����R؄��\@k�4�W��~����p%C���=�Th�4����ӕ+{����τcVec9 m	"Ɯ��7pi��S���XH"�+��%.RݔvƤ������FލG~��(�=yῦ�Y�ޜ0`i>8;�3s���3�=�������͓AZ�YrnѴ����\7�Z�+},c@� A/U��uӬeI���JA&yB_̛�H�x��:���Ԗ���[&��=�2Ϗ��"B��Un=ЋΏ��B�F��g`P������,��˹P�^�FQK�KĲ�vwL���ߙ�@������5YMT�'�$i!+���'�B�
��d׸�DsbH����*1%��;�":�	(^�F��<E��5�lg��S3{��֖rІ�_=�~c�1Ƅ)2�v��&�Q2m�/~
��D�Q_��=3�x���ݟ�vk[�F��Cj��|"��Jy���zPx�`�O���{]�j���!��I��"5���k�������+"Tu7�FD��A`�!����;��H�/Gs�?Q�o���@2Hq��c�ߏ	2%���w�?�p�˲�L�K)Ȱ���2�̷��Q�F)��,H���t�]־Pܜi�i��GM[���*��\�3���{\�;�<�S�-K@h��v&ӳIk�$��!׊�6��eaǑ �2a?���Y�J�\�
���XvbO��_G�@���~�h�s�@;S)�ӂPvՊw#�!.���}�j��͕XA�x����q�o��NuO�ڗ�#�V����=N�H�Q(Pf�HW�4Z�\n2F����9��0�rJ�_�]À��)/lP�H�������STs�d-U��!s~�5�'/�a܂֏4��8��1)Ւ��!5E�P�O�y3T4�· Q�H`�&?��Cơ��C;��v61edDC�we��w��`�W��;f��7"y�/��7�T;�FZ�hZ���'���@�o[�5��*ړ����1����~Y�] ��o#��
�o�޵c?>��ī���޳*1��)܏/XW��S�	:��A�/�S(��-��(U���:��QF6m�*����DT����Sؙ�,�f���-�6t;;� jV��۾~v�n���6{�N���!2Ԍ+,a����?Q��p=�~pښ�MDu]y�>3余WJ#�J�k��&MP���F�j��oG�hU�ѹ����)�rQ���`j+7ݻ���P�$^���G�q� L�:� {T��L5<��~'���?�j����+���\�n7yN�Ǽ?�����Y+v��s�#��b��8���A(y�Y��N�f�F�6F����j����^�ܽ���i��(00��+%\��P�AF�8���)s� ��5�nQ�~�I�O�M�M��,��n�`RZWu��Q���.l�(� f���t�a���{tE""ڨEX�mG�*�{RR��
��s�~���fl� 䄬������R��v�����l��j%.��?w{�9J�7@��An��<w�{N��h��&� #�����R�dG�gſ�Ŕ�Va_D�Ͼ�C���e�`�(	�˵@�@��wM�մ�����N
���6�	�tK���s�L �l�hG�ȑH�������D88��a��i!����ÌN{T\o��ePT̌��.�|{;���[�]��� h���-�=��?S������e`M����)Vzr�����S�u���S@��6��_橴���z�!�eW��'Y*51����=�xU� gv�pm	�S��'(�
�x��A�{����Ye'�.P�k�L����t�E����+R��� 
�Pؔ:�b�XW�4�|v78t{�������a4~vD�]�cz�-�z�8�ɢ&�jy�%���jZo}t���FY���vg�9F6R�	Z,H;�X������_9T�B롶|9bg݄q���+�$���q�R����'����X��׹��.$u	ې�Hi.�������4d}X5+���\~���;AX@[E�V~s__�E�e�}j�$`-�n*��@����;8}���c<0�ӥ͏�G<j��"n*������vQ%�2Z?Xo����TC��i9���"<�jO��m�L��8�	��ִ �G�	��@����3}]����R���Rj��{�!��xDԵ���F�ùL�8t ����ȟ���e8��~a��?�Μa+��Ι�_|����Y%��/��PM:j��wz�A���X?�${�؀�Toٵx�/[V^2>|y��]n�UW�W>:���
�б��Ӎ��e��$�8�t�ksB��:'�ӫp���cgA��Gɘ��~���'�:�JyWIg]%ʒ8�v�4_0�\�y�)|nm3���T6�� a�u�	w��������G��*���o넶>M�j���,w6>ϫ�9f΀���*Γ�.l�ys��K���Ll)}�>2��"���s��>T�t��]є��l�stB7BDp�t�$��z�ѻ��v�Vr�<RWݛ�%�16�҇���	������Q.2�5>8�U�A�#G�8�Ak��Zz"F�a�w������h1�o�1Ch",>,Q\ ��M�g�ru|p�	Z��"�)o�gY�0�;�S�n�v#�:��1�E״3�2zD�t��^a�Y�V~ok�vAw�� ��A�� �ݥ��+ �.]�~_��
�{
QM�O��&�L��b+7��[�"d
��j5 ��u�9�X�]�;�4�+����p��%�4�d�$�8���Xqx��s\���6���xU�	��]Ԋ�+����~k��n����r!k�FD�;!�a�ا�s畡�䈬�(�Z�?I�%�ږoQ��2x��I]��_���!�y�N?�~i�����<!��w�J8u���_r�)�E� ��������p��Q�c���»��+���L�pg�,��%�C���6���}�!i$>�Eނ��<�850�-M�V�W�;����&�u�h2x�3�b���V"��cug�6�ݗ�7�L7-�b�*/8��jVߨX4��u
$8�>� �����zpi�T#��+5b�e�D}��Z��������C�~i�.��/��Y	 %U�a�����������ȧ���+<���'����'�KӷZys����H)�OD�^��A� ����qS�-)e����t�` wn��Y��6w�����j(�=nnA�:T?�Q��E�Y �H�ʽ}!M�|��S%b�*@n�Q��ոD�n�I��V>Lt�/o��X�V��+Q�����Z���uO�v���>^�X�?$+0������^=��/�l�d�-m_��#����L!�P Z��ڂB�t�6�ʗ�;��Y_GE(���N�9��.T@�� e5W�\^��ѻ��z:�!�韤?Z��F��"n�1>h$��k��B����U������ 3u�3���#����������B~#+ȕ����g�˙dn������q_��m�d�����emc�	�w�S
�y>@4�ɋ�����䎱�$0c��� i�¯J4I���H�-dx���Rr9 /����e��pUw@����z�1*Z�����P�.�*� �!��5���<�N�̫��!ZS����1.s� n�Pk�G��V>����(|�B��__�ا}�8��#�f�I�Aq�2���
����&��4$�票!�FS���������ȗ�μ���۶����o÷��Tf�s3���� �����Qͦ�~��PC/9�I^$�}�/u�uJձSB+�ɰ���A�F>*Z�e?tBt��)_���Kl��_~^�7`CSc@�4@vel�HC�ϊv4�X顯��R��	��1_�b�DRj�3�3���`_a٣O3����]Y�� �~ht"J_S������;>�����Z?O>�F\�Q�����Kř��n����5O�#�;���7�z:�����_� \�P��	������
�eѮ�M��;�K7�α!�R�Q���Zy��o��!lP8\���dW��$S�j�\3qIK��.E��V��J-��8~��a+��1���$��4����{O �+_��P�T^j&�a���&��$�l�B����4�3'�.0雨�=(���Mⳛ�]�S�h2-j|���$/�:��Mߖ�d�B]�	Zށ�|�K��.3֒�t.��,IbDU�/�gf=
&-�\����/��ɓ�s}Z+�� {�%�q��y���A��S�U�x���z��W��ϟ+��BA1Gh�E��7�X�pC��e�����;6Z~K�յW3r�d۫Oo4"��5zRQ��"􏆳��˨�ז���9�G��a����LxҾ�n} ����j8Bo�ޕ�t,�0�b� ]~�2[4� c2�J��W��UdՅ�;����T]7�ꤦ{z���:�)e-�7'���H�e�8=u8��Oґ�ጟ��tʩ�$���3�Cah��e�h�D�`�\��C���E�]��[��́����� �CQU���q>3�"�)L��'�[�\b���z�|�ue{�$K����5��+��� ���z"Y�E����1���U��IZ2�i#T?:�*o�����w�)�1g7�ӹ�z{�K?:S&�8��`lH[&�<�A�9ϴ8��ږ/�`n&�? 81O9�(�pg�?A�Y��ߋ�Z�۠�T����tn?�R"�U��1y�[,D}��i���yH^�!��4/�A2�s�����*�0��������$(T���=��(-G�112�"����7�}���Wmqb�`��X��-Y�`o���3t�`B�R����,�q]��vo�?�!B�Q��:�2��w�h��i������hM�I����җVq�͢�.��G�(Y�ݞm�����\Є'R��M뻱��N@�1�m��{]y0�����*����n԰���~Ü�h��u��0�ز(@��r��fȝRQ}IN_�@���++�<fi�n�������+����p��3�p�]�I���U6M��B�-�ͻ��w$��{4 㠗y��VF'q�A :򻙧���(�2D�Xݤ��#h����9p�}���w���O����J6L� ����!��W��]�\���sC"��� oYjz� ��8�1o�&���`�#M �ޡ��"�4�ok��-Qz��X�~(�x��ߩ�4�kD�����vZµ��c��JWPZ�#Gg��m
��_D9!�r5g��Ꙩ��]��(�ӻ�ҖU�4l�b;������٥!� <�>�����e�T~�2+�Z8Ӈ� �S��,	W�S���t.�"	"�� ��#Wi������4�i���q�ǈ�KS�)�<��P�w�:O 먾���9�p�{�Bh.��ϒ��@��Q �.� #A���ؔ7�A�I�0BN�M�qF�C�2<JGLו0�`g�"�"����,�_����Q�P����C�Մ.��'誶��&G�\�Tz<�-����^��V"e�$.�wP�4czZ�*���:�2�L��!v�;���n��:	A웊ė5�5�6�߼��v28�.:���*s�D]��r��h'��f����<�(:�/HIl�<ѻ607	��o�R��?G�~�� 0����������-B2E��f\[w��61��?{��|�����FFy��
� �n�o�W��m�����c�`<�odʨwu6/P��P��%�?�VB`����6rv��'¿q ���z��pY��r}�8F���(�J�?j~a�0O�Ԭ�o��T�mT~�=�����e)>��vM]�����mb�+�J���@�%���)��Oc��P��9�|����p�^a�[bo���a�'���r�[��QGf��1��V,Z���	�F(ڌ{�~Ӣ��\�$;��{��@l��ʮh�B�zu�Zkɹ�5x���EzB����p�^SÍ��<���OX]���o�/�v6/���54A�Y�<��"�&��(�,�D6�F�$�
ɗ�ۺ���G��)��:?po��}�@�R�x\�e�ɔ]b%���WҎ�vE����Ԯ_C7����9�<sWֶ�3*^^s���4�=IHT-[&����A�D��&;t�hm�njZ����1M���0	F����I���wՈ�!���M�F���M�)	Ap���<)�r�!i���F[]��a$,�H�'kÖ=3�O�I���{lGۉ����2%Jc����2}��Z3h
p�`�Q�	�T@,JN-V5�<%�I5,`A�c�m�bT���	�k�j���J ������oe~��
(T���$	��-V;bEL�\R�`���1�Wg���PH��P�0�`a�J��_n��t�]Lf���� ��
��N��=4�UF>qh.�k��{ɨx�|������A
<�M������YG��T�KJ�&,�����0`�q���P�?y_�J�&��\8 C���j� 	�Q�����6s���ч�O�h��ئj��a���r%rn�;c�4��N���碰��O�D��­zRV��r4��@���h�ϏQ h+	�I�۟	)7�G����O��"Wኳ���
����w���-f�{tҜ���kw+���8�L����D�B(���s��n�&���ѹ?�p�)DTO��UXҺ����� 2��P��&��oW�S��F���ML��+������L�o�r	q�Mp^�1�0�YT����)q�n8*����Z,�Ķ��.L���K.2��*�T�o�����Zk�2�DeA���f5��<	��a �!��G'�ό��g��]�4\��o�[Q���׼n�-�c�t�����wF9���������v���zd�%�+��ׯ����m�)��m��)�Y��+C}����RGӟ���9^��7S��f�0��)�>�sP�/�S
ޗ�k��`=�@:�+��b'`��s�K����[�s�4f�ӗ������2� �ۭ��UZ6,�S�ل[@"���0+埚����k�5�ۯN�o��$�i������oCʙ=���#�u�i�.bcn�GT*%�^��ᖬy�����*c)�뺹S�	7Ű ���I����c�ݰ	-�2�X(-s��q�~�+>R��'�bc�Y"/���p��$�(����AZ�ͫ~M�Sb^/^hx8ݧ@�ݢ ��z���H��{C��Տ������g���6M`��y�� �F�3.������������~,�������������x�Ceb�>�P<*�m�q�_ɕݐ9p�{ҧ������V�)t�t
T���	��Qj2�ڬ ��O�Lzb���Vhb�)Nn�X��%u����N�o)pZ���i&a��3]�1h����b}�  �~�;B�s�.��Q۾����@�J�B �{R��'����:;m3��X���O�bu��uo(����Ug�!��',�"�MJ4B�#f�\i�ʱ�3�7��,[p]3����(Px8�����`�Ɔ����a˦`�����տC�8H����lA2j���ԥ������踼HQ�����X+5*�$W����\`����qn��$�
Gn�	K��]-�m]�A��q�)����a[42�����)�p��_4V���r���D�����`�$�9O�k���g/���=;�V�2��R�ø�뭪4�������ƿ� �`��M��jR	����ԧb��od�\$H�� �Vy��ˎ݄��	3�
�L�a�l�_K���DYow��*B��e�k0�լ��MҴ��Y�KM�k��=��4P]�1|��h��$cK���?�X�HÀy �-Ӕ3������\�2x�w�����&���o�ʮ���d Ƭ+�	����a���65b�+<��Y��B� �F�h��n��\6b;R�G����9��mn����q�PP�!�/�`yI���U�BX/�y�;���U&N����1} x���[��od�P��sXq�4��0����Y7a�!�G^�PcӍ	Q�IrW�Xe���Q�<�u�Sj�q�����EV�\}�}���Q4��D��E�M1e�RF-wYh�8��+��,+t:\��2�h���^�d1�@�V.>��T_~y�i>���u3q0>7�t�����du��C������#��&k�y1h�=��2��>�?��_[m"M؄
�mKV�é�%T���� K������5�P̓B��>_<��������14oJ�y��m`����+������|Ǉ�TN~����`1��@�U&RPjA�# ܷSA�_��M~� �a!
�ܮ�en�M��Ĝ!�D �Q�KxM6J�*ޗ+�y�\�� 	11L�ΝWe͟���%=!����.�5���O�A#)A����������䥥��(w�4Ɇ$@��t5D!PAD���=�g�l��D�h�|�	ڒ.n���]j��H/��aj<�)fɢ=�w]:p�M/�D�X�7eJ�x��uSq�&�Z�?`ILh)K�Ͱx�����ި�s/w@$/y��� �aq7إ�0Y��F�@�"�x�#bo������"4��;�[ȉvĭqJ��h���;���{����.!H��T)��g���q"p�-32f8J�$�\��>�n���`�a���ú�"��3>�U�H��~�7�Λ�.��w瓂}sN��.� F��e�e��m��7u�H��<1�
��L��y��|�D�`�M�=I��t��5�&��i|���>,' F𤂛���<���g'���/�nʗ��;AL��
b�E���6W	��[
)�E8i6ιO�� ��b��י���L��|�r�k������Ó���ؙ͵^�b�<t��?�z�'�����xJGХ��-J�c�P6��zJ �,���E�sq�@�r�1��1F����|�0Lk;J���� 3�g{O��g8l��������Ky�.�@L�� ��G����+#T-�|�nM~����}����S��s��)���f�q�Y��8���J�P�u�_�b�i�Z�+��x����IlVH�����X��l�Is��2z"VuҤS1�YCAi{r!�]O�1�w�.W���%�FA
Y�#�b�$4Ϩ'Y��|Bx����wҜj��7�٥d:�����2�WU�������k�2�i<��	׾a�ϫ�U6�
�]/K�41����v ��l:q-����<@y�z u�p8����>y[���&_T����S��Z@�ű��Mx&�`�{OH��n"pw3�����2@�<_��-q��88���E�"s�_T��[�,f�e+�VT11� �XF_���X:!�3վ��!�ݮ��spn@���"n#Հ_]I٘�N�i�. Ya!2
`";;����J�+0��Q�|T���s�����0�Ӝg�Y0!�L ���%����Ek����m����;3-j�Ԕ�c(G-��Z@Pt@�R,���X�	�p� oV'<A<ֿ�K>���e�+��wB����������j6-�C��n�<�G�d�Z�qR�f����<��UF���4Ck0	 ��_��΂1���C(�7��Z��F��ѫ*�:B@�b�V�r@ۼ���L�=�TD��i�1�;G)��GҹW2o�Z��1.�aK�X�&��Ǆ>-5�If��y�ȑ���ɨ��'���~|��f��"1"ر�16�(�"�=Ah��,���$h��/q�8)$^��?6�8��t���en��aY��/��,��T�$_CO�零���T)P�%��vE鲷�YG�J��h�YÕ25�����X�8�R�_��(�,{�i��a��N�MN��{��ݟ 9!��HF�K`�T���@mǇ� rg�9���z��2g�������Pz�K�`��11]-��.���?�pn�HV}�@�$��z[bL��b���h��|3WK O<Kw8�X��s���ֱ�D���J>���B#�6]��|�dϤ%*�ٯ�h��z}��q�o�)��J�� +��o��z��=C��=Y�����E����"�n�ǲ���p���G)\7����ٔf��j&��v�]���������F�ƭ�¡$R����M�#����-Ԡ���Dk�tE*�Y^Ny'�|�'NrmqsʁW|M6�l,��m��S¡]Z�P��7��YX��%�%wA�X��	, r1�@����~Ҳ��v9�Aa���բ�����v'�6��lD���qn�Uĭdd4c���;񘥻�����$�$޼�~��u�ѹ#��o��Pw����L�!Ŀ�/ �����0���S��5�X�Ѻ�ul1�7He������r��:J#���9���v��:�9a�-���H�5���/hҽ�Y�������%�4Q�"�o�����g���P`��M��(���k��o8�g&\Ll��޸`<�c4Fl�w"�C���|>�}�=�۰��>�����m�2,j��mp��'B�ҵy�ڰ��+A���8���xv͑���\v�y(���:��#�bJ���q���B�	�`d��bv���6��%���Q��f�� �9j��f�c'��w�e:Nlpp����%�wƇ����vP�Wj�@���U���t>[u]�µ��	#~�U��n�.��5P�	Z����!���ϡ⒫�v�y��;b�?�̿[�w�:���*��$uO��Kfd��~��Ϸf# ��A���ȩ��rb��a��4i@O(ť��pZa5�t�ٞ+q�h������:C<΅������'�D�?L��� �l,P���X��+ ��5�s"�3�d�Ft���Z�����6�ـow�S�cǵ��$Gig�ϳ+F�=�J9o���V�������^�����Hw�GE�]|ic3�L�ٷxr<qܹ��s����v��=���x@�Pzg�6-$8jg�ɚ�|d������{!�hEn�ص�RL�9���Bq}�!�8�$W�S��������_c�.��+���㌭C��xy�|G�\��Y�<��$_|���1������	�?1S^9V��5�N�\�a������?$J��,��2�>��f�n��]�R�uj�V)�c��12��B�T$"���\�)^���|e=uΡi:8�;pr�&��Ű/�5�ݏb�E &9�h)��ވG�i2il9�����z�G(
+�5X�y�A����F�qHnt`�7�~��{tgNQ��&�e�Ań%��

�o���U��>bV
l*Ť�Ԗ�(mBH��a%[��!���U!i'�d�O�w�Qڢ��mp�ߔ��]J��_�%e�F��oյ{�q�����:�o����VLR��A$:�YJ�+}|*"��|-�u���.ˢ"/.	1]4t17�� ��E��s�D�ֺ�bx.��nn'� Zҳ�%���u�"66o��R=��`g���a��1�%�
���2�-]	G_c ��]E�1��w��� ����)��������&J)� \hm�nDXZO�*2�^��]���1�|�1��_�y�F�T���6�ס����(�]�0��+�������� ��f�F]+����L�f�# �X�`��Sl����`P`��1v_�6/�=ԍ30��՗�rqh��Eי%5qI�xG���PY�njZk{V&(����^: �kg�02�F��� �{$�_�\�FH͉5(��L'\��ݿ����Sm]��$ςO��1g��0�,�#�̐G�ɦ�Ҷ��0=�s��<�x�i���R{�M�*d�c���$��P��g3���;q�;� 	�`IP����rN�}qd�����ߕ�µ3<���FҮ}+d\����p�͟��xXL�G]��cc�"Z�����`�KЮ�#�%����s �ccS]�?��r�����/؉�?������^3z@bf�M����(k;�dnYz!��ۀ͛־��.Kd�s�&"A�[*`L`KIc�$���9�K�(�z�8�Q��f�Ь�Pb�j)�f�cB�M�C�|nK7j�$�#=�Q�g�a
�ӝ����;"*�"p��(n�?V��60��$��#� d�|&���n��g�I�HX��:6Ks����"̀�R���l E	��|F'�g$#J@ql�
��鿨�����G�P�N�̙�$PЮ2n�����32��Dm�U.�ͯ'U@z:�N�1*�h�� ���v��L�N�ˇ���-�F%��\��p�[6QE�â8\��q��P��Y�k��:X^�j�(�s���|#�-CD0�~���B�} ��� �7o?� ~D��g~$s�����Y�	4|�TK5ItB������'��U���;���:E�;Dpou�2~��%)��w>=<�>�J�♋����$@\�O�b�tXU��I�_���M��Y~��u9�ѡ2<�v ���*%���[Bt����@�S�r�~b�E�+%��U�/*��4��+������+�7��eUtnZ@ h��Z�(������c�����\�I_p�B7�eU1����-�۾�UXo�*�5<��&���$ˉ��~��u^N���[j��WC�F�����J���|�^B75�vƜ n�ӄ�6$����>��SUg9~g��^,�S$ѪG��e�fv�{O�	�cjbk���Df����B{X_ ��}�]QR?�᷺H�cڤ˚���E�����8�H��x�@4gZ��v��oO�Av�)��Ș辬)�o,/kL�(��^�K�%NO�.��s�_�[�gF&bR�. ����
���g�C�I�3��X��*
�x�E��?y2�@��ܣx��T
������?U�o��\l*J7�HQk�OY�����WB��rٽǒ��(w�T�R���ֻ��c\}s\nw�� $���9ϑ���b�	�~N��I�Τ�K2f��?�V���L��\LS��p�Gq�-E�b;:��,�L<f�zrȺ� �|	�L��4���ޚ
��V�\���Z-�dX�,x,����\��e~��L�)��Ծ�_
�!�Ny�UU�_���{{T�~�\�b��`�%��?�9�?1��nа���֛�5��L�6����{�����B%��=�����	���#���X7�Y���h�R8Gn�I��V@�z\ç��83c{=�|�8��� I�{��/˨S��v�bS�H����i�{��/m����;�J!��E0��ž]��@X���sA�S�KI�6��:�2����!�`E�?l�<7AD��d�h��t��g���դ��˅���k/���pE�:i�3IU�9(J3��c��w����@��Td���*��y�6�Yx4w/%QVπ���c� ��X���{�_ԉcM�FM��9av����&��H&���"�HX����[�E�3Ab�0�����a�>��!haA��=�����Cb�C�t
����%�=̶�3xj����	�|˫�p?K�q����F�2�&�|-��1�d)^lj��L5�]����z�ٗ���mj�f����p�u����K\&�Hb�'��U*� |/Q3/����XL����u�9Y:w�|ţ�cu�s�AK2��"b���,��� Q�y�|�҅
$����Xj�N�?[�o�A�����2Yy�+k�pp"%�=�縑,@YNUF6^��R6�q�����L<ܚj�ɹm~ĥԟkȇ5�����g�d����д#��~�y����ʚP@���� 5BD%:9��}�JVc������Ч��NB����;��5�e�l��f�Kc�/
�_Qt�y�6;���&���!]L�̭�����L��w%�ͤ�{l���7׾Klɼ�D��΂K3��E�Q��tr�E䱢'�E�k�X"E���3�E�l�2���l��.7��3c�K�˱d?�{y���ҕI\|S�����4�h��`��[�,�d�w6�,C3o�eE(�l:�}a�&%�.b���s�y@����H!�US̖GC�3��)�?b�o�7��qx5��x��GÝ=�\���Qgg?`\����D^�Ťf����5���éI�N��ï�I���B�V�+���Иs&�jc[r0e��X
'c�'�-���4x}]��Tъ��B��j��W�Wg��aٺ#�ъ�t����*
�,f�qh~�A㦗h4��6P[��|��W��&��b�֙��Etu��Qf+�db�9�ITN;��6K���8������z�ф�C`Q��	�1?	��Vq����4��C��Cm��	��3���@�q���iTZs뇡����V��N[����UCJ�O3��V��i��2���~?���Ռ,��2��VD+�j²W�i��O���n�j:��'�`��*�͆�_��z�-�Џ�1-�vhȩ����t���7�-�%����"r�~C���}G��@���]趫�dx<�%i����0yqb�-W#��x[�xm�C֬#��|7�2��Y��p���
�-�����]��؃�©Q�1!�Ϣ�(���yc�y@�U�`&S�*�,#eꉏeN�N&�p��6�`���"h�)&��2��~T=c�s�4vr׼J'�X��|$�P�� �&��c%���.�J(��������X�)��a��x��]	�_V���냙_h#m�_�Wu�-J�y-�g�R�Q�K�.v�޿Ƅ,W����P�X�_2�O@�bڵT�Y7��{�K���Fz����-�L���M�!|�|:�A�È*�K��$�QYf��hY:��Z�p��E��?l�G�00�0bH�E��c���ekm�Ն�$&�J(�4 �%�dN?���ۙ]�$�U�T��8+_~�0�f�p�����;�[��%���f�:4�l�n9`�";�s�+^A�̈�M�<�^/�4[�^�̊A���� �c�P�+ò�(L��_���D([7�|E���.P4���M����d����.2��/=x0�Gs0���V�6����kI��kQ������#!���p�iD���`%V#>��\$��(����-��혛�5t�rRP�m����`y���,B�;���`c���.
Ξ�&�nBy�`��{�g��h�}��-5q<�&m�l�e��~��������b����j		̞or�z}�_GT�������amklܙ\6��h�I$�k��F?��|I�xh�`�o������W�jtT����4A�#���j��ų{�9睊B1U�4p[5�M���l�h��N���B�H,j�ɭx1�+;F}��ȅ�}j,qe9�!�O�g�o(8�.� ��T.�6+2@|�r��\�C�z��dN�SGVa�H��\fĭ�`k[��wVD��F��3y��R��AJkA$\,�1?��S7M�+e21.�L���,G~9��v<[�[&Û��Ùj��������#���
����)�>�Z���|Hu:o{���m:����]�(�z��������x�;Tِ��;8��񎷘lkd��@:8��-?�s샠����)���_���"	�|�z�}]���"T��UN��tcD�n+������h����g�kX3�Ԛ���7���������H��xAmUH��Q
���!3����n	�5wZ2Ml ���E7���������n�F�^̊4��*�v�;zH�ʐ�I��@8�葳܊��H��i�N�Ftn��{4ل��y�h����L̂���O��С}����g���H�R$���iM;����RJ2�~�zjcp�߂��i`����+�H���y3��X��VH�5�|�����u�����.����Rٹ��{�0�Ph��%���ߠ�GE�$cIS�P��N����D4�/�l���|,Bσ�|t��w��#^O�)��)J����t�U��["�s!0����`荔�/��q~�"�aoOJ1_�H�WP�N�,�Jj=^�c�p3H��M�'�]~� D8���^E�ǹ����k�V>�\Hk�Fyx*�@Ǧ�=H������R�ޞ��U4ҙf�o=jcT*����H�E�\~��"�L��xʘ�rm�ʚm����\J���Ms�*:�:E��kaX�ƃ8I 3n]��`���ՙeP����t�@[�w|*3�8��Q�(m�Z�S��e�b�I�ũ��^�؟f "���-��7=w��+p��>tY�c�#� ��d���8*��������& $��T�9�J�&����h{�:���`��:����2!W��8O5YˁD���Gb4������);���M�O<�H��63:�"��h�_F����������=j�s�^�0t��o»�v;R/&���]q����M��b�����Ā�	>�u_,h-Ҡ��V`�z伒���+������yF�Q�J�)�Bj���Coj��E��P��q.�(�W(%s�uY�y����Es����3���u�|V=>���ճ�.�3������^��ת�J��,�����Y�����PX��'0���B�Oo���hO[������RAU]җ��ȸ/�M>7���we$��gd�U]'��L@��.�q���=�t�B���D�;�B<��bLJ3���S̏�#�� ���1#��ϙ����F!�B�}O}��[j[B?�7�-���F&d�ِ���\������i�·����y��];���4�d������9y���cko,&�����P�˺��K�j�_�Y(�q��e�~�2�2��������K�L!
� ���N4��o���c���P��= _c�Xp�ᎈ�Yѫ^N&�+~9W�:�F ����"8_���\���L���~��_������T�� �{��U�!��������%4�rK��e�A���}#�� ������ֳ?>k�ݍ3Š�wj��̙"��2�����A��/�H���Ei��$V1�?E��i02MH)�oDH:���EF�O�_��<�[��-��8��,8�Y�.T�a��jU��9y��ŗ��״lR%�<��-����`}Z���Wa_	(1�E++�	��ʄz,��\�_���J@+J�#��G^t�<r�2���s��Y���~�T�!�S۵�ꖠ>Y�V�f��rt=��UP{|뾮�_��qU˰���=VX��,��Uͱ��!C���:G6B�_��~S�l��.���Ecɢ��L
�`!h�V=z3�.mN���{V�		N2���!�xX�� ��4����F�h����>��2����A��t7���%��Ԋ�_�f���j-�̛B�f���<IO�!(�Z������ԍ���_�UV}���m��a���T��?��m���Vrm�o���.�]��9�35��U�I�*|��>�E�^����-�O�=�#L
|�eVA7�R�"dR�ʲ��Y�����#<��[��6�͍.h�p!�>N	�fdBl�XU��Z�'�������6-^ƨ�ޅ�E�U��ܭR�=�V7cԮ�3���PdZje|�ׯ���	2�|��AI���~a�^`R�EW�k�!#�w׍^��1�A5��7����U;������J�oR��S����-���������H��-���Ɠbr8a0".!�����t�	�!q~���r�~z릩`��R�r$�(�8���f"0�TJ���@�;Y�Dm_R��YMrS
E��� S�lnk-G����Ś�?���\Z�i�I[(BPO�_�+���*��Pl�����0Yi%��?�J��`���&�;�8;�FL�_S��b4	��IBP3�m_%�N�F�;w�5�^U�s�GM_$=����󜇎@��iǧ�8<�ٳ��b��asх��5$�c���?���l�`+$�I��>~��UYeƚ	��Q�m���ƈ��_�16�������&ג�����Tc��ٹ���h���>r��oAD���	�L8$�%��T���sA>'3C������t)�t++��|qj������m8�{$��w0���[)t2��"���f�&���"�������\ף�v�l��1�����V�A��@�c�g�50׫O_!�~珕�93%^v��ԔM�Ώ8�a0����t �×�-Lage��B}�~Φ0�w����qu��0ķ��`؂x�i�ouB���ʍ��dR�3u2gC	��7j�� !:#J����X:du��?�O���q��t������ �u�$�̽�z �'��]a��_.�2`���qĤ��|��4u�{)���7�f����\rhK]�,�_�|i�l���ϫO�^�`�(�_zE�ͅ���dv�nN2PQ�+�D�؂8�J�7k]�}%b���W�[��]Z�6�Tn�#M,���/H$�1�Q�w���D	E�+������!����O��Ȯ��V���!�9m*�l�;QNq�����Qk��o��C�� jUS J�m��s;Ơ����8z,x��d��/��T�f���L���(���98y=����R�"�}*k�k�s��M�t�4Qh�X:/#�p�D=�qXq��%�eCU�Ұp����\E s�z*��W L��͍�^<4�����ƫ�$���xS�$�Z���m:&]� M��*�KI�i���Đ3B�<��P�0�?��7Վ�Xn{�$G�H՚o,N0����ʀ���ɤK�.� LuR���Hrj
���>�V�n-�� w7h�\
�j+*��́h�D����vr[�p9�g�kO�(�&ܖ�ޭ7{�`uI$ٞ�{�Br<Lᔎ�����@�LW�F�;��.5v|(�"��[gV
^a�HФo� ��Ok��q�݌ő��@N���]��Ww�����aO���z�F�4��x۷�j�9ᄏ�߅����1g����^�vP����g�է˯�E"�,��J�8�~�f�Lר���������ޑ �e)�EB0���jt
�j"{^��eO`1�N�xcIpY���ݖ{����쵿�����G� �9�F�}6�H���)����R����Dx���Q2Ch���<���3YD�x��>x���_8��~��$��a� 8;��mkZ��ʥ�BGb�A���q9/��hU���K��]��*_���u�+�4��i��\!&���I*��$i�,�����+V�J��+���9y��N�CD= {���Z ��wڅ�S�L��EZ�K�J�!�����Up���wm���z�-4S�B�������l�eI<��hv�����تg������:bo-J��H�������d�� LD\��[�i��mHF+q�J��v�-q�%q���g<i}Y>����ְ�4�݀_c��z!�XO�]{���3��ِ�}m�o���h޻q'S�_��/����,�jڣ��ƙ*�c���^i�n�,����y�D8}Ah.�ઃHuS�@lkdq98�G���W��|z0�_��n 6������g��&��V��_PSBj- �na��C�uY��]qƋ0t��>���[��h�XC�������>J���h���kJ�:����p�G��=x�-ۙ�a����˾����62E��"�P���Di`����y�A3Zlɣ@N��ՍS��g�p�����V��#[
�o2�&�g�r^���4ؙ?�Q�.������ֈ^�%�>��0���j�<���q�C�����<jr\�7��5���Q&�n��؝T����c꯿S��8�M[(*K�sb#F�'t�n��[l���M4*g�|���Q-�oi�������� t��ϷXg�J�C�DfDQν��,m"�p��Π-�g$6�0�xr�\uH��Ȕ�
<�!��Y�L�l3�����Oi&S~��������W�X-�.�]o�����.����)�}��Q�AvRo~w��ExLF�*��l�5����6�.v�iY��U$�]�Ɍ������_uz���x�����\�2R�R�F���/�����
�B��{�j��#f+@Y�$��5P>�S�ݓ�j���T"XKh��hg\z�O�!�.�6րK�i�4�w��������</��}�dy��J�V4v�2�w�=��"$	�_&���8d������`ʈUu��}j����;d�t�'GD�->�.
� c-4w��,�y�I�Ľ <�+f��C/H�"�Qۨ��Ƌ@�z�Gy.�ELT<��0r�����h�Ki����Ԝ%c\���H}��)�2��A��!��>3K�"�I:�)�t�=*�����\w�g��3E���ʟJ�X�12:�uȳ�1� v�t���e]R�i��K3`�t��'����"��v��ED)�ٟ���4@�O"o韝�����]�/�tmT��t^j;t��F<睢��\]kP�� �4v"j��>�1�x�W�i{_z��Y,�a�=ǉt��7?�����:��|3�7��J���k	h�t��۵D���S�1G�7n��. EatJ��)&vb,�'ͫ��{�����z=�K�;6��ִØ�(�՞"��o��B�Ĝ�G�/���J���o��+�r���	4
��3�^��O���SJ�l0��O_S����5#>�ǆv�%h,`�"2��3����D�jث��k�,���e�w3���G�TC�=��6I3[��[���<������#�/�T@@�R��[m��<�s6J��f�4�&��NѲOʔ����tvl*���*Hi���]�b�/%$Hʹ�^)��V���$�=��������`0��R��D32A��<^B����Q�e�@rݔ|�4��C�1~��n����j/�h;�ǈ�b�q���0Fɗ�m׋���2�
��҂*E�3��:R����[�ߓ��s�Y���"�$��q	'�&����_$�:qz�p�5T��幋��{�Rs�B�xFfQ���ϐv6D��������ѳ�m��1z���L��k6��H�w�lHs��\�Ĵ��
�ϓV��`\�  	�7������2�q��t��K�<�x.���[�"1�IO�V|���baQlU;VE2�@��K�0v�����_�D�3�\�[���j��˚g@<2.�.�z�U@�h�y�d��������e�裗�"F|��U���h���ax�aӍ<+�i� ]$�,�'b��~�3�!o��  x�/sH��U����]M�q72�|Ջ��ͮi��7.�w���@��캎!�J��W��W-޺N��i��`��j�j,��yc@�V��Ҭqv@a7�R@��s]��ʌ�C7�O��CYY �L�^ۑ���sҽ�#�&s�"�rX�g�_�	u^��	����3�����M��X���,HCiN0�S�����B� M#�^q0c4�b�ak�ۡ�$O�q"��L��]W�/��"(����d3w�祁E�.��>����;�.����&s�1փ��B��弄`�d�����Uu����w|�B��iA�p揄��qL�:ӡ�������`Q�}Y@�P�co�b�*�c������mZ̄SKk;��������w� �����d�}8������L�X��?�mp����ߑ|I0���tM4{^�=X8�~:��� c��/g�v�Js&C�l̥!���22��ջ�/B�W���{	��,�|E.����odZ���	g�c
��f���θ��i;�<*3��<mJx!Iw���yŗ�7U����/��Rg��%㯘,���������ժ� ?�#=�u����6ۭ`���UĜkP�*9��v�\DÊ2g���1�@2��d'.9��L��EQ�-�f��kPF�.�;�h���`=���Q��/�.����s�0_Y�f�
}OkgU�'�p[U�������E�� I�bTU�P��B^67��[���a�3?i��[�C�؟3Y��`�G���J:��m����I��,Y35��P�Fj��7�G5�T5��>60��k������� �n'�HB�q��s*�N޿���szzV;��.ḣ�S�=��l���ı�S0D����j��?��&ry{VT}?�@�;���*)�|z|�
�X�}�,7�e���}.
LܔxXķ˫O�`?��Sк����VLdK��N�ώ.���2'��p��qļ&�>���>ԍ�O�Ж��E%w�ֿ8��̍I���/he�-z�<��>Ial�����{��=hp6=��pž�C��BX~��=+��Q₞�a���W��a�a��]7�6��TB�Q�q�)&��Qt����P'�P�, ����|@���N��]�-�#�O4����4K�م�������B$���w{:Knn����0�B*I��`\C�n&�Y��ڛ1�Ib����4��2"� ��>f�}��h)�=&��eUɹeI3M�I?*u�>y�h��L��.�ѝBi�l����R׺��n�w<��Y��ŋU?���vuC��s�_j�/�ܨDt������ۛ\���rؓI�������Y�	GK�����V}2�0S��������&��>�CA?)P������-�t �{zK��~�Q�o�A����~z�G0�z(����\�w�.��[��hlI���F[�=���꾝�AO���xO�	ٿ��Jw�jW�;_´,��o��SB�b�n��(����%�l���]i���� �<��A�������0g T������T 9�y�pe�����?�G�{�;Fo�?�����}8��	�v��K�
4��B�Lǆ@�тq�+N'c��(q.̐���n&jb�WI&Jix1&�.?��׍镗�W�R�����1:�GB7K�X�C��w�����4A�;'�:�q	6�ס>�S�$�'M�,��T�%;Jx�d��I�%��.��E@}�R�E֌Q����sğ��#˩�U},���.�%�vg�j����k�)i�^�͡���`��G�m5�C^j2W��Q�q�_���#o�W^ͼ[�yD?Ԁ��_�2��Z�0<�t�?[�N�d-���ۧfm=�b��pE���Nq��;�����S���B<fL�"<gB,�mG���1�N�p1� ߨ4�XE�8G1�0V/�%��0* �Dk�˿RX�<SM��X	�N-}�oҰ�QaT�E���g�lq�P%(����\�#���R$I��@�+�'�Z�ӵ����+o�@u�"����T_����<�m����e��|�N�-p�[����
��]�"�Y���#�P�3�����[���f�o��h�'49?^^�sUl5.��є�Ak����k�����I�Ã������I���6^-��ed���e�{��ۀ�W��N,$�9R|�z~W�%R���ҡ�~�"���)4'&G��B��ՠ�qn���vs���0���"�"T���Gڶs*-g)N(��3��%��v�i�b��`���dE�Ѫ�ẘ��г����T�	�#Q"L���S��@,��g�����)8�|�jR������u�����[���1�ŷ����K��O�s`�����g��z�գ3���ie X�J�0����֧�{I�̈EO&GwU)Р�+��Ŷ��X�II��
:w5S����X+Q=\*%
��ٸ��g.rqY(grC�d7��w�����"��һֶ����c�0�O*�BQ�r6���5G�_����j���ឹGF��L`�7���mL�3z�1$�����GN�ʯ��ԃ�r����*��y��*lШ�6���^6߼���,1��\q�-�؍�;2���SD��	kc�J`��
QTj�R�����	�^ʞI��D�b,�̼�pJJ�|O<L�y�^E�L�<h戛��o3zi��c�;�ۮ��C�<c�OI�(�2�@�P<]��/Ds�YE�[Y��A,�T���1����䁏H��Kh�vn@���e-�8yT56<	��j�ʒ?�9���0�n%^�0̛`1ϸ��/�
>�����3�LS��ۂ�k�|d�����*�e�ʅ,�l�!�)7�J���Ƭ�GnE؜*��FP��3��pE���m\���-�F09)t$.��nrL���)'��&��
�'@�P���g)�y2��_���b[� e !d�3-Q!�Ӑ�~ ��j��I:�,�ԋ� �@�
�W
�i����n+_��w��JA��#��%C��10dڋA�"�Q�z!N�$K�Mv����W����A�*|��ͫ�骋�_�h����oL �^��9�g��{��6����ɤ���
n\��}}':�1���{%�X��^���C��``����!o<�2��'��!&�r:�0�7��%��/�BOԜVUY��Vuc���:�z!���n ~�Z�>{���}2�T�آ�vBͯl���������E�P��c�9�rR�;���wz�v"p�n�hД�9�`�D^7������J��L�z�����,,v�)��1���D�Ne:�1�l$E�h��Z�.=䊂{����Xgs�2�<Qxa{��Z�BL�4G�a�&("�4��ؠӾ�1�M��ؾ���'�
�[͏ʤ���br.D<H�NЫ�u�V�B���̈́�28�w* /ύ�4Di-C;�9�L{�,;d�7c��~�u'����2��C�S���uhST��r�~d-9'��?����U��<�~�=ܯ��(��kr�\�?H�ӆ�$�hf;�_䪸!������2t�]�,���ta^D�g^�0��n�6��(׳<:�M�"J�G)U3��ʴ[H9A'5:�G���/ּ���Sq��wG��U�-RW,��Ry
"濠�������WeSu�Z����ݐ�|dU���Ta=��e���Ll���a�jc�'���)�D�[�*�D�iV�|-"�q='��#l��4����)zذ@#]X,|�k�5W5΀�����Z��N]Ǡ�|�|��Cw8w�l݇R�x�$�K�'�
���J_���ʰ؜}*I���� Y�����.��p���ʓ��U��62K�c_3����>�[us(���B�����2�?��ѕ��J��g�%�t^���c�-�X��p4�I�lr)e��@�A���-�O�[!.yib�C�<%\�����U(��z.�8\	/H��\�9ڃ���pT�WX�Mv<��PH�LB���3�#�Mw`�G�h�6:�bQжC>$��� ��?ڥK=��"N�_����U4��ݐҴ�p%ˇ>�X�}ܗ|+L���?��"�{B�^_��"�B�E�x�b!8��q�q�W��T:��A��~�jH��|�>�m���y��
^�c$i�3�;=g�-�1����۫��T�t��d��[	��
@�w�hԻ�\K���ꅠ?�v��e��0�4eF���[H�d���,��@:`δ4"ơt�I|:�mRV�+��E ~�[lQ��8>I����Rˏ�ٴ�? �'���c�z��V%.��μ�׉�(�lG2�4,X*�cճfm��䅡)�M,��X�씬o���ڎ+z��RU
�+��jԢ��`��Ϊs�~���Bp�a�)M=@T�ME*����BW��½ws��E͞Qgױ���B���Z�
�b<'�TVc��E�e�t<G�/4vmS�AB���e�P���S�����/5g�O
��+}<4OV�5+��{ڨ�(�J����{����S;+zpFɅ�Hl��< �dh쨱��C#զ]��E>n
�L�Ƌ�ri�?�e{�BBӷ�c .���>�xE����wj�rV]�b���#���A˞��*i������I�P�,��_���:H�.+"��k0Kj�VV�J�7� wu���6�b�WT����^}���G��3g�z���SJ�`搠SSJ�5l���<�˷2G��I�&P��O�Lc>BZڵ���Pܫ� _�n�]����:o�Y߹2�ळVO,������d�m濕�.��n\�'J�o��Գ>\/���/���+�� �p+&��:a&��L�B�@L<S�I���b4�J5��dO�����_��렸\���(�x�=C�=�BRp�E�J���b�p8�0�0E�����A����;/o�A���<��D-��#b�vX�
י7�n��W=�8� ����-�9��T��G���:՘�_�[�
Ҵc����Dʿ�j��{F	xw<��e��Ky[b�k��Q��%�F�?E-��@���՚�����%�j�/������»��L�l>�(�`�%>`} �|xL܄d���)@B@EL��;-V��G�7�y��mz�v/�|gW�>�sk�K(�zL,;�����R��͘��A| ���P�Yqx\�s���ɚР,�����ɓ��>^��k�ZO���ȡ��q�?X���j l�1��iU����O�-z��	��v�1���Y`�O�gtƩ#�e�ӟx݇���'��1�8q�IB��ڑ���՞D>W~_����9:��+ȥy����Vj����i��;8cy4�������j����%z*�0�13�"�y�}�0��$-��R��HT�I�X��|L�EI�н��G�m�-�.������S#�L!h�#�I�14 �g�Q�5ByT��0Xq�3�Y/�2qR���R��$�C�ng���'�>��d4��7��SY-?[�/�ygd}橼�d.�f*PoP����0^56\�(�c�����vADf�"�������G�-�z�_��O���9��sN��M蜻�H.v����Qb3�VU��A�=#��bV�^����Q�^�Z� �^���P<a���vgv�bkΠ!�y�5�ӓ��k!��eA3wQ������	u��)7�?���F9-n9�`�#�7j�(>:Llw����[}-��5]VXz��tK��n�l%	��!p�5>)X�>���T�P5�~j�=_��x��U����K4a���}��a`�>�N���瓗�$�D���f�:���u�G��A{S݆���.���q�6bp_Jfoc���g�;��?��s&�;k�P*��C��_�K�>�^L��q����ֺ\���\��"�O�e�/��)$4�U�^OqAn��c�§���~�I�ӹR��U�;�N���dʳq�Y:��U��e�u��u�&\����w&��S��P�ɧW���Ȏ�
�P �D3����x�Ţ����h �p��Ӿ�A%��yR�l�v�_��q��|�A}Sp����_�l[
 m�����*�"S�f���v;YV�^R�|h��� '4"y���+�[�VWČ�߶��g�KZ�^{����Z����:4��z���#k�H��TCX,�Vl�HC]���v��!����s%S$�.Z˿���9���p�"���d�ܩ�Id ��G<��‶_��'EΨ��hB�y&��c��M*��W@J��
�1QM�%}e� ���v5�Bň��DH�(w��*����􃻞���?x=���������~O�Km�$K6N`W��	�
��U�=��Q��ڈ�~�E�"	�I��rX��#�a4�e�~	:�Nj�	�Y$�;�~^�Z��ޒ����@�}��[|����̎��(�~�`�տ�_���n�R�9���S�E�b��Lm��;Er���Г�H��.���Ȋ�w�=5�gQnDaZ5�6�c)��֣4vQ(��U�(f����Ouا�e�O�*���!_�i���(�I����l����?C $���4`���s���^�~x�pDݰ�gJ��y�Y��qn&���1��̃[�@q�X��&�38��|�d��?�f��B���t[T�h�=��v"��$/5��ƘZBy,y�K
��g}jM!��E���p��$z�$4J/��'N�=#� u�L��H4�gmYv�c�'���B&�c��њ<t�Q�(��}�?A��������Q���<	@e�z���y�%qR(b������Z큳���{|�P��v+҃31;`Cx��x3���B��ltR�4���|�����y5��p�8�L��B���9��Cir����wK��Vm
��nXP�q6R:�+�#ސab��B�{+ uj�ҫ��M�
X-�f0�A�������PY��3�4�\'��(�g�)��ZZ�j�O��1����?D��J���Q��� ~i!�A B�%8�Q��o��:�@�8E��qG��^���o�d��¡Nl��3��Y1��L����*�:	�ݽ��vj-B_����ńG���B<��"+o)7T���f�;�ý��0��c�l������?J�!@~*[�/��6}�:dl�P���O�N��π���@���-����RbeL[w�$Mq�S�p�����@�&n������H/�e>�������i���y����M���Z���_��O)���[��~����d]��n��GA��������NNO�3:m�
��m�K�P:t�|8�={�@����:�/�wl����`�����w]� ��S����@tO�	4���}?�
����em^�ݞ͐�+e)�{k}4�Π,�άy	�D���x�J��)i�߃v�3W��d&`ܧ��݅�c�5�I�	$��8F�����p�����]�c`��D��{/�{��F�^���^��
s6��X=[���]Θے�2u�@�9R���<'~�N�~����8%�S&4��kO
�3���HL��9��Y�1�����s}XN��I��F�o~��U��Gl�Y�\�%�*��;q��V~����[�|�+�Ã�Jvaȉ2���H�@��B��kؗP�wp%N�a�H�� �iqI��p���|g�PI��b������z�{�V؂y�k�0X\nDH��6�c��'.����k\2��Z����t<ϻM��Ɋ�͈��q9@��=�=���+0� ���9�=�9�6ŷ0��O�,!��^��X�p����%U��a�ƄM��G���,�)`��d(3vR����p�C�J�̭�>�F9j�^�׿���2=0*s��~t�T�9���*B
��-_�t��2_����u�qȲX�����J+�|:���渨|���9����uuU��V5͡�`��14���Z�4ࡅ�V��d�*o[c�>V����p�[��x��C�[̴ @�2�LP���ԑ"�����j�^�<�s�|YlB1+�/{�h<	�c"q��Ԩ�vǦ�O7��=S���VԴ�@E=N��MD�����Ϸ���O�vkFCW��������;8wJ.�ax�PD��+Pj��Mj��Qk�����k����f�����(�}�:�s)WiY~�/�b���E=�܄�
MՄg�_��+A�J��'�h���¸�ݟ�t<�ZY����>/G��KM�'+6��מזj��=�Z 0���Z�@9�� ��~7�E�͔؁�հ��fU^M��� �oy�@�r�68G��X9�`����,^�T�e2vF��gV��?`<��xe��_�b�����#ݢ���?i�nN�mEܾm;؜�S�8#�ų������ ~'�z���-�a�7��\�IMF�6��BM$�Sn���ogJ���ĩ����	�Q�ENWi�Ǩ�J�x�4���m_�i'#�t���x����yE��:�mƭ)���3E���H�ɟ�5��O��������/�2g�� g�$ӥ/1��p���"�UF@�E��L ���]�H��+[�*xN@F&a�F����?��rP�tr2�$��xɛ�`�E�؀�QSɧ�֬Հ+�>W�G@~jxDx/~g
��Xbg�}?���GkUp
���8��9�G��;�IY�I��IN�*0H���i��b�9�B)�t��D��nʣ�"�T����4�q�����j���.z��U��N)m�o�-����:_"/���I�]�*�:��M,t#N,�����P�M!�V~����>�IZ8]�S�=�0�F\3�
�PI�?`�t$z�$�ra�(�������lFٯ:}�^=�����I�.�0�:�"�Y�h���K��訠V(-�ǆ����eۣ]�3)qQ���o��+�Li�aѷ�D�N�(e �;;�bK�9��;N���o|D�P���ĕD4;1�>8>Ooo�(�a�#�#�II��I6�-���!���tpA,��^�}Ϗ��+����MF����>�f���g �6$q�(��sX1�X�f��F�Cw��C�7Yw�n��E�V��w�����+0�2���(�R��ȩ�^TOci$+�+�+q1@���Ҩ���B$�n��)hq7�j�R1��l'{s%c���SJ.��͇bl���m��@苔*Hd7͙�@_��{�B(�'<l+GO7�
	��nd\�~�C��/�~���W�4�I�H�A0f���4��������e��������ZHB"D0��᯶��u$���@�w�Xߟ�6��z�-�5���🏌ɞ�	�K�_�&�`��'b�DH¸Y�����94J�Mh<�]�+

���a�M?ݱ����&�6�ޮx�)���^���?(U@	��#{��|q@�-]odߗ�M��QRƗ�<��~�\����u��`��(�g�A��+JY?�_�;ӓ�/�L����;j,�E���q	�Ql���QWU$l%�����J?��D��'���~��7[��d}�b��K<���-"���F+�ڒ�L
��R�i��׹?���Q�Ơ`�, yMM�N	K��PBTN����yS^���VGB9�Ry�Q�Zb%���\������-JC���jG�3 �;:��Ӎ{4�9�\Q�	���Uh3�ZHŖ�$�Ѿ�z@���׮7M���M�uU��� �7�Y^��d^���Ef�h%��ԅ�R��~��,���[��޾�����{�~�>��B�W�.��o|�L>�w��BȽɨ�j���?�\���H3jC/�:�D��V��@ܴ%��t��%�?N��YCTtim�ZA�^ p�K{��(ک$���5I\f�iDTߦ�^�s��ǲ>���E~�LR=��pڴ_�k�v��_�JsRq=��O	�*�.�CL���ӂ=Qz��6���~*J(Ǵ�q��y���bze���eP��[{Uos�7%O���g�/5�46��絆s��p�l�.��qi�Cц��uќ�-o��ǜ��Dr�4��6�'CG����I�!m���a�����h1���{"���n��I��v�@�FR��`��<-�W���~�>jm[�Z�fq��|�������OP3���X|�9\Jt�����g	Ya��-;!��i 6��Z?Ǜ0��~|�0��	�g�)m��S��3�F�E�@8��G"K��J=������O�go+��3Z���X@���|
���Wf��u$���.��<���>1��+���,�Ww���>�m�� �BF�����L�W�Q51��x�4�݅������-��T$��,��p[?j?�;l���������i�{�uր?ҥ[�[�f������g���=B�+8��Q3U�8&��0@�Œ���tRT�`�d��=Ig��ǏY�sJL���C�P����z�;k�!�	�0���,{}hV�zt�S�r���p?�5��E�R�k�Agx�fF�jp��@�����[���Z���.��SAV�@��C���z�5Lm�҄�	��iyl�uT��t���U�T"9���x�8�K�M2�/�٘���$�Ԇ�1���Z��%����D���A���������r�mODKe��e�D�A�bh���kYӃ}}�T�\h�(���+v;�אjZ�m�ᱴ�Jt�0�����f<cF~;Yc�G|m��<�Agdp�T��8�c�GQK����,zH�l�Q�l�Z��+=N@$�'u�l��KB ���i��B�(��U���ȚUБ:�y��_7�WJb/�܌߼} �"���� a���b�v*3�d�NY(�}��ߪ��e~HBT��i�������	�!:�DADT-�U�q�z὘-*Vi�]�}O����7T�d�&�e�	G=+��#s���a�(���K�'�����'fQ6��>6%�3Y��Y�0Ԛ�q &z(6�<���*|^ݠ��N���d���D^�'�d���x�[�+P*+c��l����D�"�J����������v$=�1Sph@�E�
��[. <v�Rsb�^�pJ�iJ�g9D�"�k�3��D�ؿ�=�bB����x���]���5a�
$�G�"\���"lL
PZ�R$.�/8���=;w��E��Ҽ�ʃ��HBȢ�jG���Q/����zf��PH`������P�&��ɑv��o���Jme/�Aq�A; >����l�"�Ul��L2����yո�����+%�F���h��t�"4��8Uq��0��T�Zu�#	��2UI�,�DHk�U?�?�z�������:�~h1��'m��+fޕ7��[d�M�߈k���7o�Sԥ��[�-�%(������(3�)Ν�REt�C��U��9����4"=�����9�]�/F;�+�
���u�?C5��Q��<D�ڭKy4��&`�bRO��,���n����>���3�tB�º����?��ydMh%�]����q�H��(�+\g)X�2�������.j���f���2bś���oy�0w�<:J�y4�> 7�s�����Y���}0gս�+A�=�,��ņ}���l})��>@�
�T���i�a�`��u��d�u~F\�W��cj:�V��JO��Su:�n���� i��cE���h�1`�8?n��oe�����Qg?������� ���Ag��<��C 8Q��j	GLt"���u�j��"�ꇀ�/�I������}mB��-}AN=�#K����6� ��u1]�F�#���LX~Ybf��r}��&8����Q���jcT� u����:ʂ�L���g�΂4z�C�M\���{^�f"�e\
z_��F�
WY�_�٪)+$ CӼs����v�K�⢥���Ɯ1c(oi�>>��mbkz��;bթ(�DY�xk�H�S����h�7�_�� ��XL	v;.����
6~)[�� rthݨAP\*rG�>��Dئ��o�V��_�e��:�"@�r_<޿��oء���O+GN�sy���8S�{M����!�����i2��`�/{�$���6�A��� �	�tm����gdy`��&�Sq��ǎv����B�5~ ��A0@�DSe��VK�(U򙫾��3mJj*�WW|�f f-��-��B9�f��J���2}f����˂�_Xtf鄙y�>���yOMu>�QP/�Y�(��ci ϛ��%��1��ρ�S8Gv�T�Û�d��-�f$���UX܈ɏIϬ�(
�oҴ���c����x���74}�{r������GsΦ|?�	ن6����sn���u��e:����,P�Ww㕏F�l�ˎ�Q��f�3�e����2L���p]�8E�|��Ӈ�x�]�:Ht.��4���v�îI�&=p8*<1do  .Z��2�[��C}&Р�\uD��cę��D%d�McVJ�e!l�M�Wh�J��ߤ�[y޻����%mQ�F�FE����	F��]45���FJ�.\o.&}�����F�y<金	h�]������`nłr5�����4�i���]&�)eJ�L�[�&.������}4�����}�x��19�8+�Fo{&!����{!�=��=mx :�b�
AZս$a��D�v��>5�Q���\fG��8�I�&I*Z�U�,o\��?dg���E�#����C%�@��&_k3D��s"�R�Q���N2DT��o�$�*�dyuN��Z�H�^OG���n�Ɖ���?��!>t��� 3�$�/�V�G��߻������"v΋��iq�g���������Z��$�L�e�ǔ{�={�L�*(�U�-�n�X�~�{w��+I�̄,T�rw��o��X'�h��:��J-в�&_gs��o��W���%Ɇ�fc8LZ�r
L�Sj�+I���MFx��������U�&&��U=nqgW��ef屪=�Y���\��L��b�V�_Fd�Gy-���*�md�Z@�Q
���܄�Z$x&C��њ2����&��|LG�?���y?cI�p�C��	Z�ro�ْ練xL�����)�Vy���^@F��e�������Y��a��&�ڣ�l�:7��#���F����;x���k���n��pQ���Ո��)Ҩ�aj&��QM�Bo9*U:�Qp��}*��3��|̇m	�s�Xd0�e��������;��}s�� ,FQ��g���6� &��&�(aӻvH�3�.|L�Ѐ���oe �N'@�ֱ�"|ʁ+�$%���\�k��zq���W��o��{��ݹ�j"�JIS4m��?^F�����)1"�s����tѮ�@�O#�~[�ҟ�"������A+��3K���O�fez�mq?E��,���������)϶|7mIVT���Dp��D�$4�ը��Ji,O�%]J_�}��a6�Z�r�}y��XOǜ��0�n��E!�a���H��u\/zaG"=�/�����	�U������h�숒�"x����=�@��d6v�0�(���3gb> ݎ��5\�%�0=�g舭�%�������ʻ�2�N��u�2��6�aa��=����ڻ�L�D��X��]�(z���K�앮6����
�d���QUY�o�aS��U�#�+}	�0��T�v�Z���Ɖ��!5Ez}� �0a�+���!]�H�QZԡcW��D����ech�(|�}�c��kw���D;�˳t��tv?<ja�{A6��g:�C����~>�ߒ7N������T.������S����X� 2Tm�y�@}PO��
W;m=a4����F�O,I�w?
Z	��W#��d�v8�����O�����/��9{�&�j��1���FXcS�́ Q��>���qQ���{}|�nX�Y��Jt]���XsB��=����B������r����������8נ^t,��+�F������el!�+��x%�§� �� �ؾX�Z&� ������F��Q�q�s�����|�'����a���X�Ds5wj�c���1U�P���̷����.� ��uȒk������;�y;s�v�]��+�#Bo-��Y^��P�$$rˋ3Vg��Sĵ�b`�(gt�
m���D���0%@��N�-[��Ю=�*�v��{���ı{x�*%��d���u�D���Q�r-�v����2�}60�5�[O�>�нP:�]|H4�n�q��1��h�3�];�
�2N���8���l?e(��A��B%����K��x��;�n�i `�������I�')�AoM�N�)���ەX�!�U�x��k�k��(э��*���ZX'����{T��SR��Bx�rOD�������pNf��,�����b1<�/Q&_�a3�*�ۦ57���]���D��	)�q��ǚ��j�Xk�|x)+�uy���)S-�*W���Z9o��c�kI^�*�d�%섘��Ũ!u��q��>�p����k�7l��^�|��wB�������?�-1�y裏��<WD��ȓ����n��Y�d�D���)w��o�0�gQ�y�'5�$5ZV�b[B�Ò�8����%;uT�t7&�����  dm�o�R���˝Λ'���D�m;p }:�$��Y
�`(>��>!b㌞�����;�FwV�!xE䐤�dT�����o�B���쀲���U/K�ľcu!m�2S����R�ĽU��XA���8��`�C�fdǜ0W,�K� Q��w]*�̍�B��P��: 
�T��3!z3'	%=T, D�qA�Y���<��T��� �BJ��pA̗��s1V��t��z�Ĩ�%���*��I������l����Y�O���:��Qh�g�zL�b$}�+����,� �@�~�s���P39�I�����69�I�I�Ubҷ�1-�[yպM '�ݛ�AI:�d��n_��7�����cJ9R�U:�ဆ�{����~DTF4	E)s��Ȭ�0��ѝ=7w#fg&���>A zo�M��i�UO�s/�'���#w���`((bp\�st
�D�F�
Ь���'j~.U��[s5��D> ����`�����]���Y���lIA<�-���;-���?N�&?l����n�u\�*ӑ�������}_�-���nt��g�6QLt
dx�h�'�
I����,�{ʒ�d��М��3�/U�j]�Y��7��A ���ѱ���}���x��0�E��gbt�S��mA�ݬ ���G���y=x��-�p�%�C[�2��`�&}���>����;�Ho��<�;w
�� ��+i@'���i�E,��y�L~W;RR#k�Q�Ɖ�؆�a�O ��k���:�7ؐj��2���|.'�V���ӔQ��%�� Gf���^E��p�s!�&�I�!�C�$pj��4˟��	�+M`c'���6mo�g��MB�h<���g�s<�ߟV�ŕ�k����A����:�$�,��'��,���?��P�� �l`��; �u�<)t�z8];��"%3�$	f�*fJ[\>֢��2=!8�n®,�bΦ#��'#�P�@�>���HQ��N-0����@�@`�dS�T1��jf=n�H8�UDS���rZ�N
�Ց;�c�vx[��6�%-�����@�J��=�q$��$~�@M^�Q��˺8ܠ���8���p* �(��3��"����	���!u�J��O�����px�����f��|d� �e(��B��(�T2Z�fc�+Q8t�tlxP�!�adOZpÐ��ǿ�uFnM�W}��â1_́i~��Q6_�ˀlmw}��΋�d"1k)u�ŎEɥ�� �l�M�W��Oİ2���!j�V^���P��)�m���aZ�3�bJn��h��<��Zo�ƿcL,�ܗ�p�؎�]��V�.;�kZJ>:Ϯt��Bŗ�I#��na8�& Xe{��XX(�o����-PY�H���L��Ƌ|m\-)��p��Mnk����Jxb�j���T�
�W��=�g�	�+�Ee��w��^�����?[#�	PxN5=А����/Zk�:	�=�\9����|R:�P��y���E*�h-��A��>�y�t �x�!�Lhwx�c�E)�#�T;���0+�d/�Ak�*�H'���	��V��@�:XpE.8.8������&�"y[�ϩt|9�Bu8W�[>i�����p"MfE���
ZY��pX. {�n*6�2Y�]c�� ,�FE��#U����T���$d*���H���'��c�I�����?<�F?���=��l��(m�	��wh  c�H���9e��T��g��n����Ay�Y���_ry�A���v�ġ�A�`#���[68�u ��+��-O#~�߰����B���(h�����4c����� V�W���z��Ɏu]+�D����ia���Q�_%��h�f<B��c"���+�U���(�� U!���K��\�^��,��t�(U��[x�ώ�T��K�@�ٿ���_��Y�d ��5��e�Cd>� ��o�����Sٷd)n6��!��!9@�[:�� �s��餴�z�xk�oF��e\!\t�D��*����:���-<Qx��� dT�W1Dȗ�	N$u����0<9�h�s�O���rq�+q>���O0nӓ;���U �e��������X�	 �;#D
��et>xl]!J͠��r��-�jjwm�	M����S�ODj3�y��-ŭ˃|�;�IyQ'�V�;%��͢�5n� �����?0�-��I/Z�j���M�Ӕ8�7���?z=�i��èo��#��P��5�a�}bX"/{7"�d�KI��SeE)��F�§ӊcm�׋
R�2��*%�r���%z6@����)wD�i��Jq�@�;����wD��%�0\���Am�~���-�w�!:��L��d~:�b,p E�*%'���
8=<��d7P�*�^���!�r�K�����&X��>ʽ|� ����>vI`���'���I��<T�M����'�K浬|�bA{?�����po2��^"�����0MT`�t�]�Y�*sytd
D�}�:g
o�����=��=�R j�G!j�aT��7*|h@�RRgN��_�q������\�\�@t����[¡o��Q��#FS2�~���Gx�b@ט}%��2y9�K�q��d���9�W�+��K�s]�<Ū��]�G>l�_�"��A%�N�yR����3� ��m�t� Wt�K#��ĤA1�p5Q��dRC��]dI�Ґ~f1�-i�vO~��v?o�Z���~��2�T��D<ԴގS��]�H��Z���i�47b�I1�\�n��5TI�:�r�3T�(Z缫-J�II�������k�y�ν����`vy��T����E��3�y��߰��C�����x'3����0�C�f�D�?_���#�CL��FSAM=�WK�1���6v��Y��w%24Sq@%p�G�䟁��65��얒��\�V��%cԴ�*u�1L�^A��"�n�9�v>��a-≒v���HA���t��L�!J%��[X'���`U�˄6�m����w�����մ�[
}��8�J��;�W�?�n\���Ԏ��!Vr��sQ���8�j��o�)���#���$
I��`y6vJk2QF[�R"#����Q����(�LR|�ƒ����""���q`�����p ��@���:`Zh��5g���Û�,���Ը*�_}��wt7�)�G	��C-Qa��"���y�]�}.7��B����*.�a���
�%=�)�7v"���oV�q^6o��P��ɳs6
�����>���ȏ��U���ٻ���iOZ 7;J`Q܂-#��^�6�������BɶQ��㴤
�L���6�	�y9�,�d){})�إ'qոd0���#R}>��L�s��Y 1�TS��2����p7K��0��N���e�N9R{�7��p>�[��n���&�%]��p�?2C�0���T@�0�tiJ$c=����Q5�]�l@����}��Z���fm�E�:{ʓ�u&Y�q5|cc�V�NV�rG�ʥ,v
��2�% �,2��j�|�#T#9w}�v�����5�m������4�_ �63�^;e��(��@*Tn���3$��r/��B2^�p�)
d�\����bi9��-���z9pz{��B��1{��ܧ��Z�Eb����N�$d��^�UT����N5�E7:�?�D�/���{���]�Vu�h�t�[H�F�k��%r�X���ü����[����^�^����`�M5K�7�̍��ھZ@w�6n��ZS��y���*��`���� ��7���	mU�K�,H�5#sL�)�ۦ/ ǉhl0�lV��*J��}�s$� �3ơַ1��U�X���Xj�w��٠*�B^�~Z��<��Q��ĵG�����P�0�mCpP)�	(�
_��;��]�؀{��&l�b�-@��EA���7�S�� ?��]��/ټ��퓛�e�k�i�|��n7��U�L� �^aT���������Q��pf���� �tw�d�� ����e�x��Y�u[��2^lj�W��)Y���OCMo�Y�}ucS6�h�	@����(�}���"Zr̽���l�\ua���<������V��f� +3��2D�a^)o��;�Ulh4w]v�&Ѥ)��Ǭ�㇝����g���(mV�%�`�O�
��92�i�J�>e�*Q��Ri��;�m�GX�U�c�OL��ف��KKZ��-�m ��9�w@�����Hk��y�N�=:�w�����3l_�x� ��	��	�M��
��#�ڣKl͢��R�YbuJLxī���>��z=�M�U�%���]4��d͏�ǜEe��Z7,��⿄c��;_yP��>��1]�"� �o��PЩ����#8#sqe��?��V��qp�8�Me	
S�+?'��� �C�֪��1���$t�3������Қ"��O�2�,�4��;�`�}�mC����+�!��H~�W'�]�W���:,�7�1���xN�ܺ^@uX����&�Yʅ�����q7ӓ����1����_'�sQJ`h���1kXQ��~�т��{A�Q(ƽblc͚�y˂WfL�ɡaX��œZg@💲���A_�τ-76<%ٿ��&X7�
?��Du�N�����RV˛����b4���HAa�]
����;<��`�fs4�L���v1��&�R�+�7���O�D.���N�a��^��1�	�'&���PPW��z�~=<�˒Q э�{����m�&���A����D�W��R�*ҔJg=s��,�Qd��A{κO� �B)ؒ�j��m
�W�u%֫bhTVz��3��+�wm��).@U��]~���Y�1����0�j�5����β�	�*�0:c �D�/��)��q*��	�K��ьʝ(����jʶ���5Z٨����y��>�pl76�rz�_��7X"F�z&K�,	>��d��f�\ߡv �[�E#���������$R<�!���Uz�?��������{������W;�B,��ǌ޻J�nO"P���u�-K�YB��z2�Q����V��E����;F����j�9�G�3�H�Y�-���M�;�3~[BJ���o�dW��v0��L�Ѿ�Cߍ���H�t��L�O�n�6��Ԭ2~+Q�|l��G4�u颋.?�&����4�g�+�H��Ym#�i}-���d>�|�?p���`Ɉ�|������a� �4�1�K���k������U��a�G!�@����/:ߪ�~-i]�v,��N�ݹ�
���C�\	�\���(����JŐĳa0� ���H�Bٺk�<|� E��3n��~sf}V�/����2z�ɽl:��\[�tͥ+`��^6�ؿ@��/�]�'�����
���|����&�2k�v��.�E�UuN�� =��\����ݢq�|/��1�t���J��6�Ƴ�(��4�@u��]���u��0~���g�7?B�xm�:��?z�5�&��n��PBV)#S
'&���B��k�j���QB}��VU�b��FK�^B�n��<�����!d�w=�$0��O2�h����&%���8�u@��-��'���u��xZn�@xt��s��lha (���b�N�~��m���^p��!O�_i��-�x�p��ҖO糝���)4ۛ�z�r�Ɍ�rJq�u4�5�qoJ	�H���̏��R���75Z�(���0��*{�Gt==���t�+w��d������ݞ�J(�"�!�1�����g��@��b`�и(,���	��Nښ�.��,���yg�l.>�����c	�O������`?��J��{*�N�z̈́(�ꉎ���O؎hjP�e��7�o��b�NFs�aӸI�F��
�b_ϙ�����0�N���	w)��띬���r��(�OH�u$ƍ&Ptޘ ��6S �ʂս ���k���O���۹�z������ct���$v�����=g;e��T��g��S�F������q�oa
G�y/2��5��C��?��o��.��Ss�-仫y��;JYE�K%���� �CG�MF�%E���S���6�o���0[����/'B��ҽE��YjC^u�;�)VIs<A6�9���
t��$�{�/��1QV���\.�XP�N�5ф��>7���K��?�F�8B�`����`�A{��"˕���"��(���
�M���B����^���8�@ހ��K�yo�?�����n=Wy�_���j?�zXE��.%�h�*u>�Gj�T1�c���R��r;����,g���jYmwC]��Bx{L'��F�I�3�Α��C	���31ǧ�O"|Ĩ���n���Ê�X!^iʯ��׬�,.ު5U	�`c�Ą���)'"��H6GO��R:3v_Z4+��f�5ΣF��]
�)>`�A�,�;?3�.��v�
ĔՉ��8&�C>�6��*��h�m@�6�D
�ܽr�_ˠO�j��[��ށz�5��S���
�/�6#GƩ�t�m�*$�'������2Y����G#�{A�w`"
7��gsB=G�pWu�b�]?#U*]�I�_��F½/pHDPk:x0mIZL�v�r��_�pJ~���^or.�!h��LGr�Ui��7��Z���D�oQ.S/'ة/�m���5�*'!��mA[|���"�L�����[l�������g]�DX�5,�Pc�ǔKPҎ�yF���<�.�i?�N��'Wm^���Ρ����U�4:& �;O����/.]y�	�ʐ��k�Ű6��<a��{�"�{�xU�A"A;ۈH�0)�f��˥��	/>f������ȝ!�HG*f��2_u�^��Ϻ�뺩a,͏�5��.OE1�Q)byۈm���0���Hw\�Ee=�p�����]v�95޿� �M�u9�Z"�M��,c��C��B|ӻ�m<{����V^{�L�<����_9^���"B���
A[��m��a��~����dXOu��I������L��K��=_� /@�����;��C��1:%aob�և�x��]yj�|����UL�ڴ�ΟL��R�ExR%/D�w�a� �V�'S�ط9d��E4�����[\ݺ�]� �.xm���k�cH�6���w ��;ˋ��f1��q�`�dcAnc�����~�L����8+�������n>��bfWm�E�����1�9,�H��F�Ar�ⷒ�#/#�^�Wh�h�>���D�����"�����Z�z�����}��b�5��8���\c�X3���h9�^-�T�U�Ҥ}Ty	�.r�p�u���1K�w�϶����'b-�`�l�P#��+�vX��k)��\��F=D]*��7���AD�܋�;єmZs�R��?�G�����D��_�9^�Ytf��Ӊ9�R���k�#%��ՀW�Y�|⛇ �_��~`�Toq���i^ ��SЗ��k�o��z��7�L^]�n��և&91}��O�uɷ�m �f��y�o���/���0�DcKw�ew6��:��*Y��G����@\j�� ��k� � ;�,��j�c��JvY��y�g�LœVu��U�O������̠��r�7�0}o��OV��N�O}?M/�S�D�ޘ�����|��`xc�s����$�rd8�U��N���L���%\[�0Ba���z�u�*��ks����= =�;��*��fЭx��
��J�t�sg�����2P��791Ι��p�O�J�mJF�}�<C#�����������i������@|�ډ�	Ԍ��0d�S��3M7��)�g�vAy
���=�:�!�\����S�#Q�JXK7�{�k���K]s��֧*��@�5e����'�1H�h3��}�"�FC��;]6,譹�J�`|*��Q���š���\�OeQ���#W��s��u��1Y%:Se�ŏ��	[�l�f��(����uW�2}��3�(�}}�fS�:9���8���H84��(��|W�Y�s�90�
�9^v6Q���<A*6�6����*K��Dy�R�ۚ�
��[1P��ҽ�2b6J`��nH2R��}H�6���%�/(YY�}�Mk�ὠ��Uj#�T�05��P�n�܊�]���:��H���d�<�m�����נ��:����zy�z���a���zގӶ^Xc�A�>�������6��4�Ű�{(y�R.�u� �1�.0�ד��-a�A�r��KMLg�NE_eTf���s���ގ���q{[3/4�1N�]X�8Oh�a����9懷���>����Se�������`�@£�����b����&liD��I����V@��&����_�O�:�Ͼ�BilE��$d ��5Kn6�2��=흋,-�e�Cf�E��K���j���s�ld�Y��Z�{?��Ѹ�@���4z5�b֨�dsj�(e��ጯ2>��=6���[�%ܔ0��I��j�2>��շ�N��E`#m^4W�6�P���,�^G_yN)+"�
6�2��$����н[�M�D������.'8}/M�s	�-���f�v�����YR��D��K�6�*�[�K���I�C�����o��*��?z[�J	i[����ѳ"Lz�����0'��1�������[q(��8�؈O+a(�ϐ���@!�z�&��Rm�cf>���
���Ơx�����"�U"�1:�ZwB��斺���zN�vk�M��<d���a������*��9F0�΢����Aɣճ?��٣}&j9CQ�Ҍݕ/�i��="9RμHKo ;;���&^��?�2�	�|�gwg9�bʈ{F�z_���80S��	���'E��Z/io�]OKMO�ȥ�/�~Hy 6$)_�3�=�IИ{O�z��!DՆz�[����L_u�V��ƿ�������N�`f���|q�џ�<�a�,�&?y���8:�BA�b�p��@��8^.��E`�[�+S�o�u�@	�m/H�t\���<:�p���S�8Z��$���e�ܝ�?���7����ճ����y�/�Sz�RV�:���s�e��D��E2�B��b���7H�@{{��&�M,���-�w``��}��:�BV�C7�������鐂�vz��oڟ�4}����N����e�y���Q5��3h�c��h�k�^1)��4L�Favvna�C��IV}�����P�����Ap��Ũh�B�=�ueh��	{`2硓��Yem4�HW:ovˆ�˥���m��]|��~�ɤ<��JCv&''�i����$��P�\?�ʽ���T=O���xə8����4�ؗ!�C����Jy?t9�������h��
�ϵ����s��)�C�h�Z-X(H��cR�� Q��͆�l`x�@w�폆�T�����Px��;��"g������_	
&��!�� Nm��� BR���?��
A,ew.H譇ͥ>��?B�S�wG�� �ȃD�!���Q�x'�cAU�ǎ��6�3���p��P썩�Wam��+�մͻr�Y��X��޽�.�:�\��%�*�qZ��+k��$�B�oo�s�*��]���o�js�P�Pe��Ҥ䩼j�kM�E������Mvm<�Ї=/�&���8��I`�"�yOAxS�d��	ぶ"�+o��g���8FZ�ST�_X�~��/,a9-��<H����X�v.�9Q��%��b��e6�s�ͱ�Z�FJ�e�X\�MP��"��kw�TP����A��S>�mlgA"�de����*V|Yq?p!j Bᝧ��ɝ�t�6���:��������p�@�B���Bډ��-��S��ٖ_m�6��~��+���m ����%��z��#s���o�mZ3�3V��O\[�DN4�]<�={�ȘAN�P�D{��ve�'G��&���e����[J�w���a$N��μ)#�&i�ހ�|9L�M�����Zh�})�Ϯ���a\M�E��U&���DzP@���'6�\D��Q��YI˭�K��?�CG���]�&H=�m�p�MAG�V�G�(�Q�����uN�^��R�����$ϴ��Lr^��c��6�j����7�����R�$�$֛1�'���@�������1>���l�� �{OW�� ��n7���iB�ɅT�!����Xo��H;/����<9O!
ʕL�e;����
t�U��P�C�6.�~�{�����@�z�	)�Wg6�;����B��a�ȹN��nam��w���J����