��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ����������e_1��0Qԑ�@	�2p�E���,����9y!~��#jU��ާ����H�fu[�sp#����D��Bf�t]��A)*�e��J+:�"�$���8�����{} ��Sm��ش9�P�Zb�H�F����/3V��rrJ2~+9�@�=셽T$A�3d�t-��>#YᵶG}/����:o�2�݇�d����;;(�]=���R�^�%�~Q`5�>bEq]$l��=i����mWh�裈���xve�r�\�s"������H�9dQ|������ʎr��j�u�Ka����.D@`��w���bZ�}g�X��5��͚����*��]]ɉ��Q��P�����r.`�5��,�cc�3���2��sxf�/01¡�8�(s�yŷS�?o���i��C�X�x�dͩ��q�<嵫i!�$l�I���`\H��8�mr>S���Vh6V,��	L"���b��.�i
��!�L[n����i��,
QA��/����+(_0�>$ᇁ,Wɷ���k�`���4�7H��H�z{I��m.�	1[x��i�6!�h�q��}*��s=w^��N�Z�r`8؏�m�]��_�($��(~*�^�	R���p�g�1�e���!C�_��r�Y����G�!T����R@|Ǫ`��=�Щ����m4(}K�����a4�	y�9�t����2V��&|Qo1й�q��o��O�Y~>ُC�d���DlΔ��
W]"���u	1���\?k�c�@��%v�=��բ�|�[ސ���E��|iR�;��#T��P�v��.d�O�U��;��`�h��NDZcgw��/3�m8����_y�D����>�WD����;��;ʛO�0 ���-�������5�{�tu���^LE@͛��_�Q��!G6�)W�VJ=~�^��oq�s4�(6�A�����Dt��"s����c��`ʕT=�[�o��ysj��R�y�HTcI���Ԭ�F]��D�]������c@H�� �&�����[���Q��U�L�����%4�$:�t�ʽ�6���;�f[e,�`�G`1�b����/����%��1"�����.����ǈ�{�n�K��r0<� ߉q�EJ�e��>H��&2�wx{M�W\�2�O�OE"
Z��O�m�:��wƣUϱ,o���tBR�9�G�"x�V������#kOig��_rj[��˷H�4���Kз�ocu�{��qHa��B�Y�;��"3f��GM��̽�sO���M_~�.#N�:��:I�)Y���qP�L�N>���[ɉ���?�Y �nX3U�Y��̖�G�M�]�S��dW�RՇÅr]Zs�p5��<�@�j"V�p��2x~��=���)��$!:�6�Zl~/t�9]��+_ǆk��,E�Oz���5P]��p�I�N�6l��{*�oz\���1-Α�\���\�y�,��y�~�׿ڷ����zָ�r�w�#ؖLn@Ta��}�5v���o��9��F ث�j�5��S4u��$S��Vښ�Ĳ���b0>���⨻�������V��kxZȎ�ſ�ڵ�+� �,��� ��^4^T�v�Nc���p��Ky��U*��1�ǆ���=��\�~n�Δ �n�Oy��K��Ȳ�'г�K=m4y�x
�2�[�=�~� @/}U����O�O�r�ޕ�f�e���"6�������:�/Т��������U��f�!S_���T�V
������D��3����s�G�'����3��ǿ���P��c�4O:����6G?���A�h��{]���j��h���D1p~��;�k�$�SĿ��	���3���Zz���S%g(���IiC�jQ{d���l�U=KL�I�,YhM�k������.WCX# c�AdA�O���F��rNB��i܋��L���O�@)hة��0��/��\�Xͱ�ٴ�p�����sAH4�Ҭ��^C�ۇe4�s�W���@A���t��^I���>):��y ��F��c�s8����Nv�D��|�ȇ�?$�4�Dy,�����]y�LX/5� 6�U6��'��jL��h�,�Ѐ{�����2H�e�s���gpf�]��,���u����j�o�R?�#z��a�z��٤�s��HPpΕ�bo�/��p���n�ȥ���y_�IFXe��J��S�>�w'kH�U�b���0d]������[G�~��]W#�����_%�g�d��J|�Q�#�ɗ�"�ݻL8�1����r�.��(x����C�"~�h�'h���*Af�ɯn��晄c4���b3�ʣ���g��Ĥ�����Cx��
o�FpRQ���_N�j�Zȅ����,y�f6�!z�UD���/]���O�k*AeݎH|$,Z�YJ�_�!��g���Y��[�L#կ���u	:[�v�������j]iLO��`#���f�{�c1HJN�~;����!8'�9��NrqU�2}k����6�M\���*S�,�3��5r@��&�E���X���n.��$�
/���	���j��L����V�֡�71�'�M�s[��J����\=��b25�m�\o��ĮTS��A-d���R�*e�T��C�� ��}`@����ޚ��Ƭ1M	�t ���l�UB�D�����k��	�,����a���N���>����.�T��߳]I�{-���K��1�2��{��v58�$m�\J�	��S�=Y�z��Ie�[W�r��:��K'�U2�:�wd!��x����I��%F~p��E@,��몳�X$jE�Z� �3^��|�����t����}�����b�YБ#�܋�%3-7_���J�0�՛*��<�"�J[�������k�8Ԣc�.���(C�a3�I:HQ/p�|
�Dj�q�|�O�?f�v��<���a�6�m�����6�� ��k @)��$���V��'7c�ft�z�4mG��揃	q� <���NˑND(as�@���g�h>��R�~���	�Ѩ����c��_����n=��CD��/d��[��@v�JY�B"%;�*2L.�(�ȝ���m���#)����i���O88V��t��]}a�Sf��_/˙%�헌�%z�.%g�Oo�Rӭ�O+|���x�G��Z�M�Y��������i��v��V���:1?�j�VO&ve4�m3�I�3����}�~�Rr4~	�,Zc:��$�Z��������w&܆��ńAY��H���(Vy�;$�{�bΫ4�e�}�4�,AU�H�6��w�ًy�|Q?�0[� �'%��r�:r%���k�6bi����S�O2@"tU��NKV��[y[���5C&��-Z̄�$�'��:9�7r�����I�tΔ����DΎ �P�ݐu�p�1���h�A�M,�齒�䲇�$U��X�ݨ����g�B���i7��X{LEb�d�]uv�ȐL�a���#��𱕞#�L�V�(�ѯ�>�8<j��hz�%�����&G�sK˫m����/���rS7�Ȑm	o��ؙ�$�&E �����?8MG+�+���S����3e�k�#.x���L��iV4�A�E?��梚�U����٢[a���TD�9Ix;6���ӧ�)�w��z8r��W�(�T*��;���k���-��ͽ�1��,;ޔ��HH�J��P�:���фN��l~�z6���a"6�6�Ja'8���{Æ���W*�y��M�!"�)�R�͟N�!�uܾB�U-�}��%���|����O<�}E�-�����:K���Pg��~f���.����x,��KM���ޥ���Д&�)*L�k�s G{
������7o��+�aeyz2Z�l�&�~E���颷+����O����!Y�:�/��y���&F�i!b��ד��Q�D�s�b��`N�� Qp���|���~,��������k��a��ª���[^�BxhS�D����_L5�Ҍ���u�\j	��'��}\�%��m�x KL6h�7M��U/s�
��7^�O^e��O*ߒ���;mr&#h��B'q��� RN'��\`�RN��g
[���97�si,�jv���L&�$��u�2�nW��6������UV��I�H�z�2I>.�c��Um�]ց� �#B�=���=��1QY�z�udMG��<�T�O\q>����+�ޗ)`8���f��X|6U8���e\tTd����(E#�HDTVR�9�A?j������N ��d�1�-4Q�u�*���1�
��'�'P��`�e�	�/��ҥ3�����zvf�LQ叅�ظ���Z��VYu���]֍��m������
�.�O���g�*�S���[)2t3Q79;3�v.7�[ȏ����Q켆���,<��Pk6����v@T�yz
;{��ָ#���=�/�6ƉcԼ!:��P�JC��J�p�ÎL[�IT���'�^5^�g�w�Crj��A(��u�]�T<4�6���ʕ�L8ߍ}��I��7䈋�٦�~�Bq�
m����
�>�XSyT`О������
���s����l�l��%2�O,���hm���<	N jc?jA�t�,B�D-;iv�~�B���3^�\~�x�N����f#�?�i>����������9�!�����!�?"m��J���`=��𵮘N�Az��^�:��͕_��[�ZBR��٦-��^U��xE�l>je�y���pN��窶8��ͩ�O7\U��>�I�}[�����B�D|m4��ƹ<�!f�Or.gڌ���~���X��-��E�:�tU��vĵ�y��X���ʼ�����J���(d��'����?�TB~S)؉d�T��d�GC7��1A�P����G�i�"�,g�kLξF�6a��ț%��("�q�[���o�wb:��(�&�|a��b��lSu�7���eN)=��@
eO�	u�W{�GV���q�^��!��l��ۆQ	F�O� �t����qhauC
�I���˜�@�âA��ف�{.����7�II������ݪV�W�>�|\&�d����]�}�!q�Ô��#�]
w�9�P��N+Ogl�d�0>�*?��.cc�V�I�yO�ypS3�6���RH!�;~]8�c�� ˛8+F?��`i��TD b�~xaLb���>�����w��׌?()��:3D���RD�K�E�ꔎ�|��'.�9���3��(�TQU��b��s6�^���Ht���Tan�n7�`�'��tǤ|���������I�o��R��9�e6`j�K���}*�^η��ݒ^w��x:A�'�q��Ƕz{�ɭ��O[d�]�H(FO#h��/��J�mn�^�����Я�I�w�����js�ݘێ�+	7�x('�z;~�E������E��~��	+?ho�
'���S�%�1$���*�v����d/����^��RXy���8)��sٗWn�hU��uc�wsojM�ȵ��`+І�\��wH��H�̝4��=�����*P/�䒑���pϹt�t�f��2X���wj�d�J��B"��h�xt��6��;�i ]�<�D)�C��W�0��/�j<E������ �A�2���zY�v�6�e~���8�d(�ꄋ	�h�v���Dh�c= �)C�Ȃr�de�U�6�s��Q�
֝��l�oV����� �)��i�l�@�O�L"��+z�v����4l�dU�r�51����F��PX�4��S�M����W�� �ו��ah*E���?q��Ae��5?��΅�w,�?�J,!�f���:���V�Ŧ��W|�i"��.�E��E�t�%�蟨Ϟ1�Z�J}ܖ��5��ﱐ������YF���V�֖"�+�����XGw���態�� �����D݂p�-�a]s�Ѹ�����A� ܧ��ލ($G=e�;���D�����[Ir�JR�,w�Em�Xx�#��@��ة��[�s���j�ɣu�.�Q{�Rn���ǜ}�᦯7���:���t��ޔNˬ�Ħ��@�{��� ~���w��z1�v	��6I��E����tIȽ0���c�P�ퟖ��saj�ƅ�Vu88&W�$�=�,�0��N�a�|^H7՜u�49��
1��P%��,
5c������>܈RRN���m�k!}�<������r?��3�v�k�w]�	������b;\��l���%�{!�����-?:������� x^����fm����,nY�N���=�gʉ�5}09ՕE���~�5�[�y_�ZE#�D��t��W�s�e�s�㊱�`�l_�0a��mr����M��!w	x�k<?V"����W������a�/|�{�b���RqA�/� �Oy��/a&�����%c�]B�og��2��ܪ<2�����$�����$E䛝D�t�[�F���K�~{�^�G��꓈j�z�|�Ed'��.���jue�����-�:�gi�GR=sD�m�@����gآ���O$�A���.�H�]n�4��0�0����؛7?�����(�1�G�8U/ǘ�M��.���u&��@m��
��!�Q�iD���ڙ���w����4����i_��� ���֕혹��4g*VϾ�AqG�p��i�$2�g�J����ڇ��n$U�b�;%U����t4w33�v�"�LE�p�0\�{�������~2qN�b��}T�#%��G�=v�v����4�ɘ�A��?+ӻ�4V�)Ԥ����A���* ��R{���K�N���3��ш�6�����Y�f��^<K���fG#��_S���#9��]������]�3!�	m� ��{V��J��rȢ@t����Ȉ8���Tզ�H����br����ӡ�ho9�U�Ҳj=/�]n凋�����.����"��X:�s��}��q1�� eI:U��' �H��aU�B��uoG]O+&�߼D��x��x��}�]��%��ɨ��a{XzFƓ#�]a
�x��}�z�90iO���8������(�|.�Dc��8xzU��[�&ƌb,�;�Ǣ�SP剨� J
[�3���r�Ao��A��c���x�>	cښ�0��}�����崗������D�6`�kU"��ŭ<W��=. �Uy�?梍�%稻�"e1����B�B�,��:v�)T)
���r˺��X>���V�F�h�*��!�t��4�Cb�{�"p�����,j@��s�U�ڑ����Ew*��h1�T
�q茪��v.(�g-?��j�T!��*����V{��o��J,5E�H�G��E�'��Vn��ط0\"�g�#�!��8�I$Ɔ}����HX�Y��ܯLD�[�@����|���+�~�I""J��I=��Z��-㹏;��vQyyU�K���wE㔔���e0��ut�����g�ɜ�l�'���Y8�0�	%��g"Q�w�u��� ��Su��h�c!Gp���rˠ���}ɭ԰ⓑɜ�st�^⭄�U�\��̦���d��,����l�8���BR���0�"�T��7�0����'���J��{B���q�,�XŪ�R{]eM�Ƹ�t��1%�1}��C�s� ���ia>�f�Ls��=Xliv+;����Ah���5U�²�$��ȡ+@'�����p�vK��\*�WH�U��@����(ŭL��Ѝ�T�j�[Җ&�k�k~M7���  L΂���̅�0��\g��{���
LXf��fR�ʕp�*�9���I���y7��R@G��/6���A��̍������|2C2n�_!��?�!�{]��
(Vuk�_Fh*=���mn�.�)��i���O����X����(Q�`*%Q����ΚqKkF+�)7|Q�%��b�	�y�([j//�<�~�O@vc\��p�Nżzt��v�^�Q0�����̎
��>s�>��t�{�q����v�Y��g�:z�		D�e���Y�ͱ�;�|߄��