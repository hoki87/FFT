��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E�����>_�.�*�(e�{��?�4���I�x�Z��iWڲ��~&X4��-k��l���h����[��J>�B��:6��Hn9+}���xUU�s眓TM��Vm.�#�/cm.J�߉��UDX�ةo�!ժ�]>���>|S��Z�L*�EM ]���JXmk��J[V0�A��Aǧk"�\�����L=���7x�jt��Qc>�Sv,Q;���h�(�kHt�Oʍyh3p�0�����t�"��͛;<��'�޲S	[�^�E
����;	*��q<�[�`��{��LTPW��ic@�Y�Rxb��hI���w�7O��n�f0�E�m!��l\��6>��_�Z�5m:5>���C�p��P)�<\�.�|�PC��d���3����f�4�p y|M����h4�)R:B�b��#r��iH�t ���T���>��)C��+�$kz9n�֨&��~�����4P��H�\�Gށ��#P�fq�f!�W"y��Ӌ�眪|i6/b'_�m� �\��؅4%v��omp�i�]����	ԯ�P�.�pK���;,��������pSj�'�)��l���Z�2�1�9].��ۢ�u�����Zh�SI�W�D-Im��fՙ5���H��xE�*�vYm�kEb��<3q$:���{�vyN�����QG}�G})8}�����zd2�Md-�q�Qz��?�t7h}8�8ID��9dOZ�U�*Q̰I��2��PS,�O��퀿�C���-�YF�g=��W���[��gD�w`g���n,s1��ܨ���2W�`F
�D�c��iW�.�W#ځ���N��R 6�-�8��.������2�y�H6R؝#�v�����s&*A��g�Ie�Y0.[��Q���%A����X�G8 �e(o���Wu���-*-�Cm���c�S<T��<�@�+H����K �y���Usc��akr-���X/`�2��/[�:����Sڍq-�8��8��q��C=B���!59�BF("����C�H��y�+D�WA�d��L_ʔ<;8x����Z�-��ek��{N��ݤY�;�Ý�/�Z���uk��v���=j��kѰRUe�k��e7-�[�/δ�:��L�r"��E�Pv�5�Bt깽��M��C��g�9�!�u�sP��	g�BD�ʮ�R�וB�p�"A�e�kK���!whɶ�����E#��?�:&��IY��8�@͊.'��[������gȄ�8�$�d\��K�j/2>r��iӐ�Xm��ؚf�:�,�u��6��=&��CV�5|6ɐ^�BF�����Xw>�W9S��\N��9A��F��[���cF���H���7܀U6�uܽ�D�ݐw5��2�9��t�(pO��!��E��]�k��kA��;�'xUJŌ���HA6wq����GVu�榚��E�ϫ���\G6��.���i�~}�9�są7yҁ4���a��%Y�(�=6Am)n�Z��r�V�rB�R�Ǎq����4�6B~��Q�YOWj��M�o��
G��K����l�"��)�B��<��DC���?����?���v��=`^oU/B���;:�����֍��rX��J ;�ۯ�9�ww��C�h�b"X�IýrU�L�в����V��PL�����0֜�jl�m��;z,o�@�?.�������u��Dn���B�z�(��(aeY���Un�ҩ��;rb�����G��U)��TY�Y(N�y��x���7�8������s �^J�FI�.xDs4 �X&�R��,�2��G�y'��� ��т$}�pfO���R���K��������4�Oз#ϔƒl5S3tf�Q��?�����ui�[���P���h7���Qq�ǲ���m��e5�l
�z53p��W6��g��=��爆�����VBxVE�<�b��o���{��"%��^DBľ�9gͶb{,%,�Wx���i��L�ņ[[�
*��9l��؟/ǦoM=Wnx�_sf��LX#(<�2&޲ ��|d�mqn�M���\ާ=Ta���e<	q&t���I��O�-=��?n�CZ3�WdJ`T;MSwڲ����np�0yh���w��qB���#���&J�1��!�13�](�'$_�f7y��
)>	�FͺG��J�R]�W�~�6��T̜Y㠱�}^�(׾��Ħu�-��~h�ă�����T��s���uJ�7�J�5��~�1ɱQ2��*@-9�lOkHl� ��#���9�;�',H���W3=�G;�E�Y�цo��hNmya$�G�4t������"\����I��D�,�j��0�D?-�07/T�33'����O���joW~���I�{IN`����Ϟ�t
a���wiťZI�ZJ�tv��$@�I���U-'��3ݼ<�d��a��n���z�YC-����s��@Aǃ�W�-0�:�5��ƕ�^��������2���u����� �64�^/�K�b"ܥ���(�畛"�X����ȩ�e���P�\�D�&ݑ�P�	�M��ug�©y؉m-^�sCǏ��6�բ��t�ߛ'd���r�K�A�魔-�۟p�JYrI>�޲�UF-F�D#��y�=�nl�k��������|A�5]i��ֹ����2`
:���&�ͭ�){n��#���Z[����}�v���s�������B���JAWưK��O �=-�0��s�+�
�D��@�[��f�-i͟�<Tʖ�-ƕ�^}�|�v#)���T[u`o]V�>Nz��7T/a���lT�������G�F����X��J��=������H2&(x.�Ų��!'KVq֨�?�pp2��[|0�2*H7�>+���@��^�'w_0�8U�:i�<�bʳ���<F#+Й9t����v��z��������Yn���P4t3�L���;D�� �`��mJ?����b�l��2",$t�6ǝ���zj聣1����g��V���(#���AzoV_1�	&�N>�2oBk�� ;mg�f�{�C�2/R����lI�&�M����S��� N��ՠQv�2�y&�8�����u�2��DY�VcUL���$�v8�2�}�G��&��/�$A��w5���8+^����fS'�솫e�SW��'����j��H�v���'��\�3���[���B�;5���37aH�[s��rp��S��F�ϳMl=�^����=pbM�T �/��,I���Xpf��;~��S��bI1�)���������'F� ��L���ӚuլL�~U~]�v�eQB�~�~6l^Dw:}��_?�U%����8{����.����娉UN��Un�>-E��6-�����V����w�����Μs���}�~v�p��h���X��P����V5�c�m"�/+6
[���T��CB��i�6�w���ywW�a�0s '���ܯ���ћ�/^���{q����*N|%��y!����\���en!�1�K5��Z,�p��1�X�ӄr!ZE�������#Z�I�s�.N֪i.��O˺� ���G�Nt:d�O�
c��n�>�ABX�s�����Wa	����Y��r%�	i�+�Jo��v�T���}a,t6X2HÃ7E���	�)g�Mt����e�X���/�<[��A�A��tq�Re��	
<Ζ�C)���?d}�|�DJ�QF�h)UQc���јW~��ra�/-��ޓr=H ��Z�c�? fȳ��jJ҇ՔL*%�lƈ���+*�KI4N��*�wlv�� T����)���ւɞRJ�����Rq�Ic����@0��Q3t�l��V������c?���7'`Yxn�.�@�XX��ռO�Սd�Nm�Q6���e�G2!��<q�[P-�=�՗R��V�����&��=����u]A�/Ŀ��4sK��SH�y�O���,�)��U�p��`U|�V�����7�8�(�
�r���+#0����a�+<�<��H�̱�.�9��3��v�
�x*��w.<E#���9R��S���.�w��tĹa�5z�����M��Q8]��n������:�c���K��	���O���d�Ԍ"���̄>v�p���~T_4�mD#t�)J*)��S�N���X���o���(�
(?��w/��G��ZS�y㻟
�R�#6�� GR��A� n�3�W�i�#�bȳ�;S�߯ =���j(`F)�4�,YǪ�p�ԕ��)x|�y%����t��ӛ	7�z�������|E��&Q�o��r�ޥM#v�S>��ڗ��Y����Z���Nɬ�:��#��S,�.��O�ah�&>9�0?�%ZsMp�ٟ��G�8<n����"��W�-����Y)R�Ӯ���'�3S��<� '
4��҈�;�H����i&$;�'�������iֺn�VW�m<:���� �mg�F9����9����9����y�s�t,�5w'�W5<��ҷ��m�p?{I��q}��ѻG蘩L�Ք��?��0pG�`/�԰���>�zYhKS�k���?0�;�X�d��|�mM<e�h:G��ⶻe��K���.G:5�pQ��Y�MZY�?t�"��\ ��E���sэߎ�\^����g�tRQ>�E��e�j�N��ؠ�n�\�;J���ա)���5F$ۗ,cb��:�kb��'�oI�����s=r�	(�V�m���(k1f�X��	M��9�S�S5�F�Ga�������l�?U�����<{�%�x!Q�ґ�P�`�W^��ƴ�e��\})�G3��)1�\��
��ĺ���u+[�\eC)�^ɨyØѝKHc�C�A��s!Uڶ��#؉ s:/K���JŦ?XB�y?���S	���t)+C U
0�4{�NR�3A����8C���)V�����N)�TbԵ���b�r�8��^3'�d�2	z%��������b&�,�NZi3^֖�B�	Aq��E����v�A��v�*����v�-��vR d�	1Z)�l� ʼ��Y��#��Su�v�E����T#�{�逊�J�.��]��h��{_���_j~�u��[�i��D<&���,�g,I�����" ��0ƶ�b��a��C6��Rg�W�P���u9ԫE�i�ѹۃ-T�#(r���?��ƹ-�J9��m���fC��G.��4f�Emm����3b�ӁGOe��(��!��^����-�����=�M^LR�g�-�,��O��&����B&ۛt�4�Pj�e��IF��g�xdvqY���G�m8؋F�Z��a��v
O��kk�z�a ��窒./I^��p���ā-�/$�T��G���G��Dsz�j�v��wv |/p�q�';�:�ɂ��˵�Wi�����,:�����s(��$��-[���}a>����.W�E�Dw�`�]��V$�gu5B�����r�SZ�%f��u�죣J`���	�y@��*�8����ǭ)�D����xA������Xd�-и�O���YĈ4�c`@p�$P2�O6�M���x^��>g�$*[� �z^I��4ܒ�\S�:?����	��iN�v
i����o\h(��ݠ~�y���<��k4�&x��r�/�0�;�=��G�J��1f��rsR��I~V������<�H��� �2�?�����/Qp{��'D��ėU����t��-5�V�vǣ��!A���';�-��ͼ��w�gd�ډ:°d��l��M��Г�0($�B�k-�|�Vb���6�������H: �����-����t��V��%D�6�a3�ݸG!3/��̧?����削_S���q	e�k.D�E�]R�����1�2L�j���f؊����N��M�����z؝kk�I(�^R�6�z�]IoG�i>�����1���4��|Mig�����)��"\�{V��0�'|�l��lF�h :��j��.aϑ�6��&�:�K
V`���qqNDb��YE�q��eqX[CC��X���0�
tAc�ީW��|z��s�[��"��AH� ⍁Dg��ߜ+ᵨ������rin�G',>{�Pǲ�!�� b�a������Y3`$VVR�����	��8+�;��6�mH-��FX8�k�'xN�}�aθ8���,c�Z��nj݇K���z�_'`7m� q<\�;��G A'�����u������;�<;�F����K�����6�¬��1���e�v _�&�!���3��0�=��=xo���p�M��Λ��lݺ�7��9"��$��&-y
w�@3^}�e�&�,5V�!�;ׯ����ێ*P`.����9D��y*LD�L��C�+W��ov���#�+8ұ
����1[M��G��w��DF�P��7�m������ָ�ݩ����lhf��{�&$ '��6F$?���?�.�(�i4vfg��7�Ў�4��驕��Zڒ�Wq7����K%�ee�w(���
���!���K�a�ë�d�vμ>�����t��A>��|����	$w<>�M������Sb�IA�6���d��	�q�4Ljtw�3Qʡw�-�5��; 2�	�(�"�1�4��N�����ܓCT�|���_�BӢ�J��z	ؐ�˙PrV�Z{s����h�������u鞠�T�Qv5Y���>.o�P�� ��#S�,��ҩ]Y��li����y��%�A0����Wg����<�E�r���cX�R)*$H�o�z	���B���0�.{���QL��Qi����%"�ҵ'iN�Y$A(C|*1���%��)/y�� m�N�7�����N��<��Sw9ޟu�"tVNh׺��f��G�|A����"���~�-�����༶�s��V`�������7�6��w�sږ��@Uu��~Xjl��3II^y��3m�*�`(Y5ѷf�B˫��u/c2\��[n�����#x�,o�%:�.��vcpK��G������� oq�B���6��?_2�x9��P����d�	t���%L�O�Zhh�W�xD��J1Ec�-+Z�#Y����Ji߆!�� ����UVy��~�Q=d`�F��B��v����t-9trn�'*�YH$�H8M��~�9�W�g[t؍��D��F K���Y�~���GXD��n��D�M͖9Z�5$��9ĳUO�>�u5�*�����l���Yh��w�-敠�@�N���e��tK���������ݦY��6���}&oi=�EQ{���	��>9��ьw�Ԋ�+C�մ���bEGN�	�݂�����Ag�����R+�G�f��G��Y���ȟ��󹡇�q�>en����&��߱�!g}#u��Y\u�0>��6��P�����W��^3���cE*�߹s6A##����
_.�9��5H�Ӫ���v�>��T�a Y�K�Q��E����XZ��5�I5\e��$E .Vb\V���0S&yk�D&	�r��Y.�Qn,��/��}�33�_56�1���1&�i���q5/�r#@П�h�y�99�HbE��W�F�U���u��6��c����"\M�O%�����.��:����j�T�v��K���S�Ѭ��[46�N�`;����b��pR~�M�ƍ�O��ӌ>6���eE]U�/��׸">�d��q�{��v�����6���v��;�ZMT�!�-MZ�lk���^g�,�*2P��{��q�}zX��?h߉�\Q{*%��ڲ��"e{ײ:]�Ax>?�Y2,A�U�r��y�M��f^�3r���LBpa��vW�)@�7��ir{A0���e3�]:c���s�%�(_��g��?`E�A�wZ�����H�ol�'l.��b|�큻�	N�IuF��{>_����]N�h���U��.L��m:Xv@�zb�Y_� ��?iUt��!��%���,�S��{@y)��~Wʧ��(r�+ŋ/9yܞ�ۿ�j	�-��	؁`�cؤ7�ǵnf�F��F��"�&ǸB�2%T�/��;m�)��b����]M����ʫ~�MEs�JTt�h�~1����vLOX�!y
��6�l�*�4cOɳ3��B�e��(gdV���pf�Y������K��>;��`R�me�E 8k�:���2c�c+���2�a�`v8i�#��[�C1�U�8��ݷ��u�F_��+uO~Af�ʑ�@��!��D��B+�Q��l��S��79>�9[lv(X)ht�AC����E(J%0�k��P�?�H�pw�t1�%��a�pX@�u�7x˼�#��e>��AVB*_WlVi���-��v��^Qn(
)�
ߋ���A����-��Mu$bg� G���0܌�Q/Oi������I;���N�޵���_^�"���2�/��0���7v�
  L���mW05�NNb�u�f��ĺ�#<.9��V��޳�Η�K�~�)!�˂R��|�;YP�O�8j0kh��$DQ�����wׁ`��u���B��z�fڢ���$i>�����0;�b;�J	��VT"��l+ɇ��^-�����r���M��^���N8���ӛ��:.��M�=�4L�R����@�U����u@V�sc1�d�4kB�/&�W������Hwe����ǟ���)�DM(#.�2�ů�QA9�MJ����Q�-˹�e������{@���j��t5��c:���Ԭc(���h�T�����=f!C��f��T��gj{>RK�b��kB�v (��w�Dv�m��������B�ڱţ�pT� x�k�����f?h�~=Q��q��J��QD��l"���$4�-�S�)��5��T|��c��b���}����Oi�`�R���sQ+�}��[������t�"��y��6x���-�����0���$ۄs��B�lw"��˚k3=N��l�a�ë�g�2����
.�Ā��0Q�,��!�g^�N.�c�; �w-�j���#�'[G�f��&l
�GxG�#*�E�����]�&ta8*�m/�b*�L^{��q��B��J�/S��e[:4�B�)�#�ERo1��Ʃ69�C�5�$7r�6� �,�\^K�Z]<_�],�ݳ����H���2�������E��֧����$�~*��+��ݭj�C�::�U��LNy�x[x�5:&�z��e��'�wθtJV2��#��X6����S�_�'V}��@�� �E� Q����hc�
��
�Eu"d�B���<`��6�����
V��+
.b~�[�����u��<�w�Ӕ�,lJ���@����z�������c$Q��8Gh�V�'0��1�F�L��bs(k�W"o�[/���D@��	H�v=�Q�H��P
�֍JE,�W���D�{�����KdZ��8CA���Bh�����E��'v�1��Jq�����?��F�Y�\�_�&�����'[�cQ@�?��-��mu�x�����'�	=��-�Y����.ȕ|��n�V�uE�="��L|���2���n�F�-���^����=qP�9w�Io�q  ��w�o�l.����A�,<��cҒ�%�5wp���4���[�&|L��m`w�ܲ�����â�z��6�򬌻�ō�%d���\���~�M_R&�Q��kM�^��Sm4ƣD},l��lX�z�d����T�n�J2��Ϋ��Z�_�vh��؉l�=\��)z�����)�@ չi�ÒĊ=�M�c��h��-��^ہi�>>���z�R�Di���a�I�a%�3_4�JF!# ����|֗�Q1�#���=��X����Κ<=ض����<'�J@��,�pZ�FSL� ��P|3��7�­�߸I��hM��e���x�Ě� ��\^
��M��F�$K�)؊E����6f�?��S�����I5ϥ�F������v�\د.��Q6�;�̘$�%��i�a^$��Sے�ɠb�m5��I��=#��t����Q�f�8*�p'��I�M�J0Yh�A�47S�\�Cl��	�)��N��+A�̶��� �����T_�:MM�<{���Y���qp�x:��{�(���x����%{�uH �Hc�9`P�~L�pɏDЉ7qCQD��� �H5��ξ�� �+<��^ؾ���g�,�mx�Y���QA��<��ئ�'d@݀�<�=d��v��DpP����⽢���?���^	�GY�t"XV��y�H=7���I%���k�UY_���A�R١p5�� ����5���#�OJ� �m{Mx�7��X�oY�a��|�9圤��:Ed�fp����p�lETS�*y��i�K��~�>��h����!����^Ǻs��8�́=#�aE�T�Bg�5tǶ�>1��v�����$����ɢ���[=0R�o��ݰ�7���t��xy�Z�إW9��U5�[q6��������ӎ�d+>�~D�!�f%_��v���A�U->>�{�Yjj3�4+7�}u��[�d��\�̲�����Ǝ&���R$��c���� ���!��K��\�Y��>�7\�I�S��B��_�f�œ�.�!����ġg�)����0
b� jr�q��_���m0�F���I��x؅�w�$0+6�@AU:CEak�Q�~km�_e�9�+yL	�ّi��JHF�U�\J�B�z}�#xX�e�1��9/1����z�������}�>�B�����<��#�*��;� ��S�����+Gl���� !���1p��	%\~«��C�L*���ڭ��4e��V�>Ԓ9�?��n&H[����,���ް����(ۯ�Ktc���y8��oK��i�C����	�&��Ƚ�ЬDM̽o1n����`��%G�� S�ﻤN�x9�.O�p��c�UU/���÷�뾤�ۙ�u|ξ��H���fJ�J
�f=�%TL���3�B� �{,�3��BH�`�«��ݦ���D�VM>X	��P5�h�,=�Ы�EoY00PKm}v� ~�o�i�Xl�)F��;�y�o�t=���J���%�����;���]�=�x�P~���ɷ!c��#PO	<�#����� �N��%\����n�1�@f6�6����(�ĻT�5n���;��|w�y���B��1-��Y>DI%Z;��MM���JK���:I�މb�~�>�1���G���n��g,�L�Y�`�[v�d��D��(~HS�4�f�0�	D	@�8�<ݾ3�.9:�[`w�1�&�L��h��i~����-���Se���NEhR&��N�����%	�[�\)����;�Tʆ򆫺iz�n��y�7�D�V��q�z�H�d~��8���G��B�vVW�I����H�$I�O�.ʽ����Ⱦ�#�ao����P���_-��K	X��~M��'�������ʊ|�"[o��,4YB�M�τ��Saҕz�O_�e�gw���^���p�	�<�R:��V����zg琊���yp�����aC)�W4 ��:��LFv$5[џ�ȰgJ��M���j�E(Q<}�c׌���tl�3��X��kQKaQ4�/ ā�u/�N�5G;4'sQi�r��n^������胠}8묇&F�K�<Xk�?��Ln�ؓ�Nj
� �C
"�	bNb�lc03�bP�����}JZ��XT�p"W1�/�2Y92n����'���A�b
'q}��b�c]��t<������:]08�X��.��&b&zi���ͼCr�U�Rs�+�'Y��V.��K-b�#�ZQ�m�(@��-����+ۺ��[W���y�6��Ǽ��G�d���WIа���UX��8����?�~����	DC+�L$�M��`kn�3$Ej��I+���*�����9<�s-�Rs�wA/�������M����vx��� ��E�1��m�7*�UZL�XD����+��f�RZ��=��� �D|���aGa$}��0|�5�V� �������]�1ZF�u�si3=k���p����Ķ���v#��G
�Kn�-��G�S�R ��\iI�%]o��j	V��>�{�Cc�sB9'/���Tj
rX�_�V�2I�V ��ңqP�D��`.���I�h7�;_a�Y;����꩸�͓IO�����~#+~r�Nn�0�I�޹�jaK|c'��&(k��f39��~Ϙ��s����`O�Ia4Krj�!��ݫ�Y/��ܢ�˥�-O���K�~L?H%��juOq�� ���Ad�x��/��ެ�Q�F���h8��0�� �ɓ���X��(6 �1�c�Z_�?.$hI?J�\�����ڿ�(��:㖈'��:��9����)���#:�s��8*��('m���k"���8�|N��"��jx��һm9���Ϥ�˿�� �:ԎP��fSڮe���ڞ��@�WA3���0��=�.m�3i�! ��2��D�,-���� �؇�S��K���5�� ���7��"��4��20�#aD�<]�i1���Ԏ�;B���9�v��O-�h[8E�66A8���|�F��s������~��
LY���`\¦)�j8�+�Ql{4�O����T�r< ������Z:*�*Ͷ/]�d��wI�U��;�ЃyZ	����$E��N�XR��~ƈ�����<���m�Ln�&�m���8��J�T����ʯ}p �& �r����m��9i�5�S"�����b� �m�U��%�o7A�0?�U�</u�~�ܧ�	�F���|�\�L8(m^��Q�Vl�K9pյ�P�XxOq��s_`ۄ����N�^�^
�eTD<��'_J���x�cHgׯ�I���U�ȸ��W�,_j6����[�H����ۤx�	�񳺭[�-/U�Z�6v1$d����a�0D��:�:�����o��j��Y�Xyµ�%���{e�7�e\R�r1 @�����Y����IS��L���e��c�+�g��h���m��`?�*��`"�ֹ�n:���p��Ez�#� 0�4�G������3^>��Q��R��W�P�j���8����-6I��Q���Xj�!2��g���a�� ���:��覱����G���<���	/Ҟ���(IV7( ��Ԕ_Uc����).
Y����*pWfvhw�B���/ݨ�mqr� >���*����7Wo_�a��+�\���U��9[K���O;66L�?�5sɡə��Y�o�Z��j��6$�����p^��u9��0[퉛}CLZG������iI���y����=�ІK_n~�a�X�a�;�,Q�ALoǂ��ܤ�<Z�-�[<�U�
��,����A�^��A��:�_��ҔD6���>����%����H��`N5�Rڦ����E7��n�ɗ�gU�J����ö��˽J�~�C:i��{x0�J���W;��½���y�0.�J���m����!|C-g��$`��w1�/��D���ir����t-他�=Gn��;6OvM���4�H}s�R�8Yqڟtfmyc.�	��2��mG��&"S+W�5�.��t8)��-��o��t�^<\��1 t4W"&FM��h! ��Śơ�f�f�|G�du��,:#�m�c�J�e����:O!nW�P��~��f�Zə׳/
�e�4�!c��Nɛ+)���7nkwh�0���o�A�7�@=}���kX���L+�S�}̫[�`F{t�#�=�"E�_�5�f�]�N!j��!�R�e�����7"�G�4y���Zy,�SV��F;*�Q��x��P��U���<�3��w4d��<�t�%ic�]��H/��g�*�rz��M��gy�A���<��<n� ������}#�$���s �+�6h�:혮�L�W�z�Re*�DU���o�o�����[��e&b�� 2@����AކM2���$))¤��d4�Nz ��6#;D݂h ����n��HO����1����z[7M�"3����Z������ t�2Xor�%˸�c�.�G�= V�~F��dõg9w
zj�������8���� ��-n���ލ}�F"�^YQV���1��rw<櫖�<�?}��9 �g]����*�̐fE�(�;�� y�A�q�t� OeA�n��;�� OA��M�1�.���3~����Wa����]�a�ݿ��W���p�W�ٹu0����..�yk��f$/�Ɍ������r�t�J����%�xmh��ө���
m�&?�K��� �Q���)O��}��ؑ�? a�IO�*jVY����<�OK�.��aѹp����q|m� ^Ȯ~�L%�¿�w�<���/�&0��f���I0��fu_�j�7B�m�yY��]��,���H���l�}��<G;���S�89�/e
�#}���o82=�M͠�d�M����].�2�6Fx��붌X�c�W	�(9_�`���������k3 LZ�M&c �/�k����NsE�5둧��y������"J��ì�ێ����B�/#PJ�ve�M��;F�6�?�^k�Ff	\��L{=�t�(�4�Q���Dɿ�$�-k��]}m�ɒzQ1��j��6/�\�����F��nG.f�+aBs�#O�LrCb��
�_�Q^ki���l<=HVW�:w`B����2!!~��#�ս*��<>�k�Ķ�C����Ҙ
;>yn����n�B�}�j'�A�����q�	�4�ƙ' ��%�ϥ�%�h�FAu!�L�l��C섴���[ ��v�\��e�C�"�G�L[���������@x�h9��!�*Ԡ�?Ϣ�s�5[V7�Ӊ���0U���e����%�b�S9�a�� $�y�Fb�$KNi>�����<��_�����jA[��<� ;!^�? �A���v�a΂���'�$3�;Le`�䂍�`+&��9���p�2�V�OG�`��k�$�r���x,� ��#B����3g3�����ơлt-�c*9n�s6����@�b���ª�\���ǆS���b����Fl���i	G>�M=�_j[�Q�-:�g#�R�V�%��[�ӈ׵6O%}O�Ⱥ΅CJmH��Ԅ��$�!�~�F�*�_m�pA�E�2�(� ����K7�o�� �b��	%m���^Ԫs�����3ޅrh
"�*.��O�׽Գ��M�=M�X��{E��3zhQL���T @�@K�z�)���u�Z?�(O�9�T9F/ߟ�~�U�tq4����]@�����+J8)��쯪k41����6'On}S&�����x�R^v5G3v�1��e��S���%�"��iC9`��5d\=��uX��`Ս��I��A/&�kg��`�+	�N�"�� ��c����N:֐b�'��9n��0/�ݳ~6+�k��ɴmn#��^��c��H��\����T��Yv���i�,����	kdW���%��w��y��Q��|1��J����[�bgj_�J�`J����~&�	=ŋ��]�7�i:f�.�%?`0Ի^�Yh��P���q:@&���s^�fo�������(�Sصzz#�F/��M��Ò��t�������`�Sn���@UU�g���7\�U[g{� ��K���W;�a8��\��֦�W�N��R�0�H��� }@�jbQ��;�$��x����
I3�d�c�K�1ꫠ�N蹈
˵�����5|��F/h}#{��"����(woWt�6��R�ʄqh8�z�6=%����z�O���
��R��95���o�Ocm2�&%+e"o�үݼmq���p���'Ԝ�v9�3H�!Z����EF��]X�
9��#�{�?P�G���T_����p�Q=t�(>�����!�>����e �(ǧ.���Z������-ݰ�u��)&��{�6KMWuSb��	5Z?�� �7��a�0�a�^�����Q��Y�Zˤ6���pu�e͊��m5��ƙ��*͋xP��,��Mf�hMŀLl@4���Da���T�9n�[��bM������Q\23G�;!b�#+q],���N�H�ya��>{�xO�HI�k�6,��M'�	���l�ڍE��;�$��<��v�^�v!�N���ر�nFt�,%�O�����6�j/��('�J\����2!�&���wʈ��V,"R%��Zt	)�KO��e�.eC�Ҝ�!�3�M�&��j^@�7sh�m�N�W�w$IX 8�  +��h}z�0��a�8r��_8[�� c����{�	=���1@���ch��5%E����!����nZ���걗ށZ�L<�s'��s)6��b��VVf*��y�k��=�0��U�>�N�CUV~�矐��g������Z���G�0*��Ŋ�n\>����H\G��z��,�:[r��_z�'�"�0����?y�A +w��@L���3h�?���xSL��Vks�HI��F �._�1���'�i��)"!�_�q��K6����� �;~�}��-���B��J�m�Ѽo�{��nM����qD&8^ܭ���UM+m2;�So�̈h'\z[�g|ۯ�9�a%��7�����[�pTSAUe��d�=c�m�(R�@+,��␟Ƒ��v�;����e��
Vԯ�x��ґ&�v�K0�CP�UQ�)�ɕ�%��(x#8�F
�;�"wK*J��N��l�f��'�;�E�f�ԕ~A�%#Cg,�rj�pPhy����<���������c�u�th�9ǎTw]Z��)��{��f�����^�)��w+Y��H 9�;{L�6�@"����υb����k�_B���:���`��~�`@�p�&�e�;��J�b+)�_bѮx�m�|9��~�ntt��}�&G ��G��-ʟ;�f��~��Df�b�t 0��妄/ѥ�.᧝Qlˇv�(R��觐���S�:�Z"h�ԣ���~�����񉝞 �i�[(1��kF�]1̟ȫȳ#g�|��٘�U��5@��o��땓Nh���t�m�D�$��5��2���iF(�ټB�z)f��Z3����Mԋ��'#ĳ�a�8_@���#
2���P���B�0m����s�7���4�����Jm�(����M�bΙܠ�	�<�����  ͉.v`��V~��_��3t�<y##jG�[�7��x,@�tF�;Cī��!�&?nt�sZ`�+VQ3٥����Tv�Ƀ� ��`��cu�Mf��@Љi����8�/z�O�FP��j݀ه�?�NKC�7��'?�*��l�bLH��
$�:3��ʽ��!0m"�t�U7��x](�W���蛛E��뜹J��ݫJE躒�ǠO ��F��c'1���3Ӱ��ۋI�zsٔS�g+��Z��ƺ�O�����w��s
9FI6�g����t�"�ŗ_�0=`Ŋ�S~��zW����q��^�y�����yI��`N����Av$睨3��n����~�gt�����}�~irt����}Ɋ��(�tk%'4NH��N>���1��cP�W��D�hū�w`!4���+��� ��D��恶]=M�9rRDB*ɤ��ڹ[E��������0.�C@�_T�����X�KJ0�+zG���`�L5�A(�.�̒��Ťc�=a\L�^�6d �=%�T��\S�4!�u���UO�L6A^�ch����`��%/���	,�(�ђ_f�Y�>�&y�o��#�8!�VL���j�k_GL�ml[�zS��x9��FEϯ�^ԓ��{K���[�x͐�b~�Y�0T	�@Yܑ)��I�v�?n��97�+�Bö`�MZa96���H^�*�g%� �Ft;L���hi
᣷?��Ҩl@��%�����&�����4��-�k��v��w��Ǌeuc:�P�G�OL�_ZF0��bI�ߝ;��H��	��W[�VX��w�YZ��q���"g������!��$:ϘeA~O
�?ϣ��J�rvF\5�&�0#^�y�6�C��y�S�����US���{�%H�^B�d�f��y�i\�a���7��,7�R�d�D�����O�O#r�0;��!	I����z&t��VRw�����T&�&r����=��ZY��
|�I�����T)��Yj)�&/y���G��xRE��-���Ϟ�ܤ�����3V�h�Pbײ�iM�mKkTYQsrP�
��e��SU61ܬߌ�V5'�����1�=Fe)�����vy5��;n]|_AΑ{������QO��*(6YvՊ��2��(��w�fNz�f$y�����T=O�A8Nj݊F�����I/��e��V�	b��l6���`Z�F�3i1�x<~��=�ݎ�#��6�\iC8�mNn�$o)W(;�De�j�&6@��L�t>���6�s֯(�5�ANڃ-q��j�Z��o`�c�{+-�0����K��| ��gw�b�*!���`(=s ����4�Պ��� 	�j��2k��H����"P��^���� ��V��˗Ҵq��W>}P�ڥ�mm�F65qa:����#a^P��-ǻ`�N���٘1��A���ړM�?�BKd�)א�~��uކ+�%t���g��Dv�Y�Y�P�7'#�l��m��@�v�d�/r¢={��_�3���W�����[fx,>��]�f��;d�	�OGW��i�{�����;�M-J��hp��#�6
y0�o_(i�.�@x��@�)�(!���Y���a�{���DZ�|���R��3�@����g�����6�tX�{�+�(K�9��v!�r�c�L�SB�ʜP���H��G>Ϧ�׿��y��'��l���)�T�0�o�$?�C�Y�B��C"�=D���l@������g��d������|Y�g�9�<���?�$�xѷ��TTc|�'0�^mE�q�/���c(�+H�%�D��{��7Լ袅K�'=�� �J���ՈL��&Q5%:k���BP*��ꛢ�
|t�ohv�BQJ1ư�f�Z�7e���5{�D�|�J�ᢍ�v�v��	3�U�Y�%��!ޙ�/ �Z@��g����b��V��d�����a}
�:�lm���U�HY�MZ�k��>+��L���79�h�;�����/�?%���>�����	����O���S�FUv.������:=3�"U��Vl���?C��}���k%gs���h��g���ƕ�ŧz��2Yq��=�-�����Cs�._���'���� ��J���I�,D��[F�j��3�Awb�� �!����xY^�)<�����\$f����@t�R���$T�Z��~�^1CKM��v]�M�P�|
%���~QȢU��b�.H�v�j�9x�S�*=?��! D[;#"��4ƀ����x�JB:���F s���Tx�wD�l�a�2�y���J�J&����r�q���g������������u�E��Ž�4�c|���.�Ej:v[��{������^,�1|�@���]�:	V��t�#v�M���od�̔���Q�kިD�4������F/� 5a�>��Vy��K�a�~)�@
Ƀ��6�5J	����'�=R��Pl��Z�#(�^S�`�6�%$�t�{��<�6vPf~v�+/���c��r�e�KU.�M���Ww��툢|?�F��EA�#;��w	����F�iI��}[���Q8b����n�Fi�!dٛ� ��g��-�<t�́��M� ��X{��9~ E֟�݌�z�`=�R��d�8����� t1�,[�3�&{$ݗvc�!م�!���^�2�j��E����,��'8�o� ��s4!��B[�X���KL�ƥ��N�vds#6��6ԋn��ߎ.�n�/3{9��dgM�<x0�E��#,����
�,�d� ��Rܹ�g�L U�}ܮ$����W������[Pk!�#@LKޭB����B#��|B���xb����ߜG��]a�y^�"���4��"��u_Ér2�}��&�������aY�Da�tƻ�|"Kk�� ��s판u��P�7O�5��������ycϓl�	��i"Qܴ�?�ɦ_��ʔ9k�0v��Џ��'����Eخ�H��E�DF�b�Ϙ���E�V��RY'kx\�q��QӒc����F��Sl��H�΋$#���i��q򣚩�D}���j�5�A7��B�D>��W"ߟ�I��:�����c�h��p��\�y_�ݏ���D���[�����̥�i)Ooq��{�r�,ol�FH�Q5TR�g��av��+���d�Ģ~�7���oD;���U"8V������!>�Ë�E�e�D��4�f���ZK�u���I��	7��E�e�KE�����η�Q=�,l�B��G��w(�k˔ͩ�x�G!�nY����p��BK�θw�Z��2�~�4C]�x@��`�Lz'<Q��M�xF�Y���N��G#;q���,ԃ���VxE;c�c���l,�������cy�0}c�/k��NA��?�*�vv��kX:��K銘����,�^�X:f�t<FWC�bo�y�t��u���YC�۞�o�Bz`�8��k�@E�j}��9�sӑ5�O�b��M��6���!��}k���v���_
�KK�4y�6�NA������c�6�5���͡�����B+�����8<��>���~�o�X����[��o�5U����D���(Q���ʜ����z�YI�F*��H>�U��(�e�l�˧X<������+����.D<��H�|?%14��tP�N'���C����@�;1�Qw��A�LZJ
����Ƣ��E�>�cy:LO����/ʎ����O&�|#�TV�f�5)@k�GXt��X�����M����A�!���,amA��S�g�Xq��
����;m�V�mE�Z�lHmV4O�.R0��?
bu�wҝ��l
ڣ?t��2or?*�5��^��Nr��u�����
~K\^[�}��[�k�� "|��{��A�쨁�}v��-:�wM�2�/��#��ޅ��d�t@Yt��U9�+ޥW-�\m��z��~*����<?��Ӗ�E?�ĳHd��'B�,�r^��}:rǤ��M��-�sL��%=�js���bW �/�q�9^��.�N0m�zf��RdK���08,,��8S.�B\B���G"�25$�>��Zݍ��q�y�R� l{��Y�`����k��77�E�E]qSz��%��)�k�:��.L��'*,Е�"�7f�h�������~��������c.�Gf�5�.r-����=���R�XB�&/Va9�g��"��ݦn3���Ԋ�4���J�v��~�����Ғ}��%�_`N�Fo3�1x>	�s)9��Dɮ�����=d�}����r��KaZ<��sIg��?�\�5�hWXí��|Lg��,��������3e�#�L����G�K� N���v��\�^�	��8\��$�R�'��䇙�Fb�nr�pQ�[���[7/�]<�"���U������%�b���&�{�B�<������^D�2���|��%�tFcr$�Iq��;��f����v���̹�{у�/������m�X�\P[��/h�G����"r,\;��� &#�$�U�hf�!P����7y�S���za���Gm50���6�h�'��Ï���Z��tQ�c9�<�Ƙ�:�\�!�[�e�w��M⧭g�� ��n:�I�~R���VN�ٮi�D_�0�~Y6Ӗ��{[��a\/�v�A3�s�h�/��<r�Ɗ\^7 �+�_Q�Is��P��d�1xf���|Կ�Ԥ:J���d�u��3�'�����5H-�do�����Swj 0kb�LT8��>�ӿԢ9E5���3x�#t�TA�1��B<�B�{�e�ڔפ�Y�2R+��@��A����緈�|̿g���Q��{��5Be8#ur%���c!3�I��>LAO][�q�爐��*irt3����x�c�F���]�K��ZhhJ��;��A����~)��_Ð���UK?�!8�E$���1>l@g6��P���q�82B��I�8<9��MB8��f��f.~�M
��x7���4N��m��C�U]��Oڋv�W`��(cɀc,k�y������Z�_5%�j4�#�m���4��iK>y�n>�%@w�Ln��I\�wǩаL=�T���c�1�|nĵ��Z�%%�Դ�I�vI�?&��� ��Z��f���.���j)Z�7�Wd�c�nА+|�Sh�7�쩌F�v�������TV���T���|��%�]�TR��7d�W{r���xp+��e4�+��>I䛴�廖C�0OG�]�.�Qʣ�՟�u!�&���`qs�f˼u4���ȰB�U�Y,��1�@�q�?f��r�q�z�DÊ8�@��,~�cA}�mtW��ז� !�X��%��:�c���/�}��v�#�}�d?XL��tR���n�3 ۿ���Y����n�m����VeiM�a��n�ö;���8�i3��+_�pi��T
߫>ih�_�ٱ����'eU*7	�£4�r".R��~�0�Y4s�p�].Iz`�L�Р�z�A�Vp��g�a���2J�YRAs�X����{׋��Lζ��~�T����I��	@�
����'^��0.��*Y���_7"�@,�#<���K�MH=���$
񉝅YE/� ��ϩ�5��ψ�7��<�"(��.F��؞We㻝9HizO��;[��R�i���!EY�VVI�>S��O:��S�Ӷ��kq�;6��^7���٨dLK2۵���ȟ]e���o�Q8�T���IxЃ��Q�!2GY�G��L�N�9��94�#v����`�V(�JC�����u�� ����� �~�¯c�N�(3}L�����������z��\�~y��N����&X��v~c����� \���b.���(�M�o${:Q��5�����ɓ�EIt��d���3N�O�0X*�z��O��/��C�|�k�r�Y=�gZ�(Nf��%~@��������'N�g���-,Z����������L�X��*VT�¬j��}�V�K����Qp+	S�����ϋt,-
a}@�z|bꐢ`�`�B�'���{;����?��*�6��3�2��#�̧'`.w�][�X�:����oa8���3��!N+a`��s;���O�j
��:Z8����G�a��_mjz&e�i��o��c@���F�px��=��3�)t;��5��X�H��n���"P%��zJ�|�0��:8���`ze��'\��LU� ���-��;p�Q�_X��h����;�D��,�5ʅ��N�k��PЧd��Iz=K.P=��ǲE���ps��u���iH����֩�x���MQ�\±�&�	��&�G�����Q�b[m��1:gdm� �9Kв��{y��6�l�oQ�C��H�0yB��o@յ����ϝ�0�n�>UU��M�|xZ?J��|�w5���|'�_D�n��Jr �pͩ���l�2$����ǜ�E��q��e��o�F�Y|�6;��.�:�\,�v ���D�w�dy�8E���Y���cX�kҽwN�cT�tC�V�`����+Eؑ���z�U�!9�>����?X��٘��kOt\������� ��0�����r� ��`��FΧ�\c[�ޫ��a�Gk�U_A�%2ԃ�h�85g،V[A�/�c�o$Γ]���Α aT�t��6�RF%x')P�`�O�]��!Bq��ޱR!`�e���6o����wזU�����k6��
f/�B�0'�3'���%�ו	g-��+
���tl��̹�UF�[�u|��FEv������ԋ�A�F쮤��_�fJ��fG.�9���ÿ\ϟ����}����n bn�F]PE�4_��#���}�{)>c!蛎B(Mey��n�c���o��(�E?�Y-_��r��ƙo`�ޒ�����(qsI��S���8����3���Y��6��@0?���+9D� ���'�����v ۋ�5;
��Sָ�������C�0�_��!��t���ׯ̃�%��~�P�0�S�JG�m��8��)8<��Z���Ӡ�OĚ
�T�ތ�0(��2,;������ymn~b�7I�0Z3��ӂ$��%yv�-#}��n�I/�م� �	������i��mg(5�Y��xܦe��;���R�.t���V:Ne����jӉ̵#���͓&jh��([w�C���c)�;��x����b���+Ȥ�5�d!�%�[�
����1rA[��ӊя�<���1�Ń�֚��(�!�tC��7*)@�i���{N�"Z��xr���p`z�tJ�$$�z��#w�%+s+�G�#���\�T�˂Qѣ]�	w+At���y��}���S�ɋ����Tӯ؉�.��B?R��AЁ��ꑡ�b�����}��HPs-k�ɳ�\G���ѭ��m|!N-�LEj�-A���ȗF��&�y_�x/˶�K�ͩ��;.�i��13[Z�΍��"<���W��n��൛$!#���C�����2}Z�}pYf����:���ɭI҈��(�Le! �-�R���Ptґ~<}ݸ�JGXN5�2��֜l� ��G{�Lt��d�0��<c�Ɏ��SM�G���ڸZ��0?�;r5u�ԛz�FHW���bN�E��9�N��8�{���b�k�f#��O�G3���TT������ƹj���F>MF�s��L��w %���d�y�Z��^��a-Q顲�zX�
���uNTk�(ڽ�2�,�\�H���`u[(�:��6��hݥlͻJ%��4�j��aǦ�^J��灊�H����h�W31<����ο�8}�l�y�U��V����/�!���}�J��ov˹'�{,`�b|�X��i}���������WN�w˝���;���/�3]=사��J�2a�]��mtа���bZ�+�����\F��^�'�i֜t�&	�0�&���2��wpL��#!^�������1�gnL�����^�OH(�/ջ�>��-b��~�Y|��&/e�������D��kL���4N:��W�����L��� �Dti�9��~���c+G���ϰ��G��+O��@.Z}���}�'ds'��ѱZ��)]�e ���Ҵꄠp&�2�BI��/ �>s�ܬ.5�՚SR�l��ޜ�(�.���5a��c�_]�,!o��)R��r��W0mM�B�d��hCO�{G=�-#�zL�{{�:��1{4�ԩ6����,��#B�c�h�#U�6�0�YF���o[E,K���*;�P�j�H��Ȥ�V��� ���`Q^m�d2#Z+(S��;�Q��4Z��Uk����K�DY�A���)G>��"�e��O���/a��`�[nSv��&h-��$/5�`�0��8KhX�g	���S�F.����Ҝ�]���4���a�	;6\A�幏龠 ���f ���J(!��>+�{��L�1N�6l2��q��dZ��9��bU	t �a���P:7�8:�_�����}�T^�j_�P���O��1�9w�Fo��
���M�����,�}�}"����IR�f��Nr�x��'�1����o{��. ^݅����d�"UUz���H�]㙨>��A-u�2�3�f'c�qQ!��{O��ޚQ��bb����v*�C[\ڈeL	ɡ�,��]�)>$��_G�Dx�v)�V�KC���'�W�#�m+�d��)/�J���7�_�)I�F�L�)��f΅k<�|O�6��|?� Wѷn���Zo]�ï����o5}�{s�l^g$f��f����?	�;L��I�A�a�D0M�d4��(�>F7��ݩ1������3� }|��>�����x
�g�K��K	ϥ�(g(d��܎5���,4��R��O�)�oJ�:U��uqr�s���T�Z�X�l��dԚ������⍀����B������|��(���2iѶJ�>�������o4N5R��qMAV2�Ӂ[�%L���G�A_x�o,[; �n�4��ٯ_�������9�_���Ƅ��)��v���v`���ay3Y��wy�@8b)����$����3�2+'M�2�e{�F�"��ڬX.@<�a�[Ȏ��;��b��m����w�;��*��3��8A�к�z�����#�&^n�6�_���0W�x�J�}zbĕ�Q�0&^Z���&VYF����2��"E�UɪY�_*m������'N��$�Yd�|#bĲs�g<��7/���f`����ԓ�2i6Ay��uM�$�lZ��u�7�jI���cD�Wȑ>m���7z�˿�Â)�?����p���C���FqEN��b��&?t�$-��@��(��:h��F�FY�[�uYa!b�����+���V`��G
�xY��ځ�R�W��m3���E�	R�����h��>�9�<�c��N�B��s���zͦ��u�?C4�M��ۧ��2{��흂/�	|�z�=�Jx( �'/z���I~����pɵ7���(�ƻ�tS-B;4jq�>M\��V�>�3�(�;O����zVEqD�p�w����������-=qAxd}��O��z/,��vv��{�Ǘ���!ǧ6Gy�4X"Mx�|�	���E�3˥�Yp�-���U0��6ӝ��3��HU06'uSEO`���A��_f-��c�1W�����h^��
��|gq�V��.�,=X���`YDA�ʬ��3���d�&��A�\c�ʦ��^�\-��*�Ͳ�
����Pp	^S���`z�'��~k�*آD\s��d�r���� oD-�D
��� ��[:���<�t��k%���a�f��y���k�j?�X�������O�i����M� ts��Zּ��EN ��i�~�*�җ�"&_0�-xEy]gG^��Ѳ��3������$��;m��T���?��:��O������x��Gc�^{-{P}��2�2vOi�a�j���|)�A���J��ssWDZ���ݏ�i�oI�D�����@��,`~ ��[����]V}�;�A�gY�K�,��	r�E �qk���'7�7��Ͷ���LV��%���(�J����3���-�Ő��e]�hq!ocJ0�#� �τg��:t%Q��D����C��_��j�l�[�;��(Q�X��y��G鐍�b]�o{����e�����J�L.aN��w���Mh��ै_=Ց�ѿG������@��C�ٔN�6����j�D*�Ç�:��g7��RP�(���W�n�K���ƾ"��6Y�]u��S�>�+4��5�%~�ߨ�Xh5z��8Q��KQ:
�MgY!;��MH¼�N�׾���������c/�T {Uf?L�[�����A���Vg�*�w�O)����ni�
mNo�i2ut��D�M4�������1�\���Vo�ުZqia�d��N-�|�P=��0F����ĝ[s����f댝:H�A��b� ���wW�~	��ab��,�TQ��[n�$���[�J�yG��8��)C}��2 ��{㫈9+��R(���PH}jml�M������s)�L�|�O#?������0� w�B���ID���~����*����u ��;��!���ol��m���m�� Og���'+$D?|^H0��1�n�����UN�K�Sa&ZC��Y��Jx��F��;�/\`]�j�>��
%An�'hz�0��e	i���ɪ�腓[�Ϭ��W�!�`�1�����R�ďn��wyReo��>jlhAL.�V�G�C������!:�����˹�'� !]�eaT���|�,ߍo� %Iq�`SI[���R��"CoNJ��쪎q�\�Ȕ��A�a�B�f;�]�}&�-hA�*[�G���B�q��)M����ܑ�2$�/�!�<7�O���ͫ�:D�8I�2�pZ�������o�$���ns[��j= *i�|l� 2��,�s�R��,�Jo����M�qCT���A�=
��^�B�笷����3�:V��"�f0)�)W�c�W%Ҁ��T�u}��K����O���0H�������R�˔X�[�Y�t{��+;�-s���\K�_�خ* �hVwio����U z��h�� 	C6������+D"t��ҡ�
�[6����_)��[�s����(��j�}�̵�
��.z����T��ll�Z���[�k��ܱb�������n���F�_�-����ȅ���NseA�2F��}\#�<����ıU�j�_��o�jL�=g�jS���GN,�B�꿮&Xvp�