��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#���������l��U�~�׏O����j9�PY���`T���x���s����uí������P��"��b%>�1eτy�<�gܰ�N�Y�	� {��I�ɍL�ݫ�G�R�k��Q�!E	�5E��.��:�͂2��y�m�-�.E��i�����YS�
��@�H�ۼ��nD��Y�l"BU�.TԊ�=�-�����q���Ǹ��j��ԋ����tr�a�ٵ�]�b	��%�ɔe�)rYOjX5;V��R�������M\�	D��ҏ����9c=�Vͼu��Ro�P�Jf�tRvsY��c�"n�XO��	3g���Q���^�Bʹ�7gQ+Г���$�-��t�8�����A���<����l-��*�|d�ӟ�'}�.r�"��LB��d�-Sa���������|.dL�>�I���Os����{���٪W�t�9�خ��j95�e�Lt������?��%*t����ٖM¿s֧�e]Q6���U��C�@xË>�s�g��	����B���I�
�-���Y(���n�b�0���F��gW�޻/U����I��Z)C
y�(÷=�c��ru�
�{�jv�:g۞��|���;{���i��I�)^�.F{�1�����q8�Ղ��.U�����jA1��$k�y`�38A<�A�Y�V"I���N�9������$r��'`�mK������������84�1�j�}�����)���'HP� ����2d�W���һ&.�oE1��F֯�Nnw�3�^���^'&h�j��C2��gۖ�9X�PG��h^H�b�c�mwx�l.0��B�n.�rQ7�n�Vu�n�,��1v�C�f�=t{�?��A��	��8��7(��PU��-���&����`6iĻFI>6.��}l�"iѼɹ�eʱ��� �<J�9���"����@�vj.�;���|�EiR�Q�?�Kxk��I�>i���'1�+�X���7Z<�7/H�U����5�⫇�4D��D���^JU�5s�>�o���'�A�&��ߒO�u���9��� ɮ�����<��hM��c�r�JG�p4��/�y��'�e�uH��φ��^�F��+�'��������1��ۗ�L�uޟ|?+Ĕ���PԦ�-�=�����h��UЂ����͌!}�e�'Nka��L�J�Їp)���$�4�����tD��a�Ι}'��@��`�����a�����9�+��qh�}S��4��7R�F���$�PHM�XA����+0��z}EM�ƹ�";\����҇��ʀ�)ʰ5���Xl/?� |���|��ёV�˱���|u�.�kf����ޥ�:;�A�?˗N��IĐ�4RՔ~@�(�O�%�0qX��t,z������P��I���Ƈ��<W��J�UʎR�OU85+%��#Du�nw�v,_��^��Hq��I_j�~�c_��|-�Z��&@@��W����M��c���$U7%�8[?��wZ.�V\`G��H5�I�޹�����X�5���J���ݦ.��x�U4	N�+��)�*:�~�݁s	�݌�!R�ba@�`�Ȕ�ON��-\�	�����(���b�'%.C���ê=g|z�f�r{s'�"���ā�X`�Q~W�&��q.[�ŭ��6͏�b����_��'�g>�21�� ��-��i{UEb�����TN����.0�^�����Q��:��=ǈH�tRA�1��
�����&�H䊷��2;>�{W��^�7�R�O%�RKw푽�W(Su�W'�/�@��MwXU/�0�W&��'�^h���=o�Y�u�,���_�B�OQBw<�T�?í�>����P��K��!���:�������7����ua3r�6oQV�Ӭ��}SC��߻�n3�S5��K8�B���xW�ti5N)Z��h�Iɥ���]s�� N�l8P��/���y�>��D;K��������[���؅XqϞ�������b�,8W���H��#+�0-�؞�2e��a�s#��/��Fd<ã.�7,�~ ;Ŗ���}�ZC�$d�-�b��KG� 
�(�o��{Lq����b.=/�
�)��HB��abH'N�d�Z�!��Z}��ĝ[���ob2���׃$SpR���ʴ�&�v�w�)~v�(➊�Tؐ0��j��V�����C�qb��8�����"3��u��rK�Yk�v�/��9lm��#d3x��͂K�����w����[�7D#|��J���\ܺi[����*�
�u��ߋݨ�"�����3�/_��GK, �ҍ�_zT+���t��X;?v�X2YVT ��];L �d{�&�x����^C���0"ȷ�]�y��Ѭ�^�`���X�����g�@�������$@�$�AT~'�zB����&H������S��C*P��F�N� 1��c�o!kT[ŧˌU�����.� �e�nZ��;��سy���ц���<�+�f�t���w��3���MgQ�:�T��F�����U��8�} Thm.ܹ4飑^���AZ]⮦#�|�%����U�ET�6!�=�ٳS�s�W�`�:cC�����!����P�?+��Ԋ!m�1��W^�ԇ@s��)Q�Q��R7>	��q��S}����C}���=Z�ƅ����T?��0��6?�$�u����l��b
9�S�<�n�z�3}ͥ�Ԅ�Жf�?X5��l<�e��K�@��|�4����2����^�
rY2�,�ks�Unk�ر[���ڎ��t_�����5&:�6d^;оV����8@MXDl��AR[�,�4�l���C����n>qR����g��qu�9[Wˑ��闏�UkT����Ѓ^����܅��G߇�(@�`���4��(��!=��	��"n��`޻b�}��T�Y��R��V��\���
گӺ�X��_�7	�쉳��Ʉ������ʦ~ӓ,s"��ԡLM��5���1_<~�`���Zכ̩�����4f�����֧Y�~��o_�x���g&�vO��~~ ��ҭ���f8�b�R!�}��Oɮ���^�G�\����
0,�N�*_��Qh������7�<�j'�;�] �}JD��3����0��.�(G5�����_�H�c��5��Ve�i�K���
���u"|�7A�L���y�`L�b]	�Z��|`�D*VB��"T����[ny:h�d�+�\MG�} �x�Q��1:�ue-�f6��{� �eYi�>�x�YT��W\^1v���P���kM�BeN
��;���vt�E�i��I� %%L��a1n�3����` B�t2mca�2�Iw:�ra��}G`��٩ZF�����,
���"P��F��TO��\@��:���a�����P�+���\/Q��U��=V�6WP��θ���׍��MG�elǅi�����pd�fz<���a�{�c��/�G�