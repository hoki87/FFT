��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#���������l��U�~�׏O����j9�PY���`T���x���s����uí������P��"��b%>�1eτy�<�gܰ�N�Y�	� {��I�ɍL�ݫ�G�R�k��Q�!E	�5E��.��:�͂2��y�m�-�.E��i�����YS�
��@�H�ۼ��nD��Y�l"BU�.TԊ�=�-�����q���Ǹ��j��ԋ����tr�a�ٵ�]�b	��%�ɔe�)rYOjX5;V��R�������M\�	D��ҏ����9c=�Vͼu��Ro�P�Jf�tRvsY��c�"n�XO��	3g���Q���^�Bʹ�7gQ+Г���$�-��t�8�����A���<����l-��*�|dJ�M/N�[{�6+�=�e�u����l�(;���d��lE���vȼ�r�g�2�!N��"̏,��ݽ�=����(��eŦT�c�s�ƥ�����*�����/S��6|P"� �o_'^�h�l�&�4�E¢B Q,��&09 7������%�[jO:5.����%��'�(%ZG�Yf�o�;w�;R���b��}	�Uy�1Z/P:�u���ٳ�b�	`���sy4����6�OHq"����pk���1�FL*Ӽ�1#�������g'��k�0�M���9��L�dޢK {����y:2�5��mV�9َqn�G�q	p�r��PK�_�ZU�������I��$C�̩CX?"�3�䪶��q8�M����e{]3�ɕ$�d���׶�������� GA�5���%��R_�7��<�X0WZ� �ǵh�I4�	~�@�B�Q��5��Kw��;q�}R����F�K�Oz��.�dB�"���c�d2f��b�D���Y�P�a���8N��h"-p 0/��6e9i�PY��̚Cxg'X,����D����,��GL���s�GI��8�#B�����,�~
�G��(�iČ���*_�/ǒ�C�������)J����Zm�����~"�!L!���X\�`S���>�1=�H>&���,�U�����W̪�Gr��^�{�叛��~�����
��>���gK����?�x:���ݝC3�z��[�B�� 9���,y�ĩT��ۡ����a|q4D�2$�漛�b�Z]ݬ��D���C��B����:�Ci1��F�D_/ˇyy���i�k,E��ܘ���]� �c	�,j/�p<��������A1��S5ƌtl
kJ����O�Ɏ����������Ƈd���e��jD|fs�|
>��I�I54 ����;:�I%Հ����uYd���Z���A�I�t7�@s��@_�YH\m����mDY����
'
<>¸���YLe�_�oƘ��G�yn�嬨�D����v��/�#���V"��� +J�|>�9	z�w��MH/b�Ydg�5���"�ڶ�4G?y#?~���Ȁ�hn	�$��,�eރ3��)��P��8��Ot+>Cj 1�Rn
�T���u;ǹ`�88�tPҁ5{6���2�dt<x�5B2)�z��TD��@"I����>a����$2��F��	Z���[�ي�)<��3��O0w�!�Dt��X��i,�_����>�$�Em���L�*�3�r�P�l���^�8�i��e�}��䥯�������_A�VD�g?��Ά�Fr���䈧n ���9N�(��8�t������dj�ԡ�u�D���ފ��qj�r E�﹊f!q��e�Z�ݙ����ߚ���� �s������:��kx=o���xǴ&�r�%\�6�j7��������%B�k��r�+�$�AOW3�;���~�X	-�	�D�/OD|�
r�����#A��k7�+@��[m~���U�����:��@�n7��SpPh#_ Eh�9ds�'�T燏ŏ�8$ex��Y	Np�������}eKx]���l��Ką�T�H���u���QO�3ԥ90h\#��;�z���| �Gf�/J#E����:��>lA��q�bi�T�z��F�{����~�-ȹN�o��V2��2ȴ�{����I���$������w���Ynz���@��ECv��>.�#'1%��N3O�}��~�9_��5g���d�yf�8Z�W�B��lg'u�RX��J=Vޔ 03#��F5���3lcaqN�͖O3�iXç<�w���k�����c������bz7�~�(]L|M���)�����hH\-������7,��qu���!o/z��1�j�+��O}Da� ػ��'|�`�8�E6�Kk��Uiv��$��l�O</>�`��z�k*aoVa
@\��͒�$Ң�Q�=澩9��`{�:��?DU��XD͋�+�"I%+�����In˾�
,Ѓ)Ho|�G`�?C~̋nی�F���09q&�$�C�ҌN��UW|�x�$Jf7��k ǀ��Ӎ
 U?�i�g�8�������,y��1t�eV������g�[	��J����J��8���d=�����r�B��UG ���3� N�bE:�(�L��|լ"�Hˋ��������r
��g����M!��*:�t�m� o��G/}w�&c����n꼻B�:Cw�HT[i�P,�/
�Y�Ʌ?=������	"L���Le��:�R����Aɔ(���Sdh_*�H
l�dQ����
Z�+ۚ#�DB�*/' {_�@O��l|,�vm��%�E��v;�ڗ$�X?�T�Ԙ���kK�O=�&����<�yKzf���B֩m�R�������s�h� �VG��s�t��)ۥ¿{��}����A]��0Y�0)���/c�D;ز>�4�.����U�O�D�kA�S�v�%J��(1I�js!x��:�M�Kg�����]a2à��N�vB&�G�N�g�U/��� D�������
�n{�Y%���T�~VGK��%rkp�uଢ଼�\It�H5L�6��Iƾ���'���(t��G�к1�4��i���J���Dϱ; T�e]HK.	̾x���*V��{�����)�������3�ķ��������"�(��������X�b�N4�~�
@ǉvYA�aᇂ��ZO,��2N�r��p�;�G�����M��A��z�Lx�q���z���&����۲��{k�_
��T��R�P���]�Ȅ�}yBm~�է0kY��%`�=�d�%ݗF |^g��)��+*��M�CG� NS��C=���)J[
�4d��k�upq�q�D���L�+(�3e�N|���Z���4]_ s$gh�VMmX}��Vz#�bRD�̂��~.�m�j�Y�"`m�M�7�K��@�@ƫuW4����X��T���A|��*��$J2X��\��K�p)O��*���}�ErWu��!]�Gn(���q��3 ��H��F�(=�/�wUM���)C�d�{�u�/��l����d'�EΎg�����/ؐ�|N!�U�LU�|C˾ �{�i޾ctiA1Xx��,�'P <3XQ�<�z	�$Y�(��h�C=�����ykx�<A1�����$b:�g�8��?϶�85��oޖ�5�|�y9��
����-�
\��t�,���p���!N�׼��/�"cT���E���p <��pL�|PE�1O�$3�*Xa}��	���=S��k�d�4�a�Ĳ#��3*]���7T3�ՠ��:�4�9�����y�77.�V��S4��ŋ	�-[.�B�͋nU�oVr<7�`9��C@��5[�=eL0eb���;Ql�[�)�})����U�i�������c�[ [E�W-�f2oj���� 	��&�O\Nx���>?@��:Z~B`�:Y�XS��dn�����nlH(N�8�YZ<�Ϯ�T��~!j�YR��S��?x½�'�n�Z��l�;�~�C��@��,��9hA���W���%6�����N4��~�˱hU��SخA!7&KsűgW�~u�]<ƽ���#@q;�}���HBֲ��m��^����[>��}��b�~�:C��z�+B�|6�㽛��n���k�5қB;�����ʨ�^(~��)NRC�`<�/����$Z�D��F����HE�%������c�����>��>Y���KI�@u�vU`���{$GQ��g��� ��nƙ�R��$�Ǉ��#�p�.���))�t�-�ɯF:G�OA�u�皜�U}��9���z5����T���m�g�jE_�uW�9q��
������O�ȲXԩ��g��.WR�&�}���7�7-0����R���I��\��C����K;ӗh��_�&��O�4Ij�wu_����z۫C���!yC�E�R�< ��X�Q���ʇ�gү?��<�ʟ�-��ݶ�\��xR50����鰺-�>���{jb<K�n�Mrʫ�-�Ga�� e�D���ڮ�Xv��A��c�V�+�H����[m�4�č��V3ʇ;v�Cj�Xv�,���5�+���ɒ;ut�I�xΕ���m���b��P�!�\
�/a�r��p��3���9OT�\�+^��+�w�|��Cli_�RM �/{�g���e�}�k�-�0����5M�}y�`���+OC#�ؔ��!#YJB�W��`{O�@yF����`"�0�����=8���a�c��f�o��bѻ�%��h?�D5;]���N��E1V��O���5�:o������EC�y�;F�q��r�]���+#%i&Rv�,AX��=n��$K�?P�qѼ��D���{i��Y�U�)���& �в���1�|�k>���ȎM��O��W��k��x}�x��ɽ�3~��@�2[�i`�0M:�����ϗtV�۱���V!���Bۂ�BA�X02��:�B����݉^�#�k��܋�k�L�ǀ��2P�m�ҕ�o�vA ���N� #XӁC���m嬤b�G8[֔ c c|_��$�m�;�=o<'S̕XYQ;�]�{<�ˋ�qv��d�-�����?5G��lᱱ
#Gsd�$2}IGcG2Q�:,ac�uҖWH+��� ���8��(<i�����v�s-���h��>�#��e��(�k�~f�2*Vw���3X��:���Q��K7�eG����p�E9ɉ�yһ����!�ї���#�U�9#��_Ы��0.p|��T�)�	=h��;l �@4�������,rqSD��Qk:���:����!�-"�c&^�q,��NC�o��	�x�W��߸|�=lc�D.U1zSBy
q@�ھ�{� 	�%�f�"}=��$��lS�Y.�[>�)�����E>�]/�2c4 ��y/�����*p��)��Y�z� �'�" d�8����,����5��i����kB�o��7*��H��t�l�w2��8���8�� ��%&I�(2Te7�C�j]Z�()߷p��@�9��J�(xu�c�������ݰu�y�˵�t5��gf��R���?!�44�ޱQG\�j�P��q]����<�&���_�Q#Ͱ6����FP�D������:�6}�q���l)�4l�+��Ή��ݭ��E��1u���K�V�1/DlT��~��wÈ���4I���������q�m|��
m��I��n���'G�J�� ��u� �Gx���x��V�23��AyH�DP��y�24 ����"�A���Op��Xx�)
B�.SuX�<}B7�ho�>�/� E &nH2 �����_���JO'�i��Z"d�W�#�� ڔ���G"�0����dK��B���qcS?�~��qz�>~ 9&�|X�6i�C������.
���J#��g��jK�yV��o g'ǲ�aO�1}s�l1&�	"���>Ƚ��Cߟ�a�?/��k|⛡�V��**C�+�OJ
r��L錒^dE��e~�	@�#��v�n�n3�8c��G���3Z��LB��jX'�t^�&�9@�p]*fM�H�c�=�g����FX.�̀�(�%���$�h��$�=.�r^�u��~�����F��*SY���^�t��>8��5
���ihѩ�2��-�3�\!&YW n�>*��K�n���J�ΉFb���5���uY&����l"o��	褸��R�zc9p����?���s���S������c�_#���[.9F?ĉ�+�zݳ�_��5h[�Gi{8�.�Ɓ��킾�G&��*2.^m��&� �[�KS�xy�)�����4�(j�95Z�W�\n��
M�tn^i6N�FO�=l�-5`XQ�|����S�Uю���{o��W#�zO\q����D�rs��d������+�%�3�=��ӏj����-�d������)fPj۰6�4��gÄO4ƆO�ilS�&8��$��rs=P��t�qꔼ���>;[��	��9���4ls4\��~���/�N�0U�*��}5>!������S��� ���c^��聿:��m>}�i�V��%�ĝ�?df�:���s���w��qB4K���l!Q-��M݀�7�d�*�"��u櫎2� =�fd�&�-�?X��(��hE%��0
F|�%88��P�5{݈���E�$�����^�㖫��8��A��Y�pJ/9 p܇�P�N���t�"6���j�^)��#�i쇜�3�w��Dvm��=ϖ�'}�n���D�Sꧺ�:�S����P�݀��A��N����մ�~�����j�dh���3�o��lA/q���鳜�S�~}���Of�M��pu��|�[�،{���^V��I�-'~3��DR��h�֛�R��{{zH�W�\����f�_s�������#���hݜ�ّ�1��g�y���:;��߇����,��#�{.)������a��Cy{h�������uwv~��->���S �Ҕ�]��,�y�W�����I�.9^�"�uǄ���F�����iS�rS!w�Ė%�H���>uKB_*s�Z.k#}�o���@d���U��<ޓ�d��+�(J`幠Ń��mR��-���"�ǭp��+>��K3����[��Q�NW�VH����8�P��-#ߐ#$l�E+6`�9���/, �h��4�Y $l�&��ȡ�u�md��A����!����H��<���{��T:LM᥏�ɕ�l��d��Eb԰��<q۪�����rA�.�2x7A,&1�!�Z���֠3+d��5�7.�FM�C���^�a�%x�p�;��,�O�<	c��D
`ԭ,a�)�6U���k�x�"���uYU*a߻.RY/��4~��X,B�#��JK����A�HL���^�:׀hu�Oݪ��IzB	�/���PH�����ؠWW2v��ML�1�	G���$Z���2V�n���r�d��L.������(��"ܷ_Y�n��@�����M6s�M��-���*�%D����t�f)�/�\�@3OQ_.]|��!�p��|mjٻ����Қ�&�B0M�6<���.!�����3��|+t��@v��Q��&\���prň��T���
��MZ&�z�.Kf��.SҿM�[.m3�+�s�x���H�;1��ħ�wBXd$R�5;N'�'��k^���+J$����j3���`i�R¥��-:9)�����owq�?^¶��%�/�z�$�$y��������'$�t��g
7$�-"�Mr��+��Kl$��V��`@Az�NU�Y	�,�{E��NXE�M�~�����E�H�c$Rtѩ.��dU��k�?_5%�+S1�����Ҍ�ֿ�l�%oY6ezO��3����7��cZ�/�j��3���f��^���a؅ *4���){� *#�<�aAo(���2~q����7n��1(�0�=$��@A:��-�C�g�s�Ca�t6��ӎ�j��W8wk~�YQUi%��߉2g΃fr�qP��`w{��h������:���i�Wn��7>�+��~�]�
��|��mBv`�t�/{�6�$;ҌM��&�5�Ѩ��N�w(��La���񳹳%��"F B�;��-�6��l�Uo����kyv�h�o�G�:�B��� ���H��9�����Ƶ���~�<������l�\��DUC�m�L$�s}'�c�["4Y4۾���I���$��i���2�¨Z��
��uT�Tcj5l9M�%7ц�\�V��|:Y�mg�{���9�j�aoHU}V�K��m��1l��.�<q�Э�W��i�
U>q7wU��I hPhV��_�[>#�9<��)��`�KS-g<����S��p��2�[��S9̇�!>��:�P&���2V�uт������DPy^~�v
�~3����Z
��ZE��	���o&!x��E8�}C�j=�ب��;JXh��II�;=P��fsӅ淆>�3) i?�x�i����	� ��lV���o}t|�T�#���ȇ[,��c�_����..�j�<�NL��z�r���V���p�8���fu���z{�[B��bC.�E� �(���W��ok9_�;����וs��İXǷ���j�O*���]t"��[�9�l�'��~�H�g�V����4�E*�l'K�(�ƅ�����CI���vV
�m}q�����/i�R���ڥ��<����_E_ �I��K����7c	�F�ݧW�Vˮ{NZ��-�x��nZ�?b͢���r�6l�8O}����������:�ݓ������W�>��Q�.��q���7%���6 <�w��~�o��6w�

ktc�����	�O��}�����WU�Ӽ��'v������S�D�ac���4��8H�ߌ��<���zc*��iQ��؏���٫��z.��h�x��W}:h�%/�E�ʹ�f�+��@eƶ ��n�����S<b%��C�=0���2ե�{�����5c��sFf͑ =IJ f�"K���T�F���c���L�,Cu��D��T�K�?�~�5�
&L�<:�0���T-[�J�\��eMW�H�U+��(ޜ���t�6�o�kpu��`�4�9G�o}��{���]�F0mf�s/�v̭��@�"8�����͜�죐�Zˉ����'4�ٮ&�#1�.��q�0�H
�`�rs�ݟB�ݰ�Ҿo[#��^���H��L�F���4�P^Y�=s��Bs�p)�0����T���JL��ޛ���bI�@�6�T�_%\�C^m ��\`�3�'� �t���md@�5���;�W��WhaDt�,�Jʷ�-���P��0 ���"�GH�9�q���F�c�a�.�TF`+R18(]�*�E��ى�a:;�ހ��4���BG��q��PG�+rG��L�n�¿�1����VȫM��N�J�3��F$U���M�H�up=�:?�]�5x���.ok�K��f\���㿤\�s����˥&F+.Q�X$~���X``}^AKb�g"��.>U{yz"fg����4=���@� q�G3$M�>�u�c.��S?��C8�	^�6O��>� �[�%��D5�ui�4&�h�m劖Z��T�͖C#o�E[w���f�x����CIx M3w`�m�E.� \�v�5����B�!�c�M���#1i9�s����a��+"6#M8qm�8c���t4�%���)�8v 鏴b��]QYa�H/7�WW���j8�`�����t�U�@U������>��n]�{WQ�@�/��C���'� �Ig�h�V���ڼZ�?��7T#���E���p�� �L]-��^i�	��K�	s�����>)�s~H�Y�����0�E�;gN{�N&h�1�I��<�&,0�����@<�r���Y�_�IJǼ�	j��P�P:�Y����G���A`��?;XH$��(��C�b0K��(O�"4Y,U,���� �1p�1����j;�lՓ#��i4x�s2?D��������Ә&Q(̾�7�ڽ@�����LR=� �f#�G������`](�^ZP�4Ԇ���������?�5Ȼ�V6 �JL%>�팄�ei|�d��ʍĪW�-zo����b��̢̥[]��
�D��
�`�3ĝg�b�&rS�v_a2���	Z�"��;�i\���S��@4`H�K|�D�,Y��5ފ���{kl@S���i&��'��	��f�P���N1����ޒ?��s�t	�Ns���g�KJx����Y�-%����|v�`������S��y��7d�ϔa^���5^%p������JP��jLnVк��4��1{��+Ժ�"�}#��<�e�ᯀ
�3$���v�s7Ka9Tq��w��ޣ�g]���"ͱ��ЗG��_��20�];2��5 �r����t�t������#���5v�}�`�uq'�Ӄs��~q�~[C�Ⱦ*��<�x=.R7�|s�_�/fb�����D�����.��,R̰�S�fDQ���!uǖ��Ӆ����su�e����°�o8�1&����u��kZi
[J�u�g�N���
����`7o��;])���~�E���uO9<z+[��1�?���>���r��/���	$�c]/Pl͢��.����7�ȩf���I\61ԑR-���N�������m�D�*�K�0m��-��f�N��̵]Ñ�m�����I�^�=pe��_9�����Ơ{��#ԉ`��ᵘ
�N6�Lz�|W���j��R:�9�[#�D��ͱ\A��t��	��0��G<U\�f0�X�z��s��4��XF�{���F��elh���zj2M�xayӊ�8�`)��ϩVs@��N0�߿����?�E����u�qD�~@){�wk�j��͚�L�޺B�0|eoN��c���F���e�d��Y���᪫s�+�+��=ɔ����8k���I�CQfE1�:o�M>e\r�G��G���O^��hJ��XO��~n��=�)y<ߐlZ�{��x���82&� ��d����+)�|����fDD	G��%k��u������ۗ�vo��׽&�5[<Knp:�+ŵ�p����.�c=��W?�v҉ƚ.�w�1�3�n��vv�F�鏔���4������V�<q�W˫�����U�үU���{ɽ�����涥�	/�����!��T�;����~��v`-�O��u7ؕ0�Z������~'Z��;<ZRDT��ydz�.��r34�ז�u(�u"�0�o��@��<>��7�z _C�&&�Q|'H5u)��I���aN.��I���ط�iZ3�0�wb��x�E�~��"p���ɪ�ژŢ���9�؞k�z�3>�l��1��ϙ� P�@�Q��  ��Ub��Cb�z���1��>�_�/a��YqA��b��S�xJ�cE�b4P)�РLd)�~l����X� =~�@���Ʌq(�"Z�8���>�� ���o����bƆ��_pÊ��r�Y�Xӽ�8�Osv�7�<�B*D$�݂��.��ј�1Ƴ��3�xg}����̴�J���&U���&�hޞ�̴��0hk9���^�լ[s|>�0�W���[��!�������pF6�Y^	]P�'#gK���'�s����Z�X�X/7�V9X� ,�yy;A�V�Z<-X���*1�zh��X��!d �k�*[�,��Ԃ>�h-��o��m�P��K�{:�Y�w��B Nc��osK:��,���6�9�{'P�
+FH�<'�tf�(��m#J�	�A���P�q��q����v��?0�ս�1^�D>��}�Rf�@EX�RC����1�mDݷG�C򾈠��R����� 
�-(���ů4��z2`�7r8���Q;�v�^��F,�F��M'�/#׬���p'�I8KM6��L
H����V;R�ϣ�$�D/?�M�̳�s�Gl^�и:��%4��J����FɿsȄ̘ ��1�����wK��'�(�COA
��
Ŏ���0��?�<���qf���?r�c�\�ǚ�������w����v�Dsێ��d�{��+(��/���M��{�gfe�#зC͈�_�G�f=I0��"*�t�]��*ڌ��e�E���Z�%M+��r  �̀N��E�������~�6�j�.&fx��m8�P��fp���/旾�j�ڪ;J,��yz���H�
�ʮ�|�p[�'.b�ț�֑���͸BQʣ�Ufk�����K�P�B�,�jܑ�jч���'FpR;��-����;RT�[x�\�X_�E��)?hW�┼�����n���`��k��}� Gzɝ�w�9tj�0G=�.��-��Ҧx=�qi��EM�6ݿ���0��Y7v�OX�/`�.�"�#��"]��d����a�z�!�c�r�Cd}�/n)�=6��ʢ�F�N��ο4,h�e�/X`�]��m*M)�ۈ9Y}o�3�bj�TlW���&����<ǚ0�v4�Ǝ��ă4���	{�bH,��PQ�O��y���6�Ũ� ����?�����3�cd�}R���z�u���+�������՟!S2'd��M~�.�qWk��[8��nP��O:�}���F�76��\;��gl��)"�4[;nZ�OF�[�d ���)�E8�[=m�	O��p���7Y�Ƞ�~ZD�)��	��^Ϛ��W-��`���O�쳈��W8�8bG�5��@�RI_@���Ę�Өi�ר�Q������ˌ�=6iY!�vN�8�T&PD�G�!&��|�rɅ����k�!��y�4�%�孔?�7[
�G�:F
G�<�cc���9���]d�M$
���d5���A`n�,0?�B^��+>E��y��q��p���çhST��	.�Y�gV>f`҉�B�*���s��pb�+@+nN-ᵑ� ��d���ZQ�_���B۴�Qn�&.��1��!Pq]��
��jBک<�xO,�n�}
�����<�~�֋��L�Q�+��xp�~��<0Ys�����G�hSq�$�HF��Δ�e���s�U�K�Uu��U�W�7�2�'���4���J���U���r���6��:=�h$m|���~���dY���:�� =��l�	N��B��2�НBً�)��h_�����V>�;T����4b�Tٳ/ݷL��%�Qs��i��J[�y�z�3Ҷ��{�ӷ�4~	��L�+�T�0�+��Ʃ�}�Sh�nIh���pX���?:���̍2�B�l���a.{a�|>wan �Mkx
ng�����иިA�
#���K�6�鯊��lgv��"�)�q��&��_�,�%�IU�G�h\�n��]����ŭ���C;Iů�X���[@US�9���C���Aդ��,l.��c�St4�o gH���i���?��b�d�3W(!�'�v<�&"��)`�Q�5;�d�H�����Ym��('͡� s⮶��d��E:rZ_���vA�)�&U3dʵ� �8��m+�Զ~B� C�SJ����5s�oT�#J��hX����0:\5�N�{t��Q[�b�⧼�@�U����.ִ��Q8���dO�����w���@�o�5�d��.�<&�֪��%bŮ��K�t�5�6��Dq��n|� �Qt�TI�=�6s$�.@��i<�a����?DN�Bl���#�R����^
=8E� ����3��Di�h��hY�
`��A�
f�vQqiϋ��G��Ỷas�F�&%e��TI��E�Gs���=��4�j�}�ʮ= �^���3�4�&m,� ��?�A��B��9Kh^�l�6��?@}��ˠ ;u��Wr��>��t�ו<����A�%�؛�;S]0#Q�$����)�}�j���?( ���?���w��X�_���
~�S*ٛ��B���v�W������G ��E@,b[Y���})/��r��qj�rV:"�bSd*l0���w,ae"�Fz��d��ԏ�-��s�!����[��7��`�M�6i^'�c�q�-Kz)<[ƺ̷�xӶC'��,xآ�o��=������if#,�i��5���f��v#9�#'�e[�o��U�B��a���>�d���ǒ^��{�x�㌹��p ̲[o�����߻--�S��u䃐�	��b���E9�9E�k����t`��s� ���9.�Qf���I��} ��G�m�-=�8
|!.�����}��@�)�.�逅J����"� �܈7%6���6IVU������O@�&>C�A��ui`��r_�v���kk���A$�09hk�2b����©>_Y�f5+�)C,1܎$o�*j�2&E..'"�;���]EA6����͎�(J�� ŏ؏�
���&��ӎ]^�C_�gfO�Z��(e]��mn{o��V-y���+?S�[ɀ�u�V��{.O�	&�b�d��b�����E7c+��7��M��D` Čb�װ-�S�j���J�&{G8BE�z$��!�3K�����E�<:�PBe� p����c=K뤸����-���<��f��O���G�="��$���lx��b�K��MZ`Y��e��\��h��g+�|��EhP{��	���TUb�8a+[W��	�9�B��T�N �3�S��#Z����E�,�lջt��2�0J2��[���w��{�'�e�U�l���^ֵ����<�,��'����h?�<v��Pݮ"�a����
��e��¤��Ni������-��E��%u��z.v�6
f��cm�{CG�q@Ŝ)ק��-EXq ��0�b�?tZD�����"=5+�������`�*��Vp��G�)FQƀn)l�{�w����O�8	����Y�UgE�T9M�c�S~����Z�XQ����Q�2$-���6<�ۼ�p�e+�9��� �y�������x��B�ܬl���
�bʜ�c�e�,V�j���&{�����>3a?@S4D�\�(頰(
�,h�G/�4-rʂDO�?��]p�ˤ��FR��W��g��{��V⪠XFwV�=z��G�`i�\]�S��ea��%K��R��|�-���+����xv-�x���M�V!�wu�%��6 �!� �o��g��C��� (�O�\&>�j�9p���7=��:�zyJq�L������ݝ�q%�dš�I��I��w1-vTɩ�k�(��MފT�r���X8է�1�\v�ܦ*�Σ`��*��O�\JUwc���{�-.X�Z/�C�[R�S�ߧ{�?x����1��'�`l����옉��-�E,���-4bO*.��h��B(mT��k���A�t�7�C�B���j&m�u��]R��`/���)=d�s�*���#K5��u���4�x�}2��[�nD��F��$�%�y�}��J���H�(q}��Ev/�-���ZDsG�����
���X��:ڔ��N�	r�]5�Z����p�):�,c��Y_4��M�w�����/y���1�um�6�e���;��JM�R݊�EG����������}-r�
��bH��n��9�����u�ч	�uZ@+nuZ.��gI�q'��8ng��ʘ�Y����uX�}��)�γp%!4��\]��Ť�]�2�z�IfntQY�e֑���&�ߝT�=��8�ᇰUfDg�1��t�
t���b%�f1S�-���m��G;fZ��<[��\��_��Z�t�r�:��S����l�׭�*���q{���c3
����׹�X�!.t`}�˧o7��ۮ_[���_��5S�3�iO��S�׽�q-�(���on�����py��zDy��6�9f���B�VT�D2�o����S��P�_�6�2ʖ,��N
����[�օ�Q����@Ţ�T�s�h~|���f[7�:ye��m9y��;?9���c�s�wX��Bl���H��k;�a�%L�D�`�m��F[�E���<��IH��Df�e�~�����%o#��C^���2�����F�a��8�c�m锵��X�pXP`��:8�}�Uv"s�pAM���
~H�t-�z���A�7��E��v��N�t��Be�_J���šY����������s�4�*�/W5(��=b�;/���6nOaV^GM�Ԅ�-��w� ��2��2^V1�ώ���tN�",�&�w'}���,o�OK��"z��������=	��j��iUDK/j_�/w�~�G]s���HJU�ؐ����Q�*�3��>�4\�y�3%�k�!�	_���y�$y�v��O��3�z�+�D��k�I���[(����K��ƕAk ����A�k��������S$8h�F����K����c{�FJvag��¢ս���6��E�D&Y*=Ϊ�C#��s�r���1�{�zŔ{y���*SѓC:�}JL�Vf�ٍ���T�uq��-CXۛH�h!@U.�#�D�e�0A�0�C"�Z�p�q]�ay�e}���$���z�Q����xRt�bK�u�ޭ��l��{xz����re��v8DR|`��^����ݐ����G�Nƫ��5t+f����&hӷ��+��H�.�Z��̡F�n
�?wG��l2.�j!w�9�k� s��놺q�)m��h��^`t����vDiײD2�1���$F��<+1'�i|6��bf<�O��0^g^�܀_���h/aE#�I�~,�S�?�7�HfX��]R����¥Λ�%
���F(��6�����<J:�ƉP矵� �g��]�ǦO��C�w3�I	/��4��_�4��	�!��:�XKG�.�KrCXj,G���ظ�!\*�Q�'��u�1��
�G�
�3�P�[A�����]�Q�`X�\��4sV�#S&�JJ�ަ��^q9�0sw���H� C�)�%E�(vD��7׭�c�}����Rb�oYn��&8dESu�_f��@�vF8�]�!"'�uk�M�ہc_�Y���޾��Կ��+���DЭQ����i|�_����7Z�f�#4�����Unlɿ��r�'���<j�n��<j/-�羗Na�����85O9��(�V?����=�DKK��#),�f��Z��{��E�s%�P��
~�`��Vh+ՉӏϚ2��ꐑ�x��Sp����S?6�Vs/�I���$j�;�o�I���|��Tc0��"R]��\��r��$��odi�f��W���Q�Z���ˇ����ݙ��5�m�U��sJ��M��g�d�?���S��)�J_���6��^���v]W�8+�ѭ,2�I�|
6���ˉ
�].��M��	[ �E��k��,���~�Z�6�P��Tt׎�o��"y���Z0>��9�Ȉ���,����S�?��<]_�yȲ�L�Sު�����G+�$��vL��_�,����W-�t)X��;4.DmP=|σN(N^;��P	DJ��aJ�4]cX"�
!Q���ʾ-�Ot�>��,i�S��ǢO� jS�+T
��X��}�G�P)�w&cj�*�{׾�MC�H��a���fO�n�J�v,>��D����S[� ��DI�8W�0��<����F$�x+7�A�3o��d+��G(���S�P�D�ݑC�� P ����|I�ˏ�,���p����:��ʏ�@� �y�0��.<��#_��p	�v~�[=�i�q�ݳ������~�>csul�;��$�o"7(n�(��HX�2R��D� G`J@[$U�U�+�4Q�$a�3g����^)�NW����~%�����"�����H0�{5W������׭��"k�Ǿh���9[`@ʒ��vT���6��a�IpS}r_0`���>�C��Ȱ���q($��&2��A]��^����c\�@��2Fq�nA48����<�C�E�m *U�tvyX� Lx$E<�?���q�r�إ��z�F�������$�YH焕��9�l��Ҵ�&��Ҽy���s��*[X\�Cļ-Ћ6�;��7�:���+�����j�'�Zc��M:�\^n[w�N	4��7���3�@����ۧ?1�a��A�Y�X���s$�������"G�#6�/�8���o�o�p��]'����'�rw����%Ep����w�H@b�"#U�b
2riD����5����x�,8
�k�rt���s�T����+N��2���2 )�����"�]q�O-�C�42�?l)vr���dm�6b5?�&�V�C����W9�T��my��w6}G\�T���-�;ƉU���-g#�8� �G���r��4V��Fo���r5/�v�{����j']9�-���K����4؉�����դm�� y?���j��c�k#p��MK��=./�Y���{7x�樝��!�@�	����)���#^%���^�I}0J��n�bJ+�h��f�8��,2&��ƀ5	�t�jpF�t���K�ן��΅���8�@S�:�m�D.T�˕YEM������n�KT-��qc�F��b˞�T��&�b�a�4��{f�(�U��Iy&�~�"��H��=���}�#g	<Z�e~6F�_A!<�3X2T�!ņJ�6�����Q���8�J�7"3�!P�U~9�/B|Sns��	�o����]@���A�ٜ�d��?��}�]���J\��9Z��tͶʔg!Ġ[߃���l��\�=��܌R�2�2\[@�ꨫ&@���kM��y��D8�x_��C��4�?�Y3{2�3D#s�����Ͻ����s�a��q����^;�$���z�k=W���x�#$/2Up�K.�Ht>1rw-a���!�ae�9��_���M�����n>Gx��:juv�s�-v����ǈ�T���Nf�M{h1>���39k!�W�4�tƜ���8VGѺ.�f���;�\qb��!Y_�Wݧ�/&$S�g�9����6"к�>� �!k
52\�ݸӇ:��l[��怢�B��j�;!q�q��&�9V�� ˆGl�z@Y��KHB�hQBE�� �G�Q�\�	�D�.��v��a����~����fp�S-SO�c7Y��ߟG����Qܣ�8=�R�ɴ�UC�e[��2o��2_�!��jS^������o�0��X\����,m��j:�������#�}eP���
��Qs��?e�o����Z��O�~<����#U���_^na/5V����g�1VA���������y=Ĳ���G���æ���_tX�)��	2��"Y��������
(��7����1^#2x�����.HF���<���u���n��&���C	�vsf]�¸xf^��EH*�9�L�t�͸�qӴd��>�%t�)e����=�����R��Q|uYG��]̍�h����f->�v��U���\��#~����C݋5�Ă���e)�>�0
�r��9l�\sF�h��#/�"P��)Y����M_h"Y�W�dG;o��Z�6;�+�8�%�v��<ћ��{�i,�|䙇��}�Z�] J1~��3@�Z�qL��z`3`ʎ��ς2Ś"��lCV����(4ᰠ" 4���4�-;f�d���\�+W����b��q�^��%&���x�oe��?,c��7���r:R�n��\��������Y���E��B�h�j�yr�X3�����a��fӶ����3l�Wc!$?N\$��
�M?2�RA�Y�n�[c!h�TrO�-!I�>�p��0����޵����P��(\iK��׃�v {�,Ջ�+k�{'�+�Îb=~y�m�ʉI�XG�L� �B�t-�P�NXUM��f�L1ί���Q	��;���2��J���{�S��گ��׾��kP�{��m�u� �&�t`M���0��o<���l���K�����2�y��1+U{�y��Wi � �/��l&�>�_\Y.x�Zߙ����{4��:���d+ �mϴ %���GH>�v@�Ӷ˕�X3�oJ^��C��z��Ȝ�?i�|>��M#��-�	W���R��H07��P{2����aYm�h���DA����کQ�VdAn:����y}��
)J�DU-B�zlL�`�r��ט)���c��Z9¿�s����xJ�_�R�*��f�~{��~��׈�9L��� g�[�ͣ���u*f]$�=�8����6��I�9��X�0�Z���\t6b��`�4��`��as��@������΀vfy%���_��i��>���"q�r�2C|�V�٘��kl��cpd���i�e�=!����Vy
��p5~�Tn�V+�z@?/K"����ϔ�b�wL�!�ml��#H���C�>�'�{*|x68��t�����l��)) `�/�t� ��9`�#�#\����y��2��jW��IK5N?T��>�t��8�	
g��8}���\{P�^.�v�a�����xO:��	��l��L��2mq��R/q�+:@��y��Q�r{s�]��p;0V���bYI��6�z��h��!JJT�-2�S�H��h�1O�x�36F��_1&����E7���v���ǔ��)�Qk=��^ہ����f>�M�R[��;g�X-�J�$�(6r_�9:+[��*�JA �ޮ?#�3��
��~���.<�6�H���#��%�x}}2U~w�"!�#�@!VI��$�W.�W>ϓ����Kk>��.J����� ���6��P>���9c��!�2%!L�E~;�����dƄQp��9'��g5��{�l�.2 yl�:�5��n֫,RÁ�{��s�?qV�S�vd�T��o�?��\����5��ހ*�똘��������r��^<��ǀ6I�I$lG�w\�	<g�5���[[�n-��H�* �.����#L�؀T`ü�-��hb���'J0-��[�t�r���;�'{��|�͵Mzw��N�A�(��$��]��z)����e�ִ�p
��cM1 �~��Nf��D�˙���q�+y�M��L��=���_u�$��J�s�Ť�p�X�vv�l�ø�g<'�~��&�KO;���i.i�G��5�P�`B�)}��I'�l�=��&(S�tE�7�n�%�s��WA�.�d?]��ز�}*�Lh�
��t!F.�l�#G}��P�q���U�����/b��6�h�ZC�N;{���~���&�1�ٖe��"�`�,�|]��m�lg��+����i�v=���P$A,DkXAL̲�c�f;�34�z'E�Ѩ ��@s��*Z��@��i���g;h.�>�����'����B��n` ����=��*���Å��9I+���~�ʊW�C!�=���|���i���/+��鹼�i:L.b��k���lH�|����#%Cͧ�"��u���� �[3�^X��w�/l�5�=@?ӥ�x��ڵ�I�i�"N�nj
��ƀ(�'�9�ߦ\^�@�L��8�]}����1C�����B�U?�Հ�+�&�>P��h�+���_�uAF������Y'1�0�pl6����?A��B?�&���痺�_Y��a�x�iNƳ���Qʗx��(�U��9}�^�t�y/���=��ජ������/$1��c�H}�B]�, o��J� ��I��o��ނ=_�{1�%ߚ���Ro�JF��CX��^ ]}II������*���@���N���W�I��>V��Dt�o��f�4l�J(��Ю7B'e�.dq����Zm��k{0�Й&!'��Ti=;p��Ѝ5�Όb���쉝�y�y�(��|��p�\�o�Rxl�Ir�@65�e���{?>P���2�.��7,A���B�"��+����W�@�L.0q�Lk�����o���/E��Ŏ�d��E����iyM�M|`�g�-�;�L!���P���פCB�hj=Ly\�B�gRT� ��(R"n�u�F�i�L{�^�Ͼ�r���eB��T<�g��ﵳF6��k�,߃ɘ9��u�����ƽ:7�x�M��.3w(ΥCVy���@��Iw%pU0 ��5-&�m*�vS����:L��X'�͙�**ZBA.@���$8���R�| ���2�q8��ӻ�/ 7�Yj��pӀ@���|�E��#�D�� �' r�����-ĥ����W���&z�i:3��E�$C�Z9�����Aܪ��8^�Ȋ���<s�2{�.�JH�y���"�H�Sŭqוs�%tۉ�yB/���n*��I8́q=�ȉ�D�ƻ,V�g.��I�����I�?X�E|����)Y�xE9�տ��$JDi�'A��x���]�[[OVvD����MTW��g�\L�hFO:H�V�wӃ��W:�$'p���9��R���<h������Ϡ'��M'��n2/]3�7���^>�׊��K/e4A�����38Rr�T<N@��|S�XY��!Cu L��H���F^���m ��SĽֵ�*æ��-�	��ak�����	]:\�a��rS��J""�������4����#�3J�"@�v\�}J|c��*	��vvg�/�h#���ѧې)7!o�S���۟�-�(4mp�N[i���	d���
C(�c��ZJl}ԋ-�H "$w�;�6*�6�� �e3��}J[Y6��$`BɒZ_u�ID����׻�[�pҫ����[k�h0��0����2���J�-��ڱ�K��d٢Y���Cc�*���39��>礆C�M�.��i>�M¿-p�ΰ��l�#nLy�p�g��B���`����¡������Hل��-�>b�j,�Cɂ:��X�\�Ƶ�A�ot��r�ӏ!?�P��౧��ͼg����N��^���^RK¿%�E�R�&�#�1�0fM�XE`�+\Uە��@��+�ĖR�4��}q���,�c8`_}���;�dX�;�QҤ�a�R��w�t��[�6m�PQ+�8r���jM��-�.n7� }�}�"}8����z0������,*sr{Jx�+`����u�Y$c��m9�r��к�y�N����a���s�?�%fFm]�%��s�1���`�M���w��	) ��(I� cv�Vo\ƍ�LU*���{π�#nԈ����C&�!k��l���3�-���QP�����d�դ�H�9�q��^�H�{X��o7>3��1R�s�J���R���J���傔:J��iM�ld��<�PX�s��mfnb�i�,Δ�6ی"��#���Di��܏�&����#�,�㪲��Q'�˵c���iz,gW�+k�f�'�>F��*�QG�9��x���,��ɚ2�	�+Hӆ����k�hc�yY,��vȻ������b	�[�@r�g �H8��$�}����7�?���w�m�Q�!@���rxm�ER?�Bf6~%$���҆��*ū���ك��.f{�����D���7�܌_G���$���h�:tHX�<x��.$�.�@0\�=� (Lc�������X�Ɋ�TL����X"�*��L�Ƙ�0Ia$P�ԯ%J�Vz���<�iL�k��.v��*:����-�;��&���-�ʙ*��"Osتs�g&=�h���0v���SѤ��􇉀 [ȳ�_����p�7��	�L�_�N�ͷ�5���wȤC)Rs"�N�^&Xe�wE�ue�p��C�8lK<{j�f�\tl�D�N�_{ɚ�T�u�P�2}���ۢ�%Y�'c�$�pol�����E3%܄iA�2�}%��؆_�,7Z登-1�[Z�;���yvY�+1�`��ٳ�R!�P���庅)6�>������D��gL�#E��kx	֏�U"�s�A��*���o��n?o;��J�{Ulp�>=v�5qp���T�"I�����+R6�`���7�o矹��ف�� �.�D�!�)��ޔr ��ؗF�^��*"�}�>6XRh͐.Tz�\S�6���_y}[@�q3l�X�nq��@����}��bd�ֱnl�Y'i��4�������5RT��VwR=n�ǥ!� (�����)ɩ״L�?���sKFi�sM�PZ�ĀvW%�s�i��:���c�Ɍ�qG:h��x<��B���&�P{��t��M^�����,{V�*��z�ͣ]�yZ��I2Is&h�W��ͨ4~*E��EXά�	?U�W�ꔠd�:ܣ.��Bħ���"F��Qd��/e��Kt`�a�����@;m(�o3~�I��j9 �:����3��K���^�N�_tsF�M�|6���7Ζ �����pd�۔w9�de���p݉��P�($SL�^ͪ���A���ec��PG�W8��U-�m�hn|������L��`	��o1)�<p̷�d/�i>�;`iO�����մR۽�a��Ϗs
H�ӹ�I���z���J^��U���NmR��D�S�����Q�/�X�ԭ�9gA+�]��K���VZ��*�-����<OvXN`��l��{�*_zE��=$C�0��t�@�b��T)�;"�wsH�r+�(P4��G�K�H�J�e�귶�R������#S0��m�P�1��`o�@���$�����JҠ�u4��I���@'��X r*��H��T��3���r��A0(�n����{L�NS�C���.@l ��M�Pxj�#�#�re��_R Ϥ��ȋ�����صj|:�O�@NK��c�X�<eV_.i4�vy���I~|�� ��,��d`= V?6�#SSW�c��p>�TH�W�����|,��L��
#I��o�.JA8t�>�Y 
�}�~��`h���U�,�����.����J�s'� D_�����D�c�3,/� d�\}�3Itc�Vgٷ�\�0fBEGb�*�'#��iF����
�,tay�4r�H������=�Y��x�h��!��q�Q��2�*I��jF�>�牁�O�6o�q��Hu�U[RR�9�]���Bu=� �ɋ�0�6cS"6�֖��g��4%��(]�TB�r*�nku� i �A��C)U�J֥*/S᪢&�������4$�xȈԦ��e���a0�pI���^H��3��N�Q.Wܢv�fs�#���8@�K���D�!�V�w��\*���^"���?K?��][�ܫ�"�z����#�<��_ȶU�-
�ы�p��D��|��9�;�$��q�XZp���W�f�Dڟ�_>�l"�m����`��oy�ը��`�?K˞���d���Z����gnqj]5�-��ņ`������9κ�^t���qLG��}󫪃���^�+/Џ�=;�������ͬ���i���kqt]b-G�J�oj46��;��q�r�h��^l��M2q�8Jh<�^���X".�O����\�����ȌQ�$jR�i-:<�Y|旎\��oX������9y�EI����}Fǧ'i���w��m��7n�O�\�+=g����z��o\]JP"�w�� �G_�5��ɵ�x7�W�ȴ��zL�DȴE��f����F.�
�F*�e,���Yw����e��k؃=g���D�U��+`����fOmt&xA:�8��'�R�ku��fsN��u~��44��x&ҨͻKB��qw*U�89J�Ɛǎ�F���r��jz��3ᶞ�P�r�h�9SO�=5rԎ>��`Qsr�~Ȟ؛��N��3L���� '�=+ӻ��N*��y�%ȡ��
2��A9Zp�{-!ii�|m���V���i|r8K��Y��>OL�tv�ꪮa�U��f�:���<�y��������"o!�e�Ǯ�ߴM<[�X���ӕ����~��?���ek������ѯ�:�s�)�%�c����H�z)��{`�w�)8`��FKO߈��EMs��*����,S:��M�m�Y"qA�:�T��C�H"h��m�7B<m�O��^I��PZ�b!S��d|����f�
x�M��=�2���'��#�ffT<w�גyE��f�qƛ&)�Q,��Uc�vX�P�d���~���^��z�Eci�aŭ�bm#��Sg��z�;�ұ
�8#�"��V�ʨ�2�QS&�mάu6);Z�-KH�8MR_�c�H��Q��w�uH��)�%��<oz\QK0�=!�v��Z�M�18Yz��14l��Q��v4��?<��_Tz��n����x$����+�n)Ǜ����d��r�,bD"g�P �ߘ��J��ÌN���ER.�fN>��N�U&��?�����-6�O�� ���z�b��xY٫c���c� ϑa#a���ȼ�� Ks�u�^(D�����=�8��� �YK��T�oZ�b\�v:��E����Օ�ؽ��_#*Sij�=YC���.�����TԝBߠOܾ������xX����N��G�_�	ܗ̉A�9H���OUG1�f?�陶��#��11n��D ���a-�:�;z쩁�s�ͷ�|�?f�;��s{���O�.�)�E�fH0�d�q�����6fvU�gO���"�ޏɞ�\X\��P��k�w���okɽ:$�s����9jb�ܺB�����G~��S���D�ZbMͱ��{��=�7�-���PV\�s�.�WQ�I����ʫA�H ��+�]K���^��uL�R�ӯ�|Ť|���z������Zly���=
��hW5�R�+n�F�V�C�+�yG���M^�gQ��x��W�T����9�_.h�بi ��1�!K�V��P�\M�!a��S�a�t0^�M0��)�$.�3_�񨴗L�AD�8�7�2��!0�lu�����|��q�q{aU�sK�ɨ��m��og"�D\c����<@�('����N�!G�y��,��D$X�	x
�8i�B�=�F𬗻���m�s�2.M9v�e�܌�I9A4(ʸn�ۄ�R��k���=m~$�z�j��1��ލ��T2���t��ǐ�AME>p&�����|����l��oփ�
��bP�An>$��aX�����z��@"���O�>v���v�Ʈz@ZH�<��uâ�<���� �ʎ�ͤ��_9���r���U��X� q[m7�	�0P������Sh��!/@�`�!�J��T����wY�{���3L�	��=����D�~��K�U�Mg��4~w��+Ev_;&�D�����\���a��?� J4����	�B�mF�k���h��]mrN��� :���!��@3��Ȉ���}��"�{3���J�H��t�zݭ��0`�}�H+}�c>�q5WHZ}fJ!���u)���%ʚ������7K�K���X��E@'I�	�d��xHb�Q˘l�
 2%0/�?%7l���N/�ma\թ𫠡���W\~�D�"\Y/<+<�k�ʤ�M�MI�}��үU3�6U��Eຈ��g@�b��Z�6U\���bޭ�J��{�d���.ã�[w(�����.W�ZzȸE5Y([~|����vhPK��;�-�Z6hpZd�����@�t���DR����*"V.�r���|rzXߤ=0���>(|�+>i�Z6=�Q��g�S�4⠥�L�"�O�Yj*)�C���9�s�i�jb��*�@K1�V��+��j:��0�<�5����E��ƚ��y%��� b_[F/|a-IY?�P�h�KA�����y\Q�s��cg�0���/��f��ϧ��w���` x�vL����f͇�g�̻��`2���Û쯽�??�H��:���_s}np~�����?��scp�4�'T�%
0S�B@hH�*Y[��2�^�]K�xv���z�DL쑟`�d��%�`_�	��7�X�a.a0���)�t�~Y�F3M�)ȶ����){O5)v�Ǔx&)ղ�RAO�����{� #�Z�:�װ�"Iޒ����\�Ӣ��;Zj��|�ՎReݖ�B�K���<"�-��|���ѿ@HS��Å��SL�%#�(�Y�	0,Ż�;��"���Q� O'�0�FQ��Љ���={�<�|��<D&WP,�eL��>��T�{��sM�g(��w�rM���T"����q�a�4�G7D�HҪ���[ .��\�юL�I�a�gN��Cc�{|FS҈���l���C/૊��9�Z��B��8���p
*�V]����W�~��z�i3��Շc� ���oYo�ʘzf��O�ت�9ތ'�!i\:���v���,�0�Q
�� A�MEο�q��/D�n���? N�Z�G����{7�~-}3�A����	ˠ��PT�0J�{6��<}X
3S�����2�u�  ���Z#U����7��,;%�
�[e��ݝ�U�"�r߃�M�4��'gP�s0}��*p��>>L9X��In���R�#������ad� \ʃ��4�zɼY��V��2,���s�`����hq�C:?��2��l07��k�:	��2��	�g�"�'�:��\�P�^^�fp� ���n�y	v�um��y=�W{5%��<��
\<٥2Ҧr���y�@6_�|e�B���Q�%��NMR�2�Ajl��h%*�(�*�\�<wFI��[����Y�FC��QYwE�����[%�3�M~i��X-j#�Ǽ�>�o�9�1 =e���-P�	�X�e	=/��	�?ٳ�_�ޞS�·�G`Pmi�q�@��#�u`^1pƈ��_�?�R4ɑ 2;Țc0օ�mI���{w��}d豐�yD��m2Vu 4nǂ���1J���(�oU�s���}�����+�����o���p႖�:dL^�'�`�F˳#0�v>xA|�*����m��!�rc^B4����>�cA�kムߌן��}��.[.XN�m��`�l^�-q����P�6b����m�|�%�$�>���(�y�3�\�0�>�Ǹ���J��K5��O����چD�u�i��3~�LY��ԒH�k	����&�����	|R�m�1J���V�Ɖ�ހQ��|ى�����{�u�S�����ϳ�M*c���.��g$�9&�ǅ��.��.`j��m���_�Ra=�+����I^�2n9��+'ݷ�Rxd�B�=���sM�U�� mٓx�&$L�c�ټ�4�����V��ڒ=�y_�	��K[[q���0-�����7��<�e{:�~���^{c�g9Ƕ��OK���yn�Q��s���Ej�& ��h�2�B�4ʺ�f��q�y��*���8#K�����hp��wt8o��=C��������?^X�������vC�C�/ʌùQ� ��Y�c-�"#>� #�$~��`*A���G[3N�G���Yvu�e�.�%�����>	���SkJdo.oY�]5��wVC���&���T'܊�y�`ȸ�C�/���c�ct^��q�<X� ���p��& �Bzܟ���8Tkh���TG��Ü:p�A�����wH�f������"v)��Q"�1���(��I:SJ._Ǉw�*	��>Ė:��s�&K����pNI�_�6�ay�3���<>	׺���N<��/lM��ۨ �`q���C �I�_ ��$J��C�i��i�ؘ�}���������������[m�W�[�%���l�@�X�+�;�Rkǘ�#U��6�8_}�?{��c��վ�	�*l
*u��8S�����XL�˶!Ғ�.1=b�4�׶��%�m˒�j L�+��?�� �|&q�j�a���u(���Mv}�#���3�+�~�xR0l_fA��|�E�&#"��|��	�հ쐿?ِdA\n���7%r'z�z�XH��I���ꗘ�JG�N��z�cv�?���Ѷ ��l����O��|Qn�/���麎8֓����o���`�sԔt�,��ɸ�H����P�'=��#�wu@����f����#_�{����S�v#����APy�1�vFt���l����#��Yem.�HU!+�He�3���eB�j��?Ǜ4�RNf�1-&������f������p��(� iY+6���.�f<��\
Nf����k?b_�Ύ���nD�kX�ڵ��}q��%�����3[� ���lq��{����Z�=hc
|U�����M6��!�I���nx�@�tv��wL��b���1(Zd�b,�TRo	�z����D�"p�2�2�ͬa���h/�/��R�j�j)a88�V�3[A=&=J��)|v-�d Q������%��å}��!�T�#�Uպ�۰X�K����Y��
C<��w4=��f�0{�����`�B/Ԛ�Ut�TM@���R���U(~���<w�m�uSr�i��g�l�!ǹ�wӔb�K�qj���$��X����Ll�s�%�D�5b�a�<h��/`8d�E��.���w�X]�TG�k�CP5�m��m%�❓�7�<��.#�|�2����<�X���n_��f��y."�K\��f��ݓ�;�ڊipU�C�^r"z��~G�jq���9,`(�ު�Ma`a��*GtV��fQ�3c���2�δ���l%�O��KJ��U��5	�S �z���O�� �K���8��j��L��L8ha�-��b<��i�m����cBɾ��$ш��u<bCu�vć�p h��)���	<U;���7�!�����~�g��ϿMY��jv�hI:�~.NL���ZRCB�Hs(�����,��FA�u���S`�#[%-���qtz����i&�9�-[��@s���_}mN�"N��G�3,��;�Y�g�S��&��𱫽cX;ӻZ��?�������'O�W��Y��\9�u�=_�^ \���+K ��w�\k���r�[f ��ݼ�Y�%6a�]����.����^�����P�$�?�$���A$�ĞѾ���R��[�He�c�6�H�`�އ��GN��u[>W�ɥ��E'ʷTm�[�ߓ�婹���H9Py`�E���Ų2�9��e�E ���+m���K�����D�NEO�%=�P�e�+�
����H�8���Q���tϠ�)�ȚRrg�\1��G��T���2�r4n:7{�}�lQ�È�A'�O�^�Uq�՜l%%Q'Ph�J#���x��	�f���:!�9��������]u.x&�����p&�]��@ּxJ�_	���*b$���}s�m�9lrUM��(Ě;��'ia��8���U��U�BLK<|�=�����E�]�|efw��!�:��ۺ��pH᳚�y\Y�5���'�4�X�x~�x�D�/%S��n�^?g��Ѱ
0�i��9�͵?lB���8�V��L�ֆ�3no�:���Nh�.�CT�E[6#�7��͑�'��L|�#���$^��x�֌v]vI��,��(�==ڋ�0R!���I.G��@]m	�I�Ҿ�x)(na��l�~tU�88z�-`�`��wRU@Q��mIņvu������(U�m[SS<���d�Oو=��N�|��-�Q��f���j��vg3�K�>���C�β�0L���ܯ0��G��bq�������Y���S8��r趫C��zO&R.v��k���Ia���k�(��U"�FK{J���$�b7�k-�k ���=��6uC>�Zb{qPkϐ�x�_v����qȢ5�H��J����d�tx8�ې�)�'�ʘBOLA�qAL�Zc��W���au ��!��pe8����	�ݴd[jX���~=o u�����IS���IP0-Žb��hI�����%���o��+������^���򟇂�]:��2�]f��{)��-�������I�.;���{d�?4�� ���� j0����o^bَcC���9��JE�}՘�?��)#��q^~�#�p<4*���_\��T�ˋhnt��B�,�!]����8�h�|�"�
7_�Lg0�f$�йQ�"bz*�Y��o�3uo��V�^`�"NŠnҘ#��Ѕu/CŚ����-6��֝�6zw�NU���3��lM�|�Ě�CL������`)�Q���0Ĭ��i��[��	Ǡ_�DA5�
&әaY6h����gҊ�[~ٷ@d<E�N>H��g��
w���W��G�Yeu�禚��1�m�F��T���x��
� [�10�����m&����1�&�Y��`Z�%�?��������
i�c���]���hVp
+���˩ � 𲹔����5���(�b�������r_� =�aH-����p3$��^� 	��I���Q2׮������mih���f�
m���֏��+6�v�u	ß����qo�����u���nn�����؊ʙ�U�a����+����X�,����;���ns1T�9ᡬ�֬4˃ ?p"�V�
Y�3Z��b�P;��;2�Ry�2MT[�c����:�`���&�3M����}�W�1���8|OD��鰉K�p�ק}��H�$L�@��1�8�<�]�G�~i
jq�B�d�����nLqŹI��*VE
	Gw͇2��Sگ�Vփ�F��%�ŧ���{�C��K�Or�0�����C~�D���{yg����穡�D�󌰺���<�<�5�`�x���Gc<��������iMG��N?�&��F������rE�-��]o�\<L��0�Dc�M�xdU��ܴ�aQ�6��D��x����|z���,�cDĩ�����q_���鸞R��@���-���<�:�dL~�
������j�H$7�c���P�I�k<�F�	��I��6���ʿ�2��r%�r�v��ѩ�=7����pX0&�̌,կ����:�r��R��m��Agg}2��������։?~���nfh�e��z�K}Գ��}�������ō�;*P�\�y9{v��E� z4�B�2�J�O� W;��>��j���:��ȸ08]A��٨���fd_8�����Ku��X<��2ف\�+@�,c_Z�����D1�ĭ���*f3,��*�xn����URa<���4G��K@��1g=���L2�����^L�$b5�p�;��[E�7�r1��؇�V�^��	��2=]��h��C+���d�+���{ԕYx��d�5,^�\���Z����&��Ü��+�Q����Fq���s	_�~��؃��hYV���C�	���5�q�ҧ�Eb�����$)T7_+� !����v\��G�����"�w4��C�s�*ҚAeF{�\�ՙFWL+��(�G��U�:PE�M�T�Z��8e��Q`��ܼ�����Β3#��i���ҭd�8/PNuc~�=!儹�O\$��d�/{��Y�/X|��L�K���.�t:~���d���
�du!A���_������T��j�O1�e���v�`D�xj��J>��@0�'i��3��F�~`���#�𶂅�=�-��e�Ĉ�2����(�j
�51bm�P��~����V�D�ð�r�J�� �u=��/��Zy�sO�Ј��*�\Z,��@~���SQc��K��K�$��	�ǫ ��:�+(��9��m�V۾<i�<�_���|#�	�Z�ZE�J۳��Z�m��y&��%�>=?���:�G�3�RT�z(�<�s&j�l�,��TWD���*�6!iq���[6�o�>wK����w��P_���0d5�S�Z�����s߿��/h�4%s�`)��OT��� �̄�N�F++-?�s�@A%�C/��7_�� 2�o&�0��YB�I��ު�n�wa?���'a�L;ؘ�HF�7��ަh�b�Ĉs�H�v6��o�3��Ӹ��x��6��|���>�D'nҫ����>�9�pQ~��0�a������^���4w�s(�/{�%g� !>��|��˜Rf���,��W*oW� ��.?���P��1�?p���',���d���Gmm0[v������T�v̘�b�B���J�N�79��g��N�o�'`��oر�~�%^�k6����U�%�N���^�p�jN�VIQ�hD
J��+}�7@J�;�u��*I��M� ��`�'��杖����LNǜ�M.9�}�`b^�)�x	�����Ͽa&MHYfتʒ_���%0�ι�W�х2��,�/���e��(��?�f��ǘD7b"�elM�Pl!�'06C�I�'=6��B4O0tN�~v��
���{x�O[_�fk�6��-�:�fؖ�~�ʒg���<���Wb̢�jzsf4�W�6��JI(���AҜ�mhY?�=7��������"2bP���x��Xj�ԟ�"�n�%���[M$�u��8�&���'�HF�~C��E3�t�O�k�fjp �����җN�t*O󠨲Ӏ���r�e���Нx}T=˕�#���2�d�ѐ��D'^�+E��Rz�9�8���&����e�]D�@M���	��� �X����;Cf�IޅS"�_R�P�K���T�y^��`�E�M�-�.��𷉺���a�^!IA�J����IH���N�ga�a�	�).� ¹rCU>���0�ԫ����u���{r�I�����2I� h�Z����(��W�ȶ��X���}�[�,s�Paul̝8@�����bYIUW��q����Y��ԯw�^����fN.+�9�mp��t!Y���jM��#B�BN
sځD5$�X�-=���vv\Bx��JJٸ��,�xW�APg���ǟ�$B6�N;�0p6Nx�A3�M2�T״L9]��\�ǁ.��t+������Џ9&�_	j�<�"�: -��g�l<�3���!���ί8��M������i�:�
�������K
>�	� j�qn6)X���#���3����G�G�Sw"=PR!k��:�=
����"уm)�j@�]S�����[d�{_k9�U{UB�$����Hԧ�u����QwS�� .���j߂@ar[��I��>A秐�9&^�1=�k��Jr֊��`�"/����'�/��