��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ�������������(�/�&kff�_���#~�+J�p�y�_0? �^/$2) e�Av�!8=��1�G�$,
�Y��Vb��3AIy����%G	��h�^d�+��F?�]�F#�G]q��x6_7 ���"c����(K��~E6��;��DcX�Du��:&NP�����C���mL�Wg��Y���퓾��c��T�"���UӾp����ú(;l�#�����_�ő�d��ň.�#3��iՓ�4��HVd�{����μ�!	!Ս.J���?Ӵ�ޭ�e_\�^q������g�,�ᫍdBV�`f��"?�6�Z��]�غ~^�( ��~��X�D�u=o�W�����^h��	��&%
��]#�si�%%0��C��N�q��E����n��m�������A�絶r�@y�G򑴒k̈n�V�~��=�]���ψ�ƅY?E����2����">y]�b��6�J7ԃj��v���S+	����	k컺�^Xt`���M�7H��t��싕��U���5���ֵ��D��Ң��{�ja`#�_�rp�#��v�������|���&^���ؼ�4c�����6��8�d���OT�٧J5z���B�F�jRk��Ri2Q{��ι8�j������ߢ��w��4|�m$g��A����O/�c����k��β ��X\Q�@�Z��rk�� n�w�5u˙��NǓ��f�2TW�y-a�]5ڃ?��:q�)���d�}4����#��̳M���)�ԏz���w�yqX�AԆ;�O:
�f�N�~$z����  n��,��
����C�}vλ���9p����2���&F�D��ε�M��0߲��%�q����4��%�u�g��.R���ub�9
�1��1m"o6A���y�Abf:ױ9k�Q�ƌy�7�f..����6��t��T=�brU(`��~�4~[�� e��{c��@��Ӽ���r)kR�C^�+��$�o	d]��v��4ܿ,���'�kM'�r$��7&�d�*Z_��*d��3�v��_7WE�D"V���������s�3����~���Ndǈ��d�N9	�k��E� C:��y�.�E�'�y�A�{�6�k�h1Y@h<-E#'���z�>n�Ug�?4���h�G����]Vk�n���\V u�I�%B`-S$��B��"���vGP����F?Wi�����J��o�m�x
\;��޼�*5���h������*������7��3n�_���oj��g�~�L�	� ��B��Vyd����3�m�E�Y����˽2��b]&�sQ#ŀ���8S�� zu	?G�	�5�}zA&Ƿ���X�Ň�9��������H|C�[�a��6�ee���W��_�tkO�'Y�![L�eVf����<�͒G?x
ق�<��=	
m#�w���F��N狗�_=����d>6Pl�(�w��f}���4����?�;����x�WwK�5O^�;��X��skK����P��Gi�4�b��0��C)�N�r_�!ew!��c6�w��LA���{C�,��mFYr"�lJ$.�7�ǜ��w޶^R��0����BO�e���R$��H��hYbjj�!�A�]�{�s#�|�J�Y�����^��])�El����� D�n�X@BY���a�i��˃Ma0"��w�"_{�l���R�D�,{�1գgc�����)8�B��*4q�fkƬ(*� Y{1�Z����g�l��vh�j����x=G�i�a'����ҫݳ�.X��N�m��֋Ƥ/�$��<YC@S�|z��AXQ��أU��S֬�Hv�Dwa=���H �J���5��6���w=�T� �Rb�v~q u���ؗuz�ez�����$v�ӵ6�l|m�E��$h`I��l�|��H�d��ȲV��GN=�6?�c�a�j
�����5<�$ž�v����俻�H��j���<�=oi�UD��&S8�4��4���'m�/�ʁ� ��J��(3�=���!�cV�������X��>Ub��-��v�Ԫ�*;d	�J��ܷ���.HUW��vóg ��=���(�;��K/���Ϗ[�7Ua4aP�ʄ�o!;-��xAO��<�,?(3$;m�N��3y�߹3�4{��kw�1���@%�S�o�����ŕ�`���o�!�idK��?�T7����&��0=�
\�j��&�lpm.E'�<KA��j�Ni�螈z�5�Э�ɢEb��*ג1�6w����Kȳ{��9/ȍ�8YhO氤p�ǩ)�c�x��sM�ڸ�_ǹ'_�O��� ��撙nRҮ���tzX� EQ��>밿�k��{7��-��PX�����D��	�V�?T��6��@nO���!7��)b��U�	�O�I�c3Ϊ:]fk�б��t�����ٛ1I})�|��[�"��ܗ	�����P{�ɣQJs�5����Ud�%����@�ۜ�opW�"�y�Kz{$Z)�\+�٩#����F��g�Z��$8��̅���k??{kxls��P�Rh!�悿�V'�gW���w�����r��Ֆ��@��a^��HN��g�\���1A�Ȕ���8alⓨ̑Av��V��-�s���1��W>ŭ�� l������3~4���Z��wD��Fa_���E�������án��b��:�"]��_�-h�KQ�f�J�sx�ހ�q��|�;P8[�CxYh��!%! A�f�T:E��n���6s�s�6��T�� �eŘ��*�?�SzŞ��r<�A�7��֛�dp�?�{RZݑ�􊤬�qI���x�*�R����i<|�K����5�5_��CfV��b�T��BZ���Q�(��g��^��P���~���w���r �����{�\Ȇ��M�gu��ҖA �����~5
���رl�n#��Z��"�-De[�离}K�S6|�59��ݴ��7EB t�t��f1��T��e�����CӮ("Ob�����	dte��\�}ݮWg�b8In4�s�C�gJe��$��Y}y�3Q�iu�#i[_�����cǉ��R� ������b�JK���uNi��j$ ��R��W!��w����q=���	y��Q�h%���t�~:E�M���\���M�0WyT�����S��y��&C��]ko�,b��鬅�֨�\�Hl��H�n-�?c(��h�RU.{���?�@����J g	�)\|�~������IDw�L���7P?i������:Fל�2�QN&*�5c�Iၞl��ߛ�R ��F[>P���'k̼���Bt�Xl��W������A<�}d��<C�O = ,�Up���l{�_�r�K�J�tW�q��n��9%E[[���X���9$��uP�)��Q�יaC�I�qN�0IW��RLt�g�C+��R��T�Y�{�,���[�F��,��xmu�������@��_3���j,t������W/m�yҬ �.e��,?\�:c�O�߯K�.�$�x�T�y��j�_E	�p��rq"=y=)��:u4m��t�����^���Ë�0V�@��r�v�Dcu�����e���' ����HL�'|�� �8{�z��E�������!V��+;y��z���H�����8Q�&k H�S��'�P��_���v]EAG��:#�n�	CtV�[�U��]���ק�aYH�@K^_�z  .j����>�1�~���
����)J0�w�0;������ �O]�Msb�k6��^d��S8zb@::�@k��D7E}��	���F&�>�@-}���[C��U$iޤ�ì����r��e�̷������!	��1Ī�x*�"����^���E��%i ��Ğ��+��g�rՋ��\���:�ڥG �٤[FA����%B���T��H#�'iZ����uyL�����B���-8>�A�B�S	���G2��6G]Uo1tے�������7hZ�4�K��z��p�[���L�¨J�s�)�z[�d�2`~SF�T,h4�CWڎ�G�Q�!+n�$;���s ��:ր'~պ"� ��믗�#[����^g���z5�)�4	���/�dl�=°o���e�YK��'��,��N�?��ɿZ���m���!6oSD��Fk��jw6�+*������R-�S>���?Ud��sE��c��Ug9��I�L�=��u�ł[4���f̾VlM�`�9Y;�[s�����c�B$����\s�)s5kDr��:�j>�u�de3�Z|�f6�Ҳd|o�[:�+��� ffJI�|U�|F(h��������hH�j�"�ڮ�,�f�҆|9�)��&3M�+A��!|@�Up�s������H�� p}�G)���E (�
&�`2���q{=\����dr���r����,.@gv�Z��"6�d�U֖� $I��aQ��*s�PJa��}���np��/0W�\>7���"lc����;����l��[.�m"���9��L}����X#�v�ro�@�v�.�6B��:O�+7�!���˶\m�\؞�'�I��P�4�=W�2�WpI1�<T�@��J��K���x�/��U���7#�*��ɾ��X$缝��֐�H��\s�^��>(1�q���`�7��i�q<��_��ꈵ,�@���߸�Q磓/�1�2�u��!�ŉ3���Hr� 0�;�S�^��D+�ȅ�k���o��\.	�Lݴ7h��z0��̣�v򧥍DBX��}׋��k^��{�ͮ?^� M[��]⻠Ӭ�mԟ���`\/j��F5pU��|�����%�RCH�t�� wtrk���*ƏK�Pۆ>��BfL�R;څ�Z�CLQj7f�h��%fe��ܦ�PG�!�<��#a&���%?�ՙ��o`�s�`����r���y�0���&��Tÿ��7���t$(�%�x��o�e��;�8[�O�P@���p'ɚ���~����$}��S����:� ��.���7���K{���,�����B��S������" ]5��
�]��c���^����Zz'������7흐�`y߹f����{���W�$��J\]���y�a�E�@��I���Ht��W�, ���m��~a�`ⴳ�/�ǜ��˂D4A��e��F��ő>1��M�|���jVõH�y�LT�ςy^���|A���{�3$��������}+g�g�l�;K������L�>h�+���n�8�!Q���2jЉbڨ��j
���G^������Qsr-����?/laY��¯��rd�������"ޝ ��w:�T|@���H��_^ج�M��*E����7L��"�C̲�uF�l��]�Y�L֒&|۶�,yO�#�"L�����񷊚�԰NUn�âu԰ᰘM�e�6%��A��T�H��%��ج�;ވ_�_�%�!a#!i�(�
��ǚ��ɱ�ZcE%
�$�L��>A�-��?����7�?��B���\!}���ֳ�����F��cp�
�|���9`���]8+s�b*L:��p(&k�s��v���C�����*�f����;�R;�^�Uq�!������y]zU���N )�Vǀ�Ժ�+x[��'C2�60�)+V[hV{�v��G��?1X�?�BѮ��d�&��$mH�Q�A�x)hI����٣��-
�^;��U�"����Z�z�>���k�׵!����=��������f��Y1?�W����]%o7Ǘ<��ާ�aDO�=��Y���,�:< ��d<j�r�V����Y�ˬ>�����b�V�qn]����,\<�f)����^��0�TsK���oOb�D�Z���y��@?H$���a�<�q��@���� ������7������0�Q�@8���<��y.i]'t���3a<�K�s��+��b���9U���_A{!���}�-JM}����z\_��/��-dx`R��̤wy�DޭWخ���p��ؽR��|����<v��7w��Y�*
�k-zvU�9�lV�#N�9÷�9�-�͑Z^]��I�V�G��v�|e�Ûrj���\E���,��$��Ժ�d�mT��e�����ꣽ`�j���1�W��838[����(굺,Ǽީ��l�f��2+I1�6	!�����U�@f"��/��]A�G�BzA�l��S��x%D�Vm=�����7�{�=;	YP�r�2$�����Wt�q��%=&)�aL�.�S �{���]�-[�h���=�xOo�2e���m��"��ɕ[��d{�h(�re`��mnJ�	��l��j a�֓��`�`/����S�GL���_���Vs2ue�]����3j�[Ei��7:tU�ܽ����-���:S�Ag$��}���;r`2P�'),���'�:���aC�G���M8@��|`�����ۂ��CP�g�3f�ЭڕE��U��)S���e�{Q1x)$Xt:��9=3���T��9��������%�|'�
Yw��敭٥�1�}��8 n
�7���l}Mf��mm6��A,L������*V_}z�P��O�	���W����$8k���Urh����O�Mͥ,+j~79p�ٔ�/�̾�R��V"c��\�,�G��{W؅��%u�{Y��[� �N�>�b&��F����]��o�p���wW�=�2WFTa��dz���_E����:�~���5p�m��<E�G	iǭl0uq�M��2�g0�Pu9rX��B�j�7a���p�1��5������pu�b�7�$
v#V.&���y�U�����R~�j$ޯ*�K�q��L7�����o�h�����,��[J��$0KY����B�P.ѝ#�?kC�f�7*�~x���N>��8J��x���5� �U~DoE��'���w�J��\�����vÁI[��^2���O%���$t�n��ܯ_�h�P�%��@��Y�o4��gW%Y�*�Ct������'?������vI�vG"�wԥ��B�\��:�J�>ש������E�v��n�{��U;���f��$�[*T�F�x�̼�|�R��u�q�Gή�[$+�wz�� Q���]%�ɱ�y�[i}|�<�vE�16��.��|@��� |JZ�/�*�t��Q��_$x�e��=ձs:�YuD[ ����<���/߾�T&E_,�߻� `���� Jq'^]{fb5z�F:��H�$�X�?%����/����fE�6l����|��L7�H4����4F��BN��ua���7.�/��	#p�����,��ߴ�Ln�6uC_��=1���.��~��Q^ ?���K���ֲ_�u���b�vK���Z�f���U�je��͌@�Ԫ�%�t��Rߝr�F$��r��^�J���u=���'�?�����q�MX� ���0B��z�����V�L���q�F��t�ق�V�îTAo$��n*=�����f������V�9��uǟ�����H�_Y-�^dMm�	smE	�cbB��cKJ�������JZ����>���U`^d
`���Æ��]�D~�gf���M�z�j�������ӟ_��NP�B�r�^��7:�N\��_:����}�b��y�pT/��HiS`Kdh&��ު:��%?Q����ǲ5�w�)�6.o5طȄ��z��j�+X��X�}��.�>��j#�.������m5t�=J��BG`21��E����1�r�_�3X�g)��T�&nγ2�������7��J���M��߰DB�5GQSL��=�d�Xm-�@��:�̰�0����#F1H��m�.4KF{���Fh5���s�\�o����/�43�2<Jȝǖh��a�^Jv�� ��|���V�d�ޱv�;u���x�P����Ͱ(�'��9��R~�RR�1��Y����ڐ�V�� Y#�#�|g�aQ�R��%hd�O��@��ĜRxw>4W�¦�?C�����z�"��5��:\\�W�v�h�j����5w���	l��g��L�HDb�̂�0�A�Hl�4����$)���*�3���1?��AE��,xӯ����/�qU1�u]��]�XX��jdh�N 3!�� ��1==�;�����PT��ww8>좊mw	0cP��ڏ�S�8���$t������YM������ROXI�#�4Ψ8����с~qv�O���FnA�U{:[����F���=W��<��¯��@�ܕ+�Z�o���w�@��>N�N����%�I��龜BvJ]�lV������$�r��*e�$�n���;�M������>��/R�c�}�Ն�|����\������y�/eFv12<�M��'��yd�`Ρ��,��ָ�z�(�
��s�  {����M.�����2Xx�|MK�W%�������U�C#U���M�O�����]�4S�O��k�(��|�uEK
�GF`o�A�e��&���a�x�@s�_�s���,W8ո�[^%��!��l53LP�k�~��a�p@T���p�]������@ֆ3���V��%C B����Z�����t�����C�C��%cA�Р��=��ɳ\�wZTh��R��Dz�W��u�C����$v��%(��>n3����GU�V������P6��FBƳSD.��j7i�j.v��:"�Xdڪz��P�}#�vH��fgp/�*����ܡ���b������;��0#nL�O^1\��ю�_�jk�8��X�q�T�BEɰS�8�����w�f�w�6��L��*����+���+��+�D�tSX�D������X{�����)8C�0@��O�8,=VꂪCwq��ڇY�����,0< j6Q���ŏ~�4V���p?���̻���e�edrnЗC�A�ʽ�D�c�� �Fp�����5�؛��q���Q�E��j�q����l��	��#3Y���y&�GQVǝ��#�r4|�=�`ik���������] �rhnt��k����C@�����r���K������6�%���#y�>s T&(3q�YXWOE������ާ|h\>jD�{�rڠ7��Z�U:�
��8�}CvVs�>�s		^��S�}���\�q��9 %�#�5ѭdk���g�&I �`AJ����:b8m��6���,������T�\�\a�Րx��[GV��(�c֍s���,�K1X��"��.x���,G�HzM�g�[���ɴ2훤2�*D"9�0�SoH�톄A��G@�@���X��.�_Y�	��I����-|��k���3y_�0L{p��O;�X��8Xh���G Ò40�3Bx������	J˳d����]���"ޟ	i��6�"��#62�g��z��P�%�ҧ�������u�F)
��+&rpĥ��=0{�?d��C�}�)�?���:�	�'�w�����E�y&�~u������Ψ��%f_�[8^t/��'<R�d�N��NX���S����3�t�T{��'�ĭ#�*�م��~E��[���.�z/R�_��_���Oڃ`9��{�L`�<)���|]�Ǝ!�~,�S�[�d��d�:�@��L���#e�!nko�W�	���@�_u�48��Q��aNo��QO�)��~X�f��6��/���+��bg�Mkn�i]�,�wF�=�7B�*�����<=��A]��`��ɫ����k��E	C�V��+���>���ͷ�n��^r��ᚶ|Y���j���K��m� ߔ�h"N9f��q瞘��7q�P�ʼ������~'���|�X�>�֩U)��w�~���^__��{�_�
��W�XqוHP��$a��"
u�������`��� ��gz�Ԣ���'�saџ����.�eC֣qS��Xo&���[!��Q�y�eإ����,���\5�|���E�o���?>�[� &J]���|�^X1$H9F)����_R����_��
a\�ԝP�u�T~���Ny��{굛�<mS��bo��ȴ�T��?���V���l�?�6��"GE�	+�; 1f���E�js�7I�_��]R��?��������a��&T�@�j૜`mOhW�Ү��{�s+Mq:�X�d3��O}%�y��*G��Mu#S�I�V_��y���>�瑂jI�	ds�����&�9?��GE�K[g�����c�,�`q��c�_�;�nH�*nJKq������ p�'�ހ��b�"�EK�����*q�⎬�_r7mh�<�Y��?z�s �SJ�R6RC���b��2-�fx��������¡����hR��)�ˁ��E�ٸN��I�O�h_��\����'ғB��{k��l@� ;� �|\��V8\]�<�W�h��Yuc���c}�YOX��0�x��2zt+f�T&t�e]�7�A��>2�L}�!^~�VC5�e�8���	\��v���#�@}�k9�dE�?"g.v�H�n�$3�hY��x����2��`I��qʿ���
T�[~S���4�.F�9�r�c>U�\\K�T�ޝ����ӾU�q�SB�,�,��^�
ĩG�Gt����)��
���*�q������N��j��.&����@'�<:5B�cܻ���/N~y�7��,��J�9~�������ݙ����LZ�~����-�t�)0�V�����/��z�W}���.��w�I'I���`�K��b��ik�~OeJp�_�3˹�u\��\ǯ�Z"mW+��FܘR/
ؔ��;}�+�+s}�[���w��~�Y��W��(C�<M�q����P�D�u5���{i(�O�n���}kW�B�I����W�.tPt���`�_C+��p+�g��^ j�m���_A��ㅙSM����"-^��_����}�W���s.��z�$�.�9�F����t�P\���X	���G�#���z�@��� g�@~�����1�N�R�xL~s?�z''� l���փ�2j�Lk{��g�W��G� Բ����:�/�1�ىB.�f��X_
�nȳ"0�OA���I�,���ZE(�$c��!#/��d-�1�m�2�c>��q-u"��^�h��{��ӝ;�&���#1�ˋ����,鐟�:�7����@=/�׭�ͅ�(We��<�n�RAa�SHԀv6��YT�bHH�D�g�f�g�2c����Ԍ�����d���B������� ���ei��mXv"�v#v|dE	 -5G�`���V.j��dS���H�6\��d,�x���%ހ@��"O	��zG��U^Q#O�[�
X��r�H�+1����T�����19�q��[/�ܜ�)�J�x'��2jӿ:۲���߱f���
�U�f�"u�>�`*�W�g1g80��dC�9�[���c0If\|V#^C|� hfƀ����X��Y�����*��0�"J�Ν\����T��O�9Ow����&p""�κ����:/r�#��9g��[�k����C�D�Z]��]
�j9|�$p�