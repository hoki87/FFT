��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ���������y@f�~?A7v*�2%�*��2�p�9��B��*����5���E���� =ǣ�І�c���v��t�2bX�C5�8 �bQ�J����d��v��!ԷE�����+V?6���nxXw'�m�>B'�Q��˪}�* �j=�Q�ڴ���Ia-�4L3�@T�~���z~tj^���B}�\:��^�H۳e����h�q�H�s�P�:�Yƥ���+�+	{f������F֠s�����N���ϒ��]�F�'�O������{�lI>1�3Y���T��H�*޼  L��/�K�>�x�r'H������=R�PsD�N}q �o�3)�*v;P˓]]S=Q�> \	<�Q*n���ya��_>�R(��fN��A��I-�����!�����CWA�������u)gt�Z
fJ�sӘ\���,�q���1�+��9�yv[�8�����k7��M�ܝ�s	v��%.�(D����k@�ǰ�
݉�[^�k�K���[����g|Q%�wT����B8�κMJ];�x�rna��P���gh[a�	�w�;��ɹ܏t�\�z�9��}�'��]c<0��B$.��m6ґ;&yq�N����(+��<xΉ������2��Pi>�!��;�[��8�M�y4�p��P7V�ɾ��'�s&���tE�Ҋ�����3t
�͵;��$��C�\C*�\}p̝�ryo(]�̉m#?�7���+ƹ��pƆ�f��5r�����ҳ��6�#�}\%Uc;��������vπb���'=�Ѳ�}u7�;\�>�"{%<�	��e�����>fn�6���7��*��!�����7S\Z&zV���7�wI��w�e��T�u���a�^�,����1���=�8�J��L���)�#��T�x7%� sDg`�����Z"@���"�̇�
!���n�ͫ�34e���Z'�+{�`;�����̾��u�P$t'ٗ�2����3��5l��^B�M�nc^!Z�T\��r��\���w�+eP8j�]j;���]G b��[3�S�S�u�@�ƙq�)�٣q����nƓ��4���Ϣ�b�f@F�Jf����W�'����d��>E,�M�˸L��-_�a�H/8R�8�a���;呻>w��l�n��<	1g�|�'�)��v]�i�Gq�H�ޖ�0�0��;������@��\-�@�)�!�%Ѱ7�8�'E�V��}�4XK��������2��+��V���I��g��7^��	0p�^��<-�/�W� �+'�������Al�C��~SֲF��̛w�m�\qMS��w{҃Lô�Φ�6�/}6J���]c 	�mo��`h
�aJ�HAL�"�P[I&) ��5�<bĥ ܄ �K���m� �$�����)e���AV���	z��\#0�+G��h�4�����
5#� �ڧ��%��q�F8Sa~+h/���T��iTѕ�\��ߛ�L�<�1f$��9���+�!�����z"���>bBmA	͠j?�/{Φ ��u���	�%
���o1�+~���Nw��.���vi�T]3��G2+��hm	n���Iq�9n/A�,��6�����Q6R�t�QZ��IPo��l$�=�O�d���A�����(��*������Wǧ�V�u������Ξ՟�w��!�ϳ�l�Q|�5��~��!\;�`*%1>k�V廯�������0E��ogf��x� |V��ݾ��c���Jnn?�w��К��[��IChȁݯQ�#m~��a�T-*�B��.�K���N棾~��F��@o�{�4��#��4���Oa���K���i�Aߊ��4m9���K9�7y2X��/�!��Sٜt�n{�e��^s{E���}��~f�ѯ��}�LsPؒ����?���lW�;0X͜��0����2|�R:opT���5��{#��k0[0�x�wZ��j�.�5Q�&���;V!Kɖ.	�5WQ�u�����h���39#�ή<5kȘ"գ�3��pz� ��'��O��76�3�/�������n�nx�9�OU�	���}hV:@��kv n!�P%o�j1�N�Fyk��|
�e/U��+�R�6��U�@~��G�E
>5��ĀlUm�21c5�Ŧ���P2l����fKd�9[1U�
kLic��wL�ޚ{q�!o�V:��$b�^��0�7���X��N#��D�Ơ����@��	f�)�s��5��[>��r�J5�y�x؛�>)g�Na�W�f8x�/B��Ҁ�3:��n�+� ��dq�ճ:�q*X�1Ŵ�$%���!�o�6<³��������O��ć|��NV�P��@���p^�T���An�V��k0��s{^^�V�]�Ob�p��Q�8 ���� �a���4��*�Z��Jl@���N];"�X�f�(@��l�WASSL�X-��	�	�&�/��pa�]%?m��P�AgO3/���ն�`��4-�������÷]@�p��|d~[.-�P��NI��=��\�H���^��hv҈M���x��G����͞�4t�HMh�&�J�V�7P/č��T�y�E���}q�)�A���CԠ�7g�x��{���X�F��+*������r�i� �]�E~��[f�������GIU���)��|u�x�P�ݔԜ�I�A-��Gc�T�$�`9�[�n��� �
�'�r�9!jҨ(X�y��[:��	ñ;�,��6I".u��$���q����$��\ ���RxXf�W!8���a��ԅ�|�!kS	��V��)�nP�(C{��Q1H���0-�	��������bW�|��MR@ěɄ;��0�X.���K�`�X��"�#�R�.�=�}�AY�]�ș�d���x�Gd����'\��
�k��b�1$�/E�0����5<uC}_a�e�/��$Y�L	<s0��Z��TUוH�s���,�7�r%b�@xDJ��M^{L��Lr~�Y�I�9K��n���D�S���t���{�'b|9}x<��K���fa�'i���%h���z`�����F���r��ȷͽI�	�����?��W��b��SI�9u1�%��l����\��.&9���t7���a+:0���L��\=S2�S���e�g�t0Rѹ^�A�ԧK�C�{�|����Gâ
gK7D�Z�]@�7���&�vև��^K���ֽ���j���b�,8{���`�� �"t�W�0.�n��[e1��n.!�׃>,Ρ���x���IU��w/�u�9(X����>��n�T%���)6�F��`Sق���'6bei��22�>ĽD��b�I���}f>�!�>Y�GZ~�.�Ʒ�S�� 3�V�TA�vBfȼ����ޏ57 ����)$%���R�D�S��z�8T���%w?�D�Z�Z��͎Sep3�"�Q�++�{�(��/h?e�� ��f3�od����}��8X���L�S@�(�ޥ�X-ױ�&S�X՚����qh�.��(�l# 8Zc�u�ʫ�����U��/� �u��X�^)��&Y�;��z]|ܕ$�q)�ѫ ��L�b�E��%D=��sXy},��S+�C�,�C�sGR�t�b��[��#��i�`h��r�!+�5=��+����":�O0GV�x#G1����e[��k��"y�5���s����Ht��ߨs�F`�]��"�-���y�p�If�} ������$F4fF5�T��
Z��3��u�3����b���7X��e��GJ�v�'sC�|eW��o{3�Ϟ3�����I�Z�Лv芫�֯D�:ػ����Vײ�rb>�Ȱ�O~�y�^�T�T�rQDdN���o�~/�^p�5L��r�������Qޕ�C��T�8����".�a# �C9�� �a���ّm�{�2-;���������`��RV��x\M�?�]�����J_w]2�e���	g%B��.oUe�*�?�%��<VGt-��e!�@s�eT�,��s�E3Hh��Ru;�ah�\��ޤ{��c�~3]�V!��$2�����,���ɉ���l��2Y�!s��k-F�����ȧVşF�h��U�vR�w�VRʁ8�^��0�L9 ��)c�)"u�����:hӢ���j���u�?"�h�]q_X�x&0��D��n�?͸s���x���W�{�>�Hb�p}�6��1�w���ԏqi^,߷�ouB�6P>W�y�M0�%���ه5ޟ����c�ѧM��Q��;2���ij$q\������=��ӛ�F1��P�?Y����r�K���Z��.8����l+��5����������%	{�ιN� ��w�ɮ�c�1�YZ}�y�C�Mv�oQ�+���x�
;u�7�t	�xH����V�X�h�m�������`Э8��	��u���Sa5��?����t���(D�?+,ʿ��c���D)%#��IeIt���u��61�i���}g�.8�]u���I���1댚�25�R�_ofS2�dU�n�!.��5��K=9�j��U$��xb�>�RD�	.���,���	������
��Sd���$`�1�2�/?m�	M�do(�N��tv6�E a�����É��%�5䷶���	W
���kB���/�����<�q$�-cX:T��5`i�k��e�e��Sf�[ �,�"$�0Q*�;줬�^��dv����;�X����:�>fX������e�c?y��ؼ�ޑ��X9�`�4J�.v��S�jYlxx�S�>��+�1����1eO�K��d�N�(!�z���h3�NA���;�a�Y�m�̅S��]6�� ��h�����]F���I�v�%�\'��;��w�,��a+A�z`���}�2���+B,������"m^���I�uM��ν��He\<8��t�X�ån�Uܷw��!o����<���h��[>GIU���Ij医Q8�9'��^rD��$~�V;8�8:!̒"2t�@��,�q���u;�۪09+߭D�}{g�L�X��3;��v���V�����b͖j'ٛJ��~��v
��w�a����bݧ�S��ɞ�f���O%����T�t7��v��W3l��sLXq}�9�Q9vk�H��,��s�FHg7e?��9H�A��ωZ
��)`�����u�@�8*��gI^ٱR�lig�|��n��0}��M��p��Һك	����y+��!LQB����©���Q�X�M=��і[Ք>4c�����x��^E��)\9C3�=s3f�#/Uź�[�C�`��T��]�rkaW�~9��+ZK���鄶6d8���������yMЃ�[i�y|�>S' �cǳ���L�,�t[�f%�p<�2��D�[w�CPda|m�i��D�x�nz0���S��@�+UV���%j[�T�����g�0<��v���VB/�~�Hh��~�լ
�dIuڃ&CyD_xPFUr`�)�&j���=q]g�q`���w��?�e���Ed�|�W�qfh-3S��P�S!���:x�E�/	���ǹo�­�S[�j�"\��g��L�(T�dP����";�X�cP�_4Q�tU����)#��#��/�k�|���^S�ֺ2Hd}H<]u&#�\ {	�ʫo�^��-aǉ]w�72�`�99&�G��|&RgAI�6��"RV�l ��R�ڹYh�q�'b����n� �IĒ2l�h3)���7���\���J2]�������%�-L[[�@�-+�[:Jg�;����3;V;8k��oj�]K�*A����=�#�1���`��Li"@^=�y4�cG�M�'�!�>�O�ĕr���PGݾ?^��Iy���׷]K��mP����屌ZH̉(:p���b���NE�<š�.{e%�x�H+=�4�Bø�v>�Y�*�fC^�T�Z�VR�@��A
�I�{O9O\.B@|�R
a�16�.<�ܡ