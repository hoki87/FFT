��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#���������l��U�~�׏O����j9�PY���`T���x���s����uí������P��"��b%>�1eτy�<�gܰ�N�Y�	� {��I�ɍL�ݫ�G�R�k��Q�!E	�5E��.��:�͂2��y�m�-�.E��i�����YS�
��@�H�ۼ��nD��Y�l"BU�.TԊ�=�-�����q���Ǹ��j��ԋ����tr�a�ٵ�]�b	��%�ɔe�)rYOjX5;V��R�������M\�	D��ҏ����9c=�Vͼu��Ro�P�Jf�tRvsY��c�"n�XO��	3g���Q���^�Bʹ�7gQ+Г���$�-��t�8�����A���<����l-��*�|d�!�&�J1l��+�Xg�dي�5W:�{0�b�c���ж��fs�=G0@��N-�XJF���DC��O�<�j�H��r�?����˵������kF�̤H��6�' Lx� 	i�>񿘱k�d鷰Թꕜ�*�~���lW�w�'m�Y���O�|M��tb���i)K��PT%S"ԑ��&����q$g9=�U��(X�6���-6����6#�ʕ5B�|��<W"J2Kk�_7�_��l�����5S�oe˸��}�wvT�;J���jD1:*�X(��*�5���|�=��s*�8�~�����Z/��Q�=���HNS畿V2����5�ovrR��#�«˚��n�
�J�+���n�����_�e`���Y�	���PS�9�WA��M�w�����JL�+	���v���0�5*g�[8t�q�iH�$Dm+f�lrNt[o�oHŽ`�]�o��Fl�"��L���P�S$K�}0Q�R�>J�(
�7�}�}��M���F	1$ϛ,�]��2&��b�v/���s̀��ѧ��ʿ�^xI����s�^��0��3�p�YJ��9��<�& �~*=\bQ�5��xS�7q����Է�X�O06t�����O�R44>��|R���(Gw�ٿ�A"��0�MN����Z��������f�����O>�{��Wh-B�.�7;!Q88-�[�H�i�`��4�?�Ո�2�)b�hO%if`����#�D��� �M%�>Ѱ��.ߣFc÷L5	MB����G���T�}�%�[�^���Ƕ��	�0��O��+���-�E��� 8�U�a�q��K�&���9�;-0U�.�.�a�P?'��T*K����m�|����bP��ᲈ��'��vT�5�������q�d��۶a������Q������!���D��v�]��%�"�����f<Q���#cRNMH҂{)+��:�Q���R��9��y�ĩX���,�d��V��#��aw04�sH�#¥�̙�>v7q$�W6���p�6���\ɣ�j�����"Ūⰰ�\�֓,���_�9}�8��'(i�����5+�"�P�+6��B=��P���i�E�?���!#4\�"��<d�\��p�F�޳ojJ�Hx�#p5�����K��$1w&k��$�C����¼삵��.�a����K�����ZD�9�2%�S��T�v���6~�RU�R\3,GZi�븉6	��U%Q�~�Z�!���{�6Ga�>��eT�>����گ5����R�?�x
~�~yVű0A~�Y*Q�c�9�ZZ��c��J~ԄB}I�J��Nݚ�;�����ک�
�%��M�s�NI�(���L~;"�et�~�k(�|�<��>G�R��L�`j�ʽ������#��
����.�v#C����Iڏ���R�a� 2�;v.]���,AP��R=1\����T �`y ��W��G�1�C2��1�p�pF��'�N4����E�񀒻�LƟ%����L�wt�{%M� �	L���2?�k�$�NR2e̡B�n��xY�&4���֜��z��z�a#ݼ�r��w��F�7`�Θ(FS;e"�T�F}��a0�'���?r�x�I�I��&���[��?���'Y��f<�6��٫���0Yi���:{�E�Qw¾���Lh6�_)�l�N+���)NMf�`eB*ODn(���!ꄥ�|�w'q+��K�|��8��:�(�p���ܿ����[�H	v�풢ر֪iu��W�Nx�h���vp�3����g��ֳ`�������WI�g%�gVO�E��-A�[��Vl��4t`f��ƷV�n���W���W8a7Q�6�L��|�T
�Ryۓ��еYߧv_�i�!�	U��T8�O�/#uWo���;�s����)�ڸ����l{��4���'��~�X�hƁ��`(�}0��H�L6Ќ1nG= S�����>R�rS��}�:u�z;�>�z��:m��)/x�O �:�-����ޏ)��C��Bߙ0�LvH��cg'ew8�*I�Ry� 5���]�� [�'��%V�lڷ�
bcǛ�_�~ȳ+<�\p��( ���������P���Z4Yf��23�$dp�����΍2j)s5A�$o;���d�#�95�dTF���捱�n��<X�T�p���tPy�==���I��s(|[��sY�n�E����<��-�W��Pte�/�y�̚>�z�|���`������:gmQ��	���	He���S%bvKc�`
�_^�F���m�c����� ����d@��k��cs�ʄc��ڡ�o�A�?����N��0J�K�QPr�g�;�B@\��Uvy^bD*�&��n�E��_ܙ�qPl=ܞő��7_.ټ����guL;��zu�
�rZ�V�_(��7�b��Z�Q4,�6���?���b�e�L|��^=`_��p�e�g}�Ĳ;ţ0���/?���N(�W�ev�^��ME뾖�Z��6 A�e!r�U=��뭒���rB���d揆������yw6Xx�M=���n�M��ƺ�JW�HK�t�T�0[R��x(gݜ��\"�+R���͈�|��}V��睻��B��'�����{�S2o�����2�d�=;�F+.��^�7K����򘏙M:� �ٙ�ޙ���>�+���`�2i���g��l�����4�i}4#�a]I���p�1L�v�s�ϻ���,�[��R���k���.JC7LF�V������Q��L�1��FZ�Nme���K�`�'�]
}}���%X���Y��Cc,��*iG/��F߀��.��w�^�H��ľ���`i8���8��3��kbA��r���_�G7��@!蠦T6`���N���lp��}������`��/j3�!�c�HmT"�W�.�3���=>�����0���fU,ɠ��l��|�^����`�dy]��z��z\J^nJ[R�����K]8p$�X5��.&��%��ꚢ)}o�L��$�	�f�s��:Y�*F,���T����l�z�]�����t�����4��L>g!ݙ_��ag\j�:�s����ð%�ѩ9GL,xq�O�ٱ9�H��W6_HAg����z������Gl���(���V�Z:�xj�-�ҁQ�L��D�l'�C���?�߆?����ƀ��y���?Mg��r��`���l2���,(�){��KCL5 dS��HQ(IL�{�ݨ�*M�C����<�;����Tz�y ~�>���}� M��n,5ߙ�x
��#�'G8�E�'FY��l�Xθ�eiҀ�n:�[d���{���F����QRy/�F���1����[!k�kU�Y�{�|b��Lp2f������G=5�3��n���پ�����n�̈Z�pV�/e~�3m��:����nH�\� U�; ����ـ��*��������#�E�UT���@x���~y):-����P�����^�i-�P w�z�)�˗r�{���/����w< W�B!���9�t�*ڄQ|���`�N�f�ɬ��rq'y@�gj�W�\q�Ú�Ѿ^%k2����L�n�xyFV��]�2�+�d�e�m*��4z���x�p A�8��𠥵��dd�h�ur�������I�.�[�{�psn#s8{'��>T�^�P�A`��Z-�����^㞷���/1�0��rdԄ�0,��C�����Nk����6�(�D"ձ�CQ<���L�h���d���� 5�!�"��3��l��{M���c���&� ۛ6>� ��"X�fo�e����a�U�""p\+�2��D��S�N�*��ȑ<�=P#��~��5T�h�+�3ZY���OU�l�h]YvN��>��3�h�#�7��!�����֡�sv�m��i�����Ǌ*{xy���`��� 8tq5M�;�cOSE(!�	�A�DL��M[��15�ٳ�@%��ӟz\����l��!ޟ@m��,I-kF�.;7P� �ڇ_m�JG���\Y5���}
��,�G��|�/6���<�y.؏ԏzOɢ�L�+EֆrA��8��D1��4Փx�E(����M�ϧ��26awZ�b��'6~C��2 ��b&b⼆*�ߎ��+-@j	N�*@_	KJ����]w.�̎��M|�-ۀ:~�R�3[xk�Bq��5>�JjZn�f	YvC����gx���4�f�X���Zb?���^0�^,�Vϵ�b)2���̈́E���^T�r�1e���v8�����1�a#Ұ��Y�A�\&�0�::H���־�w[hjAVb�W�C� �.��k�����}�m��{e�=��/�Jn��\*A��[7����IP>?�<� ��f%di��-/�g.J�~�����y|ɇ��v=�����ٕ�-:,��{j���d�Qt*�L��S�q=�:ʪϠk!�hwrYjx<�{�n ���f�N�D���`���f9B���"�N]��E0ծ��[�ByS�*iI�R�q&%|ץ�ۘ�����ӊ�kLah����d�)�I��ٲ�0�+x(������9����RgY/!��.�~[b4ޡ%~;�pKXO_�O
32zM�'�v�y�@\�cN�(�/b3�>H)sT�6���佗��&��*��ta���ʘ�*�|:{6��U��~�'��[���� �z�5��G�9��"A��9�Y���찱����P1���Eq���������i��	�|�&
D�}��h3?�4*%�JF)\얄l�[�Q�7ɯJ��&Z7�0� ����3!`c�~�[��r�π֎�y)Y��?'�w��bN�Xô��������{T~��>o�?�ۚ*X��H��:d��@ể���a���Á%���҉��*���CRヺ�663�>s-�w����<
�%F��]D>�?}�}�OU�[6��P���CH�;����5�j�N�5��P�lJ'Q=|ʲd]��`�E<?o�y(����V��qm��9u+��Ed��������:k�ϖ�Ԁ�ǽ��Z0� �HFoN2��)�%T$���\v��.Č��e_��*XMA�S�^sOW��r�:m�6�o��A�Q_�Y:���GV�m��5=��M�%6�k���E�h_K�
."��è�&��/	%CW!@!��]?>�����4@�%�̔�Qj.v^�Yĉ��$mhRBYhnP�cđ�b�#�N/z݇�#���zM
5�2�	��{������}��
x���K����Tp��Q���v����M��J���-�x2����5��d{`�.�=���Ӟ�N�G��4��!t�	h���@WZ��Bx#��Bu.W̌��>�5	�ʆ���F &g8��H����a�*�2TΑ������=��l�FC�젩��P����h�M��1�������u�G*%�}k�|��8�t�56W�np��?4����9�$V.�U{^�(�s��X��-iQ���
D�q*f��L�g�� ���6�)O�rҶ�����-�l�kw���Y��-����&C(^�݁��:���֐�&6	?�ޢ���_԰��GWAAiR6��L���[�_��&C,����#a�!f��x��$8=*32�C���p f�wf��	U"M���"�#B�K�B;���z2ぷ�V‴�g�#i�igה�)�7���|n�w�O�R�$����k��-&4�����r���W�Y�qb��gV[�9��y12��$.������^߁�Xru/�W 2�Z���w6=�/s�E.ޡ#�hU��7*@_x�L� ܋�k��i��k6o�Fƈ�L_G(�lx�V�?j׬Á�^�|�~��\>(������Pܑ��B[��鮭��+�]��x�>'�l�:x��[�cM��4k'`�7Oc�2�&��2��`���.����w��p��ψ!��b�Sڎc}'O@c��n��=z�J��c�|��.|�E�~&̌r��Kv�dAw熁�#zZxexDv����ka������'ӯ2����]�,��bw�t�c�oV)���G���6+�oo=�ɦy��I���Mb�F�(����	¸�'�kZ{�!��0"�B�/J�&+!����ų�q�C`ӇY��(�o7@ڣ�*"'�
�4}�*����B�����ğ�m�N��*n��R��6HL� �)_W�\���;ͮC��w�-T�G%�(���M�2��|�'��l�8^Jʤ�+����Uj� EI_���ff�a� ��Q,����,ɺG�۫(����������L�D���du���5lw�����-/ ���r4�CJ �5'�?���7���>r�q�od�=�w%��(dutYpJs�n��	�oW��v�� �-�&ɻM�9�	�3��~����~�h�h�[�9���iP5^�{X�V-�b�~���R��Ƒݏ�,��m�٧�R���4D�?Cw���$2!��7�J�
ƚ�`���	�3{��ؽ��YI�l6A=x�k��7��x+�����J����ޭJVQ�J������Ē$�T��w���?E]4�+�#k��k�?{�:&�L
QSĴ�
p� ���&Zfue�#��R��CI�؁�L��=ێ�f�B�&���Lc˯<`��F��5�A��W���	`)� S���guf��p���j���q��Z��jo�&�;fkm�j	�j�)wM�C[Ӕ�E	��W���ۼ����<�J�:�m���"�0d�D<���p�s���&�Ѻ�eZ����`�?�����uqj��yj!f"$.:b.�yIa-j�$�5⒧b0*L��蠛���k��gv�W[[�(�W�����#֧�q�6?x1c��{J�1c���E�������a�E+aK�w����? M�d��Cx"r����ϕ!�]v�o��u5��Yq����c\�e� ���?�w�c��%����lRZ�V�Xy���V#D�J)=3ʾo�:�����0��و�e�B�ų�`��J���)]���I�@�����H���&8����;�'�ϻ�.!������!�˺�M���-�&��(GfE:ݎW.o��j��O H�bF�{�+��,m.��kY�p�������u�.���R����E��c��O@�tlV�'��W�<�~m����@�N�(ފ����a��uJ�������M^s7L��xR��'#y2�b�~�\B��U���� �;��-sP#Dj�)HKo��d��{������ֳ�SRY-J�mhHj���΁[=��S�`�����G��H>��J%���������?�D�ی�)(�s�2��_ld�q��u5eN��9C�Z[��O�}P:
�(2�d�5�|����k�ƬNlk< �n�%��\�>$ ���a�5�![:t&c��f�4 ,!@�Mi�i��+���c+4�#ړ��;�&�)]�=����[N���H����r���A�%2�@,vcS��՛w�窌ӓTK5��j^�u�Ci���̍WK"ߕ�L����E�n�1��a[�7O'o
V2"M����GSE�䄝���C�r����+!LC1T��^Y+?L?6޹�}�]S-�hx��闃����O�����t�h�?b*����1�
9Ȕ�v�m��������U0��˱�!?�l`�\bi����&X��Ol`s#�I�PJ��"�'�3L�:��%Yq��\��ysZ�o�Y�Ej?Ė�6��x�M՝"m���SD����E�X��[e��m��1�N{� Θ�3?F���	UN.P&Ĩ�E?�~?��s�����Ux��?�N�ێ{,_x�zإ52HuT0O��Q�0OU&D�j��}��0\ű��:y���e3@+=�ޗ딀�ccI��Fu�/o�>N�wv�i��mc҃:X�?���ߺ��_ˊ9�Z\�a*=*po{��Z\6��b޳��S(��F{8r�zg���(�1\C�t`S���3����^Xc�������l�,�y4(#�G=��0we�]��*�s�� �LTa��������q0�.��^\&�o���i�0����p���1��
��9=�����b�R�SM]5[��yހ&s�N�R��8�*���y͕�!�)�LYw*d��`�=�xD��X�C���d����Mk{����ـ�P� ��d�����w�lD�YotC��E���
�!�B�4cc�����`��T���4}.�� F�6�X�<x>�	��bB�����ng�N��\@J���!��{��+��Np��0X7
7��_�hU ������4�E:��-خ8t�1I�"�
���~ُ�Z��c�h��,�П뉺��=�S�����H��i*Z�矆y����m��e�z��;8#ɣ��#L����ͲN�M��H�%���sZ�W�����纈����QM0c�F�-Tآ/�����s"FӬ6e�-,T��G巜Z;�����D�]W�шc�eu�;�����"�5���R��q�e,l����@s��ȓ_�$NpK	�m�i��u`Y�\���4�8s�ڋ���#� �=�a�pD�w"��_�ض0BOq) ��`cW�P��ʴ�;J{��3/��-ɸ����Bq�x�(��	��A��`@�yaĸ����M����L�+����a'�On� ��+'	"�u[4/~fz��E%T�Ĝ|�I���wm�V�:G0;��`фj4�Gv20����]�Z*裝�1�,k�(������v*D����A�o�7�����ƷA�Og��rNmN�E1��_r��r|J��M����$���mӳ�T�9��P(�ec�s��,
UΉ������y��mrһB(����\�o�����)8\}�K��J�ySt�%�:�JT�a7�ŗe.Qz�<��p{�V�@�����1�)�is�E��OO�'�Ǻ�C��$Ro���xB�A(��16a�\������ ���"r�CG*E4
�3�#�#�c1����N�E�K��j�ЋLg�c�W����S�5�*�d��OI�A�S����}�J��!�=ԛ�2�$%F`�>ӡ(JQbRw��
�Ț
+YpE��pq�)sb��{�>.����F����e�ͭ��mbbk��ϛ��B�~f�ӛ�r��ϟG��!�B���0BH~ů�3�]VG����l���+�I4�?=�G��1�6$���#�WiE�z�RZNg���v��� ��ۙ�\��Ym��#��r�]˒53fΚ�ֳR�5S==�봵/g��8�y�%n����:���Y0�'f�[��2�����{� �1�x�zj����UIr�!��%���l�K���K�Q[6e��pV�=Z�	B7"ٶ�ɻ;����g������]�A�n�����Tur@�`4wH%��]e�YaI�����.3�2(`E�݂�������0#��处�	�������H�#����	�h�y6��K�U�uԇ��#�j�H�o	�4�&e%�h��f��KE�D���RX��;������i~&��yX�Z*n0X�%���uV���9Qa
��@�[WȒ�,�L��5�)j�em�p\��ҟ~
砈�ʝy�39i�=E��*bm�����t_1=�K�k����CV�K�I��E�n䊠�=����lua�?�b� ɠN����z�Os��[��Y0xz�(�uO�qKF�$�MK��z��T�e�ub�,%i�EZ����$6�VA��l��=UzIs}�������RZĜ��'T��䚃LeR��<����J��=�)"�����a��:��?�) ��1֞�^]?�S*"�p���T2&!�b:��ƀz�g��ղ��ڕa6*�M�ѱ�L�-�o:��9]x�兒�m��y�c��靶lR�Hݝ�!U3���}5�����������Y��SQ��� g���E�f18��B�7����o��%��԰L�C`x�X|M�
��i��2Id%����/W㔍:-�F06@%a�i�@���௪���;a�/\{t��I���:�I�txYKV0ŎJ�'��Ѹ�g5��k��)@d�h�T6h؊��Gȃ<LoU�I��C��
�-��-�,a�-��b��{@>�Ӆ0�gb^"����V@Q������=7��*fCNJ_ �����I��O�ֵR��Y�k[/�~0!�B�Ap�N�Y��:{<q�D���2��hh�)�MƁ�5�_�� `�59鿏Yo&ظA�N��xm�;t'�Y�ʣ��=���xq�B���G�)j4�GUD�m��9~~LˋȰ0�oյ_�!wB��7��=w��)�u�1"OC�6��|D��bD�m����j�P�����=r6�O�>��x�}�yٜU�?�Pd�lC7��yA������b�:�6>�߫��1���m��n@hF}\����\�
Fjyeu��l*��Jtť�\�~K�^�dw��No��LEsu�H<�t���MC~p�?�o+�^���K����T����J��(�@��8z;�1�^��5�6w�e4�P��G=�}�*O�4h|��y�d��-�A��9����>�_�[N��$�p�ˉϙVT���i~&o��B���ב�/ ��/H��+��"Fno���{)�kY��Y��-	!���*El�}UL!��6M-88'<���v)��z��֢�N@�����	���Qw�N}q$��b?j�W5�EnD�����Pm�\�'�?X��H��Q�v0̧D��;$v�ޫ�s>�lA�[�j��	�Y�	bG5p��Q��ko���d�`�cuS��C�	u��uډ|e����b�µ����]��t�Ib�2E�*k����I�3���j��$������0�>o�m�+兛�Z�s���;n�!������vF^f��Nr^�;�n�R�y�cV����.�.H�������P�p9N�,�$�"�DL٤Ξ�m^"�iTW�~�VGG���؎%�\Qn1�����
 �/-�2�%߯q �O�«<�����{�o\?B���1ɣ㈞� )��8�kB�#�o�W&�6�ЅAg
�{���^�����d|�_�o�1�R��pP�f�E�~�K���;��֝�u�U�TUs� 6%�&��0��<�Ὰ�kQY�ڏ�<���k<����Ll�C�p}�%�?zT�e� H��ɳ7�,U��#�GA���hB�&�,�\�/��G2�a /Ec�n��쬣�#�����<nQ�b���!���6yF�����+�̣k�÷gOZ����S1�(ݼ�(7ޝc�oR�ev++I���{��(r��Us|�ޔr�92ǐ��l�R�������ت�XClOE��W��� ���m�����ɳe`}O/�..g�Z�8��?���q�l�?O	ְ#�$�ln�Z���2�&��E��Y���ףټ�Rs&�&���pI��'մ���|a� �i�
p�'��ً�4��X��J0���T1�E�dW����J��0�˩�=��PRJ�{�t�/��q�&�&M��)���e��-���7a�B��훞�Jj��$���g�m ��c���Ά��(~��Hޜ�f���3�ސg�'��1)���^$[�&����#gX���m��1��L�J�����^Ml��H�RŽO(��aU��^1
��
մ7b�ؐ�`Z})HLbm�:]��܎n�SA>Q��E���m����^HC%i���ِ��a<.��R�P���~��䵺�a�ќ\#n���l%����O&��<4����	r`�K�5�/��H����2s��`gr�(u6��}�Kc:�>n?�~+�Ϭ��2�UBTpj�O"�>������n���fC&��c��:N�wA+��䚏ڋT��U2R�Z(��>D�a��/ �2��ڂ3��这({dq"�Ǉ�U�pbD;�����RRTF��N�c`g�����%�������!�N���b�HJ�uN�VGK�Me�>�0h��x�@���C��uBv�S�5�����q��'�u\GҰ���2Ec=�Z�|j���犱Ě��)�h�%#��R�!�hK����ga�	/��u�WT�$+�p��q����`��D^c�Qb���~hӕy[���D�h���P~����GvQ���4�-���(Ӽ��;m'&�L�"��B#�Q%`v� ڤ�dI�Rg���e/�6Χ�}���6�+�:o�K�ª�iG���DL㫛�v�HYK�#���<na�6=� n�^�}mn,딃���\(b�����P�/:2�BG�[2<�&w�$U��&��G�BW^v���/���N��e��% x�(x�º�����X�<�ڂZV]gϜ�>-ftLo>�i���Q��R���V���_�������糔��'v\z�3�l	jW�Ӯ�W�����z�>P��=Շ&a#k]�=��\z�Wd6D8̭�)v!��,�=7H@�b�_m&!�NFѝe�(��;9Mn�����:��r�v���!�S� p���� drBǴ�_l'5:������t���Š�IS�M�°�]��f���% L��Z�_�'�⇩ؓ����!};=
�
/'r��6|E*�BA�4i���U<TZ��[�&H�>��B,djb4A�:~Y�Қ��S(��˾��I�;z�RoP����f��Y��#@�.W�l,=�,r2re�e�����m`���Z��PCC��:Y������^G�j�'�h�IKC!Fk��<�l����W��&[e��0�0��'�v"7ZO��-a�UM� �Ç%O��W��Դ�5�eio�l����Y/%���
T��8���Xɋ�jW��������������a'����S�,Y��}��"3����e�~Ѕ� $t�V��2��[�M�7!E�X���s۔Q�\�*���^��V60˷c~���_�p�����Nޫ��1 j�7,�����n�:�ݶ3���/?[��b�OY��N��ֹ�?��sǖ��T��II 6n =$�Q��XΪ��������ڀ��[�j'	B<�Q�';߻�gh����*CƁHq�/'%t� ��?�а7��r���!%F��{��5~�V�,��H�
��,�'�R�����k�4����I��6x'��Q��<"6��(j"� �K�2"~�=܅�����+P",9��(Y��s�	#`;r��L�E���f5ڌ:p�� Ǆ�t�e��M���d�D󞛦�'��r��Q�;�,���`�t�XX����bQJ!<6�f���N�:ϣ�׌����P��չL�q��mamn���I�h&�K ֌� *_gCX~���"-�d- �y�΍�1��cb-�́�k��M���+4���U%~'3�EhB���8c.'w�-M/��=����[�ೡ!��%\߻���&�'\�͔�f�e�����f�t>��Z"4��"j����S?N��)���7@�2��W�^<���7�6yc���������<�������'�,��l�E�1�Zل�k�ޭ��Y�s�Mof.fNl��3��ͧ�1�������Q�P��׊��R���$Wf����ɘY���R�O��pU��ׅ�ơٝ� �X�'Wb��`�8!�tB�����sI��,J�n�<n�R6����0�� mR�獤��U��y�����|��f�%�b���V�-h�Z#!C��0�ܖ�afd���o*���-�����U��Y�<JqM��LtCn`�;�w�!��C3W�X�:�a½&����O��167�ӎ�)�E~�|M�JT6G�Ϸ�<�����ʬ
'ߴ���&��&�`z(�0���/���>�f\m�$�Z?@���9u��ԧ�'Y>|	۽��.܏h�N��d^�f�Hi+�zL/�7�6"
�>��]�E�_�QT��:t7���r;R�P��m����0�i�����P�g�mG2P<��崱�:�i�A��A�ց�p�������R�ԁ@����٪� �)B��N7�d�G��i�儼;[Z6������rbFS��8���l.�>;�6�$4ؿf��^H�:�B���?C���H�O�U�TY��V���;��v 1PlY�pWz��TA�o�;AՀ����XY%��k�j�U@S�y$`]��Mr/��u�D����?5,�Ķ�&X[=u�^��μ��ҩ�����vt���$��n񜝫�@��Ř!u)�я(|/�t�12���{+�[��2������@���G:_�E��a""�YLͯ9~�1GW�CU0�A(�>�ҩ��Q?��U�ϓ
��Jb2*��Jg��K�A��Y{s\��7���1K;Io�X��gJ7�r�v�5颫3��S��Xx�<&���Ie(��I�3{襸�k���~�0"��q�����iJ�z׆�.ON�P ��FӃl�,�Qv�=�L�QJ���[S�}^�%Jz$�9���0�|/�B8O��h#?���I�o:f]�P�d�om*�Q�����Ź�����+����*F��s#�ڞ�%)������I9�#!C,f!���=�=H5>�J�)�q�Z4���q�K�*h����5����=x|I��@LTF�o�&4�y`�<����9���]���=iU�>n,>C�Lw��mm�{i0P�΍��B�9���\��Z�FD�˪�}���5'�O�E#�줈wLB&E��鑟ځ���h� �G%��kR���^t�y_)�.I�a��z�q[y+�g��R��U�q�5D��1��X8�:�j����WD�A4Ћ�e�{-3_\*����#O��,�CeL�wb���Rx�+��j,���A|�T�L���Z'�=V��r��Ȯ�qƿ���ܮf=���
�7�x#�ksN��Y*�<���{�������R� 4أ6"���-l��=VQ�%�ɪm9A�C��W���ުyn�>4Y���\3A�����r��9ږ�lH�Q�Q�c�TUw�<1��IQ���d*����ZWac�n��Q��2��-��c#���z�	* O��ɿ���4�&'_8���42��<�r�d����1�����b�V�m��-�S��1�����̞�M*X$̡Cίb.���!K���S�s��ь4���j�`��Ol'1@���vn����yI��y� �H(@v�t\�4�F����.�����?rEH4+�#�Eϸ��zoc�k����E�r�?/0Tt�:�]��$
ے��e5>*��A���Ia���5�Q�b��$L77����~�r��4����4�I?]|����n���	�i�},۔!#Gh��-R�ؙi�mg�?|�}�V<ٵ��%$�H\��� +��t����N���S>�l�@���o���f:}z.ܒ-�$��@�F��BA��F���(װ��ܖn� G���R���/;��|�3�hhu�L�^��/;� &[b���)YGf��-�ّ�h����������.9����0p^h2��/Ȥ�����4-�ox��ω�[)ȇ�� 1���X����b�?�k�q���R��&K/9������l������%J���~G����=�C������Ré%�����7�H�R`�S7��?�M~R���k�I�7bSc.�ة����/��걦Gn��MF�V�*�r��75kQ��+x��Bɋ�$��� ���T�X��M�b0R�;���ڈx��k�Z���2C���R��&�$2�E�=x�LS����k������'`��
��vF�n��J����J��\��Mv${eo�o�1r}y��!����9~Q2��B��H����m���,�ד�]Z�*9"�������N� iw�FF�>��6�g4.���?�}4x������7q�`|=f[$-n8����&��Zl�ѡ��&�]8�,=�z�ݲ����/�$f����f��Ё?r���Ƹ�QJa�Q.�𪝉7��x/{������������<u��B.����O��m��S�v~� ���/k���b�`ܲT,��4�j�p���A;�r��֦/��t���a|DI����!K�β��5K�k����f�	^sж[l�0���Hr%��T�Y�n��,� Ǳ���I��/G���T����v#�Qb@L�nS�ҦʑI��k���o6A�89�{P�q֗	�SȒSd���.���<�ʗ��$\�]G���ͣ��rN˂>Vs����ΘP쀻�D�/P/Z�V�Ӄ�������\l�'Nw39~��8激)�EH��oh�*������H�Q�����0L�ٓ��y>y��%9��g�E�u������D5dӠT3��U@�Tm0<�£s�H��v-�cb��5R��v�/׎5��T�lj �����`�70>+i�IA��� h���C��>I.(��MG��d"w�<�B���
�LGn/���r�G}s����(k�2!���-�C�bl�$d��.q���=&�y ��>P�5R��S5�[���-�)��0��@�d���'�?T�q5�����Y�f��ӏ���	X
S���c���k�@8Ϗq�v��.�]y�Mr]7OՁ_��*\]Z}0��O�[��H�#]�?��r�{���܅;O;O
���6MʔmO'WM���Ƶ����7���(p ����yQ^�_���p���ɔ"Yi����?0x�$���&ԙ1��v�;���@�����o��FZPU)ctɖ:��������fN.�v@]\ᨀ������-���6,'�@��b�5�Pb~��w��\1	�i�bh3w��h�u}7f���=VL�et2�X} L�qdJ��s�llɼ�Qu��7I<l������1�I��먃�2ï��j?P�bI�_U�ż���<6HŤX�q*)�<�@���j�h�!nT0�A�i ^2����~�P@>�)a��
Y �ץZ`ۺ�(rb$	]3w��mL�� !�oW@.I�T�ehf��J�:�'��4����Ϻ�8��IƉ�N8x�l��xF�(E�ۿ��y"{����8z66�N��$3 e_ڄEKo@�;S�w(	PZOJ��f�X��UV3M���"j�����R��p�u�Ko�N�c��,��&s�5�� �[]~����{7��;��}QR~"�I��!�j�}��!�$�Β�����IЪx���Bi�۩�8���oy�5����_��O�#u �����
d��Q��l�&�����3�����K�;%�S%�0��k���goY�G��7M���r�j�X��q$~�y��ܿy
6:��3�IY�B�6��4��|<s�b�P�yA�3�����R�4lO���~�I����$d��<쒺5x>�B��n���+�<Δ������UaD�<���cIaY�h��X�� �(Cf�۸�r�xr��$�&
�?}'�?Mѷp�,��[?�_FC?�* ��!���Κ��_��)l��Z�B��j�-UEK���+2���dH�0+J�Q|���z�����U1C^�u�,}�d��im�#�۵z�}΀��"�:!�]�p�D���V�ů���z \�:�|��v�]'��=Cq��3[�SK��.�� �8HN5c���{�>�4�8��} �)aS���>��F쪙��*>���v%��;.�|Q���o��4�j����ޒ��c?q���S4Al��p����j���ʁ*�6,����0C��� ��W-��h����R��}�1�pl��O�q�}���6{α�e��p�&�h�����g��y��b8/��t��./֒�v%�@���!����*�p�6���M��$���B1�����$4�Y��R�y���,����Ȕ�Ċ�<����۵�F�&8-K��F�O���kĤ��"�?W�N�gY0��o=��}	�����1���i��W�i��%�ت�k>2#�6���&�����Z�nBr��*�  ��:)r����� �&i:}Ծ{�[�W�EH<�[�q��[6���+�H<�{fA#����>�;A���R��d�|�go�N�I2ȅ2�����(���N�Yc� <-d]�B�a��G~�N#���4N;����c%5����T�UO�ԥf��J5�Ἃ��!"��Eb=n���${���Ւ��"4>���ā�X���?��E�?��5{RAY�ʜ0����\�a�=���t�&G+�/�.%��,�w�| ً�Oqf�yU9�����[�	\uN��/�2��y�LD��;*�8q8�#���#@������j��K�EÅظ�oE��2��?�_w�-�Y�-��P��,,[����!�;[��"�6�:?O)����4G����^��7�/;Z�����,������~kX=��=�TA��s;߰\�����|H
�7a�t���r ���a �}�ցDZ`ѺcV)�.��K̃����6��W4���K����gv�{����ï�<��N��x0D��{[΅��PR�g�����e��5�h�ۭ���5����a�Rs1C�ټd�D���|!��dP��v��9��>��r���zz}Y���"!=�4=�y<�h�¦T�9���):c>�C�~Iԫ�����������зA���D���z��Ƕ�gw���򕥣����|��<D��k!����,NM�֑�9����{J'GĮ%+}�Z{7����A|�����6Ȋ\sI��-8��iF)r'p\0��FM���gt'�@��W1�{��=��m,�_vUQ���&o���*��τ�C���ɪ��$���c�o-�����o��$��/|C�bD�Y2��7���%BB��yA��P-Ӆ�c��s�o�\�����Ua*��������;�S�>S!y���I�c���l�$TK��m6��wg~�Q�.��7����q>*Fl�c9��?K������0����T5�G����Smv���ۑ�."�*�LY� $"cpGa����u��L�V)0cf��,[��I���q(nk-��˱����_�C����v�]�=}tJ!##����r*�n(�ߟ��¤����ݎW间�Y���+Ɖ^I8��o�.Ek?��ąc�q�ȹ�J`�w U�g�s�
��\sv�
��y��zz����ۡ�B^��W7H#�k=P'�W�*m20t����