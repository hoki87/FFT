��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�#&��#�<����貖���\&�
9ڠ�D���J[�J�\bT��0�o�o�o$�t�3�A9 e��q��}�&����/	�{"'���
��C��E��;��ν6���{7��q���Q�JU�Oz���!���5���
d�@�1)l�})���Gi�y����X�>�%��P�\��\Ō5on��?�K������/f�8�{3��?�N�L��֎[��E���ݟ��Հ"��h� CAQL���AC�[�0��f�v3N��p���iEۚ�DQ�I{��ݬ�E~IG�}�8L���{�����g����p�"h��f
[�z�N��9'S���r�����׻<~����8C�h5س�����l��uf�~�����:�����qQ\��q�~Мwo�+|���4�_��auEN���;�V�_�̂�Kh�թ�6��S�1Ե)��a�}T0[(������Caŗ�U�\3�א�Rs�ߔ-�j&5=:��m|N*U���!.�jv�=�@�kR���ۄ��adUg��pR�|
HK΁�3j�߼W�6�������lL�g0Vs��L�����)O�	����)�,��CŢ�B[6 �3-��Wgs���wM�A����P��[nY/�]jK=�;=Z3�V9g$�Cٓ�\�P�bL�����I.��C�:V�i�P[��������c9~�s ���Ϩ�㴆���-��ɭWL�r��90U�6�f�|X���	-l�!���ZgS��]\{y�2� �[{�F��66�<�8v���#�[-���W�$��B�7���n
ї'��� �j����Wew`a�v8���u��{����u{�Nv�0����7��Ypy+��?�Y�J#%U<b��������S7y��n�d��k0[W+t�	���v(�A1��|]��w?������^�q�鐁{R���s��}�������P�\Y�c�P����l����#�,n��Dzh���1�w(�Uv�~�۵��oz|�`�lX��P^x��W�(_�P6�Nm���W>�+�F�K�pu�P`��\��v����6H��:�(��Ip�ls���C�T?�l���c���i�!��1�ͱv��5=�N��v��Z���C ��:�J�y ��ⓨ�>�
&�]ސ�*Qc.� �2�!�W'��W0�^K}�]�_և $�pG$��_�4�Q��B�V0���&��V]����2�c"�""
�.�FP��A�}����В%+dX'�B����6�λ���'���V�cu�zj��������K��[5V��6�C '��K��W11<��sE]���\�C��:P�aԕ�8]1�t�k���-�p��d��i��I�l:��Pe؄�H��������_���_L@:*�&��@�1wf��ukh�3$7CO�ʥ��h�AC�	r�h�D�Ƿ[���1��~�<��IF���Ic��B�Eps�g(Z�y�9_�=���	��1��e���[1��+�K�C��=�X���!7��KQR��\B5mW`�U�9	��k��ze��Ƣvu�j�+:?������a��їiar���	��n)re�(�߯Lԟ���u۽`ػo��;w-�A�w��!��oӏzi���K�w���a����j��Գ�������E��ȡ����3#4���2�CɶW{Z�\�h��@�?�ײ��0�c�a���K�W@<��h��J?4z��Z7*���t�SC�+K����j0�`���Ř�(�FQ��:M��ԋ����z�)2�R���*Uo*�5s�=.I'q��%����&Al�z6�"g�fۦ�[I�ʂqMz��O��қ��o¯��B�uT���Fmg
T����+[�j���=�;�-f��]3�10�\-s>ձ�ӓ���4�oT	j
M��_�ˌ��S8ҭ�ǨH�I٩@�����-Ύ:��4A���J���D�J� ��Y[o �_6�b.������JxX~�-[Ğ_��Ɔ�*BI&��T$3��Y<�b�� +,Þ]�	����؋���,[�߸ Rg���I٦�5  ��ŕ���V
3S��6�cȚ��c�<&S6=>��`�ϔ�3��dVx(�c��;s�,A��6K0�q��hS���G3�4ʽ�D�BT��o6�A*���0n'����l�M�h�FA���8�V���J���E=O ����о�j����W��O�I��1�oF=�T��G*�~,��}��&z� �()�{ˍ�RN&}�f�sV�"����p�I�s<�y:O���sY�����S���8ْ� m�$�M�+4��z��B�kr�b&?��ϴl�	fq �Qz��P�|�$Q��E�5LU��!����wOSl��@�-ou��rD�h���ow���[�"=�0?��?�CUŷ��Ԑ�J��d�`��<e:��rs�t��ǳ�-}��ؼv�
��>��F�b��s�|D�&D0�BB{s�>�"^��w�zCw�n�Z&�"t�AC�&�*��gY_=BZh<$y��~|>�cu�2�qV�E`y�e%֫_��&���#��S�f"7�y���H,�l����������@���縺���O����� ����đ�g�q�	���h \*�,����~Ҟ���F����^Xe,�2�Y��Zw��R��������;Yo�h�����%`�:4^��#�AԻ5ڐR�j|!5O�;HA�)Hԫ[^��ӛ��ZR"��/�%�v뉞L�:�޸�O�b��L��Զ?�5��� ��E��^~�i�a��*�B���6d�_A�3�R]�NbQH65�WBw~4��C�s�(C��J�3~�F�V���
�(�����Y�]菄�7Y���,;ժT'�ƺ\T����y�qv��Y�/�dϜqRo�g>�v��3�f���k@��@;��z��Ju{������)e$���=3��<��*ȸ��ؑ�F
�[+��ղ����h�N�D��y�JZ��W�L����"�C��v���`]�<VɁ)l7SS�K�����n��~=�i��b� ���,4�&���'#� _�[�x���v�B�g�*3�g�&0C_�	[�����f���A��̴����q����u���� 0��P��D�!��hg�@9�<c��զ[#�(,rJ�4|U_�\d>
X�`�Y�A����_��Mx���3��Z�����Ã�82�z'0�sK���7�/���C�d���S��gK�~�j�J q�n4}@�
��U"�(:�_\E�y��������à�
�\��i|3�X�	Ay�꾪��.|0)���-����ʶEo�W���P�]w�;���8T֗M��,��b��=֘9bJp���Y��� @���ܹ���M
�����1�̤�n�:�=�(�K������r�68��ءE�gT�O���8� #Pf���Cu8��ʣ��$D:� j4z-ԣSYC�9����y�i�<�/1�#��Ş��q�Ky�ں�^���d4u:�L�J~d�kK�F�'�Bx���'ȋ6��Ym}_��`S�������N���-������-@vwHe�/I\wˊQ���^���I���jƮZo�� �/�;�inK�m/���(���[e?���I=[�?�'�ɗ���Ux�-����C|��t >[��̨z}+!P<ؼy�Q;��k�,�&��=(��~`y(Znj�-�x~s�>V�DW��0�Y�(YQ�)�HP}���nc�\���}�3f��_�Ћ|��t/���K�WN�QG��j��!�};.��0o-�Q�����(_�����g�O
O��A¾С����P��v�&��5�y�+:����45t~��z��g]l>�O��� Ȇ�$0��^��j�X-�ӝ�ƞMP��ްE�r�
��P� �xVs��W�`����O��H�����l�Җ4���&y_j���x��O�3�H�/ROou�'��d��ϗ��$f�VQ�2�d�j�ݮ;�]��TH1��A�!i���K8咙��G�[ab�y�PBw�|��Y\���U�6�a�b�)��*�5�R�P��ł�Cm�R2\4m�MK�e��F���bk��#��2�!Pq��ǉy��nh�8�c10{��X=y��}?�-��m�38�]�׸�\����q(������t��+�k6}3��>�ei<�ZsScv��v�,&�B:�ԻA>��	���@%/�%G�Ry�Vg �P]��7+ǎ�!>��{c���h��E��W1�4D�L��z�m,g�}s��k��/�C$����#i֪�~�d���E��\�룬v�Z�����%�0�Is�)כ0��2��AiesV��AB�C�A�{u�ޣ���D�P �OYt;5�_^�a�<�_�C�Ε���tD���/�5���
%�P�g2a1��EO���������Qᤪ�j��}��S�n �����>�!��b�V�&�;w�P���*�6�#�ϣ�ͦ^	W��
�x�ҙ�G�9ZR8���	�Q7�%RC��恍]!�ES/[*1�C`��+j����>��Ömޮ`�Z�X���d�%��,��D/!GX��q).�Rk1��9�2ɥ�����$oJ	���X�ð�6�9}O�z6�Fo�P���I6V�P:?DLc�䳋5��K/w����+�b�Qn�*�mi��w�I[�r�Y^������"�HO4��D@���bG0z�O%�]l����ϦP��L��=m�B��aЇ���nM"��<���rS�8S�{�z������o�ˮ���fRdk�%stE�Tr-�aڱ�J�l��(��OqCi���ҽ�#nk�"o3�25���l�`������6��D���an�_�[�f���	Y��ip�<�f�:^F��
XD���F��a
ˑSR�N��e��ߨ�L9���XkU�����yl@�[q�M(]S,����&���9S���.ѪAQ]�F���s����])��h����o�ՃÓ�{���͜�u�޼�Ʋ�ZW\���%�ׇ�/�j�'��>��]�<�p�q��}y�_�O�<o�d�&����j��dS}V�Efxr����#��)gb�����X��5e�$�|��;C� �h����N��n���q��!�T�1S�.<'�@��3�L}�rM��C	ɮ�F�@-�,���`���<RF�ݸ�S�p����\BK ^�ՠ"(2�IQ`%r�(���qT�4iagm���6��M��-.9�8��c/Y�H'���X�7k�3��o�ݷ��2!����Q�kO�'�����O�U<�V2ؒ���8Sy�+_��Ng�yj�I�w]�����;�ћr[] }��/"���NX��
.ͮR	/��}խZ.h&'t_������WQ�t}��1��E�''��X0�}�$u>XEH��F0�s�귮�Ĵu��ro�۷Z��hC���#lwa#x�\{���̜3�fh��� �5�q�O_u�[���Q(7�cBAȊ���%\����q�@t=n;���r�I�g��(E���8Z��+��&�uH�X��0��p��"���Y�J�7�t�FE���q|��S�M~#��e��\���i�U�{z���qOC�9Is�=�rDza�1}j���W�4�V��E�J{����(��q=mk��~�::��;�V�-�w�fꯩ�?I�r�}���g��2�~�>Sw�#p�Z[���̎�-��H:�#����XC\G�3Xf%Ns3)���^�͍N�6�7�A�a5]<�	Q�èLG/h���k�$�G�꡺~Ѕi1uc��?�!��Ewe�W��;bLaTe���f�,�ʪ����u����Y��ƍF��N�wj�P�Ex���h�"]FH��y`/���`ft'+�ú`��	���L��Ŵ`�����*�b�#���Jl�洫])b���c����1xҥ̅/M�vl��w����}/�,|AJ�6��s��r�,>��m�������?�֖H!ٻ`�yglw/���X��3�S0�[s���gF�0�ǆ�n!r�km�7�ؚlŮ��ǛAiY(>�� �
6�LN`)������Z�`�:��i�o�Q�*�ٸ,4*�8�t�XԼ�K�w�qÜ�)��u�h�v�0K��ʹ��;�'A�̛,����oڀ�+q~�ĩ؝-y%}�fؕ��޶.��]�$�iFŞ��6��10��Ի��{U�<" Ҽ� ��q�E�c
[ʼ��� ��W��g�=il����81�7a�D��C�Eїd		7-����BlU m��r�ȰM�F�Ԛ���#a�$*�p���x>i�� F^4�'�َ�������Z����@f��A)��n��a��P����O/gGܻ�П���rwj�qC�9rA���_���Y���2��0���t!�/?K�#fFXų4�)�s�>�P�=�їJf�gp� I��i��ðC5� �$��R��)4����We��U�����J�zP���D���?W{�5H�TŦ-�ۮ҆��a���GP�����&�:�sM�-���.��J�0��kh��!+ъ��2<lNM}U}�b�c!:o9`K��ծ跗xi��	�!4ǋT�yL�O�f@��V�y��ضV���}�5�
h�W{ss�����T�6��ճg���)V̱��!��bK�^ ��+�j��d�ꄅ���&c'��S]�aJ����A\}���`��,�
 �� 9JAa����+v�ݱ�})ǲa�}R#Q���H�C�q��g��LL�fBFZ���7&�)�ȱs�W�]�mn��D&��jv#	.}�Q�&,
u��l$֌$�U��'7�e.G���EES�;�