��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#���������l��U�~�׏O����j9�PY���`T���x���s����uí������P��"��b%>�1eτy�<�gܰ�N�Y�	� {��I�ɍL�ݫ�G�R�k��Q�!E	�5E��.��:�͂2��y�m�-�.E��i�����YS�
��@�H�ۼ��nD��Y�l"BU�.TԊ�=�-�����q���Ǹ��j��ԋ����tr�a�ٵ�]�b	��%�ɔe�)rYOjX5;V��R�������M\�	D��ҏ����9c=�Vͼu��Ro�P�Jf�tRvsY��c�"n�XO��	3g���Q���^�Bʹ�7gQ+Г���$�-��t�8�����A���<����l-��*�|dgM.�{�F��]�|�b8�،��}5�AŞbs�/�~@����{�af�9
z�ߩ�P!43`P���Z��߼w�g���r��d k��a����
���ƻg5ۅ�N4�>�/+��˧�I��pP�v��Y̝�q.�/1Mñ�f��!B�{Z��@�SKe���]�W��&�?���|�E���p"a�9�j�!>���c&Ɖ���d�@�Za:��խ�2���/��겄!��51�Pe�F�Lk���9T��NP�V����c�ȇ]g��!�џmC�[��X�ߢ�O�2���ݽx�=LFn��	�9�u�͛�f�	�a4am����&T�T]�S�Wu[ĸyU5^ݕ�zF�7ч.^��,1w���|k���(_C�`���#0L[;��P����Dx�NX,�~g'K���@m�?��pϒ.�w����S0Aq>Cp5z�3�$�D)��9�si���{��p�~��k���d1`�v����ΎX�ǘ�DN�|���d΃8�)BjwueJ��_~m��k8��K'r��«�X}�t$�{=ϾZ�φ�u
^7KO;����5���R�l�df�5��ywV��m���g}BO����PƵ��i	qk��f�M&�q�0�����|���N�Xno�fb'�켅����
��'a����s&��I�H�W'
��3���-�-+�R��+���t��V�_�bkS�nwƄf�u0�9E"����k���C"���g�}.�v�gDK�q�f8�׋A��{�#-:A,�
� �'�R�R%��1,�d�+iW 1���m�І��Vm/2X<�q{0(�y
��q6	���l39�5x�MwB?䴧\�$���ӌ�[����$�q���6��얅�l�x���NQ�q��3/u'�ܒ}#�G a�����gK��#�����mI�r�~(���̆��P%w�ߗ������~��=���6�P�}���,	�_K� �墸���E��F�\�8�.
�oڱ����!��ێ<��b_���{m�eU�Ϗ_�.���Lf�H5\3	�ES@�t��ʰү%��`!���N=�����Y���t�����܍®t�GG��m膃eĽ�f�W8�X����y�����u��B�tؗpl�4��\��R�~L���v���F��p#��$���ʝ����Fd��W��"f]�ę��j18��8�ז�ﾭ�� IW�S!��BՕ]T�Es��
1��m�E�QP�Ջ`&������'��<�f>!ƺ6p�D�H�SG1�.�,����'�2E�>&� ���1|�fk.��t��GG<#+@"0�Wc��K�/�}��_!���r'�_����:
-�3���ٙ��:�6�M:�4�AF���.�}; o�Ƭ����0�w��7$�x�*�a���,g"j�V�~ʔ�~�o4�h0�L�}\;���
b�Z��J?�,$״by�V6��0������^��8C ���``�}�I���<F�XM�	y��:�˜;��5�ݯ		 ��iS���q�7��l��J��6)Gಡ�w&��%F���P��%�[킑�C���+��K�WP�j7ϵ�tl�
�7Y*����Ez�|��e[1%袢I���R���>r\��pSѩ]���]�3�w�Tk�a-��{Ҝ���J���%5[�����wn>؆%6���k���q��:��#B<k���ťg �a��eM"�4y`6�o��&"j���tl?P.lѮs�:)�K?(�����鎀�m+�e�#�O3��sP�w�A`15 ��G����)��z��F��c���/)��?є�3�F+W�V��yA�5�����	5bl%2IlW����8;��>bn�ѼL֗i�#^��%��X����s�~,��fD��ϐň�NM�5��3���1�E"T���"~$c�?j@ w�������.ݨ|�,�m�`4�k�{�3Ā��n��;���P`�ʧ�=��(�-�f�k�*�+!`��ϊH
M�����R]��s�j�8���4���i��p�]�^���3���KԸnH��́ϡH<v���@YYG�%��JiIv��Ï��ɾh�U�e4U�f��H'"8Aato��KUS��ј��1議�y�6�V"jY4�T�X$NIi�o ��-k��q��F�]v���-�z�MEe��U�a�Do���NFX�Û<�e%�B��Wջ%��VF�N��3V;ʗ����4��4d:KM�{��AV�c+' W���� @˗���L�~҄���>��(z`}J�T'���x,[����+����8�z`"`J�#p%�/��9
>M�jU~:�"�\����E#Y(s�?��8�P���LC>�(J�T�D��{y�|d��L�x)LZ�d `���liho�xZOj�?�㢮��^<!���*Ɂ�ѧ�E��3�پ���=���q�vr�!󱊜l�T�R�C���M��"ӹ%��2�[z�v�'|�q�����,���2����괴w�k0${ ���V�vH',�>��*<k��t�%V����[����, �5�d�{y�ﴓ5wx"�޲sYR\�I\U�b[�3��B���>)LQ�-q���퀠�j_i%/���"����4�W2.����QV�2���H��$��zז8C����ۋ��9뉚*d�S�@��6~��8����+z�4��lj������D���veK*a3l�ډ�nEK�l�mB\�����~
�軗:y��T��T��N뤈`D�L���r/����'Ĵ����/��]�O��O���#N�&�U��'�ч4Y?�'�"���Iea�7��3D�j2G��D���6�a�{�GNo|����Ӝ�sS�A `�tĦ~E�&�ga=vţ�1I���7w��c�%�'�U���S�r%)A+�B��Қ�e]�O��m�$ـ6�7W�u�^vs�m-'b[�c�I���J�;���,x��]�q���g�GBN�eq �ǲ�?k�L_�H@i���t�ٯ�>\ђ�7q�����G�唞z!�}֘9�D�m�jےք�?�P������b�0�9�r�����>rp��sr�݅��gFk�z����<ne��N#2��dq�%�fr<�0��W�H�<�J����B�B���. ����G�ģ8��Z��N,�.Ņ��	�<y����S�3��������6��1�t�� cb�;"(���j�C��{�f�S����^h/�����ݖ�k�XWQ���_
�E�Nڐ{bR�ykK�1&��8�� _��68=�H�h���J�f
e��w�j����~��S��0'���0"c�Y��E��cbQ�>�1�po81�����S��,&������o$Gu9[�4���1X����hnT�ܢI�!��}���q��x}���]�Z0J����F�x#{��\��EKua�������>ƅ9�[5���)@��ek@jtde�B/�����`�j0�kB~���V>��G�8ho7k������0��FBj]��	�X`\���*�q������پ4�b9qC�j֋�I�Z�D�9I�ѭIh��9W�{d�GҨ� X�'��?�-�7.�0K�W�R��3�|	����F�t/%�t�9�/�،@f�"��-�4��|_1��k�,|2Ah�.=�)q�t-�+���Gn#\�ܛ�\7��"�&d���nD�d�4��վ�-�Q`����\n0���|r8�b��ZH���[S*�GTgh`�Q�8�� �Z׺	Ӊ���}�_5m�}E�)����J#HlE��ޤ9 �{��2t4u��W��4$����v:�����PdX�8I���\��������7D�}�>A;�a�������m�7�T�� ���v�U>b ����=y`z+�4
�py��7fu�?=�h{�B�:RJ�߶�4���/r�(^	�Ma��m��ˉY����AY�����HZ!�X��MK�&+�;L��ÖN)��,�~ȶJ�U���-]/�?
13�Ҵa_Sz�c��o
��&!�4�s��iÖ/�!"��'��#����62pF-��r>��WDo.po����̔#�v��C8��O��/B�X���q��pj�J=�-��2M�`YvYPRo��`�>�L,{����X��K����f�e��h�`2�)D��	H5�~��p���U5��a�M	鎘��9�*��@�S��;��%>��A#��|S�ו�*�y�y��}|4��b[�I�����#9��U���> ����I�����Kh�r�	��S���m�r{�7�.,�F:�V}9"����1qɔ2�}�;�t���p��iHa�3!B�;p���Z�a�f؇��
�2u-4K*���x�C�5R3)��*�����S�`	���9����<��{�A�C����A�*V)d(�}Y�-H��C�Ñ���V���sX����gOXBp�m��w[";�^V$����y�E8?��n�R��Ńo1G�]q�p-t	��&N:LK.m��u%��]�0����Wjl���T���5E�S�Γ�o���Hw<'�I�����^�����J&F�/gN�]ÞE��{`�Z���	E���61t��>��(����_L��C5��F������au�T�r�[Ht�}�h�W���dE#�#A�4sr ���iM�Q|���Sh� ���q�~�
ޒ̫����g�fr!-rS�2<�nmW�徐�J�!�D��O9�!��,5��z��:�p�8��}5���a/��m�lO#XF
t�~^ؔ��N��B��
D�v:�DQ��=j?pȀ�����>f����I��g*��T��]��y�}g'�o}���z�N���,�埧b��ܑ:2��\��C~Me���k�p�"����HB���7u���Ǥ�<���Eo�L����8t 3��8N�:<f�:V�`y"q�è��<+Nl�jf��Ƌ��S�x���X3��4_?O���i:s�-	Z��93e�*B�v�0�"�	�lu�\l8��L�7���!y�]��Cr�ݎ;i{�q�&"��ԝ7��R����HO�����.$ye�:7��$�"�j���sQTs=�wن�����B�AD��F�Tk�|��b?�Ճ�>�H��2B��ޛ]�����>��s�Y�>��_�����VS-�]�gE���ԭ��P.�0oUnB(C5C�����������k�C��瀠�h>%µ�g����X�(�ssG�,��F�A||H:��P�|�[���+��}@/6~�N7��b�HJC�n���Wr��i�R��Z�]S��(CQ�Z)��N��u�~�	��uIU#�7����k(��F'2��<T�pr?�!=MM?j8��˫$��C��v$Ώ�>�Xy2�Rh���y�U���X��-j��	�Hp G�%Hjrh��L����<�7 #�|v��O{k�]�5�&�:����Vs[�W;���g��R6�;x>]�M�x���E���w�A軯�~�c�}�_Lys
хFB�G����!��M�]1�j�$�b����'SY��x�RZ<��+�ۼ��{qCF9��>3�4a�Z�>NY�ou����vZL�H���P�[�8LJ�I�"�����ZC�YM�l��5ׇ�j�r�4���%�����8�XԱ�f-q�
jj�N��+z��o��d�5�4cwY�X�&��c���E#g�6b����P�N��, 
nY��#]4�<�����-UJ�+�.�k��:�2 �Rx�w�dCJJv�Z���=.�;���h�&_�'����upX��o���.��W_�oR���8/���9l_�6��m���`���[D3�ۯ��X����8;�qv�ڎ�]B(�څ/���l�����ZW�K�:��`��0�ڃ�\b�]�uK��X�h ��������_]���մ��h�y�!%A���es��Mد�p��������ؽ*騫W���c��VE>�
z���$��T����?^��5�@�lG8&U+����9:h���1ў$ s�ґ3KΝ��� ,�d&x!�y�ke�S����L͜$�x�;IDI/�<�]YW?t�~��X`h�z��yc3N��s�W���t3����KR��{�&��[a��z+�L+���*���T<�d�;+��X��4<w`~�u�x\��A��+e��UD��U��]�]��hl/`9��|}��|�<������+̊��ξ"jlM[�7�ڂIDf���<���\�J����Z�j��Ղ�yUτ���\1>*����F܎��v4���u��e���+9��-��B%�n�`����||�W6������H׊b����#Z_7��oA�3��>��	��=�g����"ǁ�_p��l��)ų�2���3U����\�7�l�IQQt^�	���"�R���vH�C
�k���G��HUJp�AS
	{b�߇�p6.�5��0��{v+hM���.�*��BU�ȟXmZ>ʄ�kЏ���
�nϛ�撹ym���[�,:(>q�E7e")����-T�~C��`-zܧ�� |�6P�8o7�������p*k��d�2��Ǖ:XؖIW��Ö�&�� �Cc�`T�X��U�����i	��~@ܒ-Z�~�sVv��l
�Q�p�]�JW]�ކ�5Gt�8��H���	����S�/�p���uf�~vs����AOx=r{��R�xӵ,��h�W�p-�b:�A ��7'*�����̳̕h"�_�N�Y��F5��L�Wc)ӄ��<��%$*����厏��s�G�4� �Ʀ�i�X�[�E��%	6>(4���������E�e��_���HhG�1M�G�_�9 Ry� �>�*z���|���J�ZO�tF�*�UC�> ���	�]E�"��A�#�d]�h�e�a
���5&�K�5�p@f�,E��/k�^֭�
��'E2ff�WV�sF�.���9`��%��"w�p�|oj���Q-���=N�yǕtIQ�ދ����2���#,L������ؕ��.�G�)J��_Gk��n���5UPS�M}�Ms;��}%���}��0�O�(��u�˔Aڕ���)mf_W�"}�+�r	Q�T�6�+��>�5倨  QN��]����$@�VE����W����y� �)���a�"�Ǜ�)�u)Ұ�e�|!�����ו,.N_s�Z�)��ǏpW�ˬ  ���6�f�Ūm�s���������j��_�b�;�p�h��]B�U����S8��+���y,X���N)��C,��*}Lm��aB֙l���
$� ��Җ�v�\����2r�/b9���}$���v�B2x�>�� ��F���	<qo�H�>=s,����ݜ����I_�;f���V'��1�I{�l����m�t�,P��h���X�2�{)�Z8��)4�Ǌ�O�� Nqt�=(8L����C��O��t��K��fF���⤟_~{��8��E�F=��)��_�H�����v���j�ۛH�ീf�N�bzt|�p0���o��	�clю��c��W|�[��z�߭�;_&J�E��|~"L(Tv?{}��{�8�ّ�����5���߃`6�3i�N�d�ŬB���8|V�(�kwgc��,,@���1`�EYZ��:
N�]���+�C��QzI������PI�A���J�����r.i/;RJ.',�i94Q����/���F�f���$v�����:]��;Où&�7���~�#�՜��Y7�2�����^'��6�6g�2�(Na.OR��nd�R������]Q�n(70�ew����y�x� f%j���HE��<FT�����?R�3(����C�aK��Zf1O�����n��f��~��̹�!��@��+��15�gkq[��v������q�B����4�����q��/�QF����Yv.o���Q�kޑ	ə�D�j�i�$���n�\Ob|U0���[~̱Z��N,� 5�\�KҮt�G�t�bCy�**�Hu�g�(����8]��醳�����g4O�?�������B/��@���@��:�t������y��C��_��p�)%`X�3��A0?ߔ�2t��.#�³I�4��_��u�n:lk��^����Ðᏺ/Ic{* {U'�?�j�����5�	�Q�F�KJ6�k����{�R�?��ږ�
����Y�:��癐Ò`5�˥b,ԱAtr�c�t�U1������/���b�ؠ��0jT&����+��*;����L0���0g�>;�8m������p�B~�o����h� -)dK؛��rt�-jYKf�u�$�1���I�N�K�sw�
�Q
�����,�^�����j��ʏ�0 DAXі��V��I��>^���0~��� ��2�w@�f�k�ٔb1T���=R��8�#�D��6�����J	�MS���Q���0X��=�
lαq��s7B���~h�I����TQ��~˒�#K;q1���=��GWN�?6�.��d"�B�>D��Ox��_W�𤷼N�0ek��F�Xc˕~
�
�%��%h�����TQ�p>8�s�ȭ%�o�u��4N�]_S�m!�f���Â
������w���i�$/��^�`�)`H!~ӧw����n)�4�%&Қ�iy��m�eJ)���7�g�N�\�����@�+���j��cy��Y�ӏ<����͕H�wi��O\��q�x�I�U[:��M�Ҍ��G�IB6D/)�u��"��}������)F��#�B1�����#�Z�4և�B7�A����6)��]��Ċ��c��U`^�7��u�RX��'G7���1�����0�R��T�� mNW��02��ERP~�|�R�Ԛ�(b�)t����3D�f,���ǈ�
�l1��0�k����8.ӻU���S�m�WN��!�KVdj��ӟ�N?��6�xFM��J�R&�`NT�+�,���JX�vF@ee8V�>1�O`y�fqG���~����QA>P o��;7hr+}�kL�	ܪ7GY�	�6�3�ۂ��������Э�y��Z��l�Ʃ�|m������e;�TGþ��)�z﴾�Ҡ`6|�P�z�,&,�t}#;z&BjH�V�T�5Tnu�É�t��p��Y5UAM�e�n ��ä�)m	�bs�K#4A�ŷX��=t���I.�SY%�+-l�n< v��g)�{/#x��
ߏ]v��c��[����bΆ�u!��!���0���� �(,
}��KN��U������?��e%��gv��8�<�9�!��9T|����@e�5�a�勜�vŎ-�S��9dAm��6�׈��T�r�[�h��IB[��}��!<�O�`�Y��L����5��Nj'�H��+����ù��y��Rd�r�>�P�$��7`�gpkٺZJ9
M�ߧԉ|��㎕T���[�O`��� i4G������?������1����T�Я��Hm�@�	��7RDg��,#��tOj�J�Td�Pm��zJ(�q�;{��Z�ڢ�k,���uD��p�4h�iI¶�K�+�P5A��}ܡ:�w4��X��p�d�d�a�Sv�=Ռ����&m�o�OL�ġx8��?�َ���1�ѼaM��6[1��S�h���x��ڇ̊�l��ݮ��Kv&^��';E��3[i&�&�}9�@���*��HVQ���U#ڶ���Ә�HG��`�f N��Uh��n��&�d�G�&��d�U\��/���q����j�ܭM*%��援J"�E*��j��:������PCOL��R�*���{݊ň���+�B<,J%��@D�;ry�A:���$,���z�De|��cH��H($
ƙ�S���=���1��U ���5��
n�����u60��B�d|`$���K���UP��]EƄ��. �~f�N[�a~���Mq�®��.B���㇍������ʢdP�
��6�;b��tt��Yh��C�^@���#PxM�F�܊�����@u�O�Sᕟ��x`���T;���եξ=_'�#��`5���D�L1]B�%��fO��|���/C�-*�b�"����)�1;��	���:��0)��Q��iM�pT#F@�<r��y�����~6E����ZiDa�U[(;����d!z+U���1$��V�ئ`Y�s��Gq�F�~�t��-Qa��^�:����NcZA��N�\�}>�ð6`h{�JN�:�3lBG�ю�7�&��y]*��Gg���K�<^[ Id|�y����vaK��琀[A���>���+�N?���f-^>��Np?��?Y�	�b�_	��$�e�E����ze��QW�&A9᦮JX%"��Ϯ$���3��)4��D�-q�����fҫ����Ɂ�Y���\��2�H��I�g�h��&T7��u��,�B���}���� ����(��yB��&��,*�j�����ѻ�tI@�=u���X���0qR�=�R���iI~��J�ٿh�,�q�k��j"간J�M�|���Xpp�� 6�������U�Pݢ��U�x�O��xz^��y�*,��l��Vx�O��cJ�v�?��PZ��8n���S��E9��\#��7��TZ5ڏ�Ly�x�/(̩}F��Ӌ˿kء�u����i4���x5˕�B$�;=�Ksl�qE�ڊ7{Dȏ���@� ��<�g3V����~Ƙ����.���86 2�������5���[����X-��I� p���I������v��5u�y�$�����:�_����D"��n�����j 6���\��bP0���:�nÿ�[}�--�@jk��mec�,�� �Ȇb�H�u�t�>Y��e��f��S���@�*SC�!Y��;Q�2�B��>F���x�#�Z�62LnN0���'/R�L�11�!�ـ�Ny��?r�s .X:> H��)�Y�[T��#P?�����B޺�	�Mq�]`<FVK�覠�fܩZ?����W����	�7�@`>��y1@#�Y�z��Asa��t���3u�5��nDh���p�����m~�x�Va�6������a&�C����?�9{B0p�ץ��믶�W>��j��!9�zf��ע{[Ӊ�f��]C�ν9�.��鶗$3d�rIls�Q0ԃ��5�&���������ej��QGd��uQ<�Iv*�٘����?(����!������o��3��Nᑊ"�u��n^i#"��E�mn�'RL>��
��~��U>�@�9��ttvrT�	Ѫ��6���uU���Ǻ�.�U�	�{�x�GU�]�����/�����$��n%���SB"��v���[���\My%���kX�<\͌ʷ�Л���~�y�w��f�=υ�1Byp���>�����oJS���GAV�ȒY%��Xps.��=��5���m�E���?YY5x��o'� D��I��Bs��O��z.�Ŭ�=]z�"L}0%:�< ����G$�t�����g/��I=YDD���o�������!XB��&��%\�M�j��S �n��O-�U�F�}~u�̵3��!'��LX1�y��Z�#�僗��������g��t@�������dj$����u�� ګ�#��7qc����^I�~Jht��U�ab���%����TPM���x"��Nf�ۅ$1�$O�ES|-�����.��u)��e9$>��Om�]q��H;�75f�������˜�b%�h%�C ү�];p���}Aj���[��1\ݔ������8��/!
����ԫ��fحlX�!�-��L��n�ňc�����:;Ȝ�F~�{���67d���� �qɷJ���y���b�U��}�h��@:�Ep�i���ŬgN�����V\:�A;��d�=^���K�\XqO�ޔO�=,��f}��c�}���펣���3���
�v��r�ѷa�=a�dW	��C�r���C,dNCKg1��]�y+4�ax����!ֆ�E�U2�OB�p)�6�f9�E����=�i`# �2\`m�1�q��TݧŤV�.%^��hw�^�bZ��{�����y�־(�f��p��Ai���E5�D`N�_�F��]b!T'/��xHzGH����o=��ڡUէ3�쨑q�9�D!_*��u�ZzH��\f��u��l�g�0���C�G�D��y�{��O�M;������<��9�:�6h|n_�aB.�t7A��år�2KZ:4¹�}��ܵ�����
[�Dn(ܢ��p�w�Qvc!�jUW��~ɔ�����3*�]*.��N�i!���3��#�W�J|�%�';ϋ�=�ӳ�K�o��,����B��8!H OB����bI)����@/4$�!I�|j۰@��aM�B�&9Tc�K���pU9�ΰ`aGn�S6��Kt@�Ԯ���;��ꋛ�s�r!`�D[�������B�����0����΋pR�+�k[��I�-^�+@�Oӭ]��m8Ů
�q]-�[t祼��9�\�m	�.Ғ'Cv�b֔v�Ԉ����+SW RYe�d�|�0� ���$i{���/��]�K
GQ�îX=T�xB�(
B`W�����w�!v�úOF�mE�nl�q���w1���U����`!*F������eH������,A}�u����[�]sfw�l�Ʒ�.��1���_^�=%�	!"$��&��t^�@�C�'z�
����Ȁ��@�׏��ٟ��5p�b�{t�@9�"�[�� 'n���ɜ��l�0��)���Ÿ�&�[�\;I�28Za"u��ɤ���#u�C[8?u���ϰm���	<�J��8ˈ���x�V�S�.A���s���?���G������ �\��+�w��A�rC$l������:"L'�_`pj�����'�I�ӫ�Gg��4��% W�cg F��)d�u�\f+� ѡVK�S���ʦ{QF�!�|\������A��ky勃�0��mE'M��Ek���֓�7��������2u�����dъK�J�4�t1�����LV�����ݕE�^l��!����(����QG� ��x�eH�`9Ŵ����U���<P\	 �� ��P�0�B3�j�卵=�,�^8}ވ��_�NH�>N���;@Gi�kq�3�7r�'.:6�4tAV��I)!���*��9��8
7ys{�֓���7�}	+�3�fQz(�C"8`�W����~g94V���n#��HChb��@������l�;��C��{�쿇�0`������{{�5cݰ�4�u�C���>�6)���Y��8��Z�~H�yv�r
�y�}�jń�9�[.BĖ�9�pV��R<,uF�?�ӯ�CR�0�=�X���
�ڋſq�ݾAT�3�'�g�VF�b�`�
���Y=�	n�bhp��Eo�n�6��*��5��F�6�`g'��խ@~}9�Glj�B��USE&0z�����\&�+����h��s�|�^�(i�ɮ����l�oղ�'o{�%P�x5�-÷��ݪ����p�7(�cQ��N��-3�o�e9lh�j\����t�,]U�s��zS�K��~ ��<�2ԟQ�;�K�3����"!ZuH#G��z�_��X�fE~˸���B2*H(�}v�M��L���O�Z{�RvW���@WֵV�i"p��r��0����7I���-?h �k�;�͸USF�w�`�仳�h@�NY�E`�E��?��S,�B��:�YC'@G�N�P�!Y4s�6�����ƒ�^l]��@Zv�D��>���X��-������p�T��kP�·=�x]�Z��|���Q���'y����0{.r��g��to XU��kkؼr5���ޒ�;5Y P�OTl*���'~`~�s���ۆ��W�`�����51]�Cr��"�L<;�ߟI�ѡ��'d[M��՞���!�vio|ت�������>�46�ԨѬL���	�Z��'�{k_в�����K�{mN��j� ��	�b�/�.�;X&Л8_PD���I|��� +릠_�R��Σ%��a�`��zԚ����g���
d1�_�o5X_�7���	+��O�/JJEćۮ����,�؝Jrq��!l�r�%D��j���KliVb�%6�'-���g,$�XXd� ���~O�o����LP�8��\z� ������dGz�ɷ�����/����A�?Y>��Eg�����Xg��U{+9ֽ������mOYQ�U@(�`� "�D�f��9������G�lU�
���NM�̈́ue3�@̈́�S��9/��ۃ�Vc?�RtY1�C�빭H$�}��ed�Hm�� %֫,�m���-�~����r��T�p�zOF4z�msՕ��uXC��c�!�ڽ��z�%ȃ>�~]�J�&F��w��1�V�}	��4 Jq�I����q&�f������l�7��Z9��D��m��y��v�VrQ�.���v[}{�57S�^�I��>_�;�ݦwK�Up����A�����ĢS�$K�E�ͩ�����뼒�h���`�q�$t��:��r�z��Jb�pw	���`�Cv�5 ��ɍ�� ��1���P\G���;`7��5�ت�- �ܯj���^�:�����1�c��ov��0ߢ�Ѐ�R[� �>��RYh��Ʀ�/@?�y!�V��=��~��}����'&�J��`�,z燔*䫸q%I�l���J��]�_�Up�h08�w ���ۛ$r���~vD}d����qAǆ���*H�g4��u���::�ؚ�2�G|�=q����?�2��%��u��|�ҫu�c��W���f9��K��I�����Mj�]`��bQ��\���ʓ]����8�ԴK�U���ˎ�� ��Zv�ɕ�����"�>�$�\����q��p�y�A�ނ��}�ɞ��eR���nl��]��������'�!�*���U�SEK��m�OK/���-�G���F_k�!�X� �.��7�hU�;�u���=)�>ʹA���5�� �pT�&��9G���d.�LEaâ�/W�G^S3�6RL�����T)uM/f�YujnK`��X�4����N����xV���x�����4��L|�u�b�����"��n�95���Pr�zz��*6~��|��ź����׷i�8L˪��y�a?�^�d(�EՅH*�j��g����Y#xaڽ#�0���� �H�fҀ����!X�9�s lm�7�t{�Y��A���Ơ��ɽ�����g����r�H���%�.��)�
��R��6��e�������Щ�̱���Mw����OA���L�SOyT�rBG�A�,��@��V��m;�IYm.TRG�\z,?�)�^ "?*	�Uȟ*Gi��!@P��_�ۜ4(�������ʩ_X�r�NPO��j�U�gPP�ա�NmI���B��M����k����7�CX~Aې���)�ᛌ��V�跠�X�,��i#�s�S����>�J����;��Lch�o��DE8,��~��x-T��
=AM# �	b"4C+�\�ɶ~��Q�z��\�X�͕�8�iE�n�[�"m<�#˛�7Ȏi���"IX	�H)1��,K6 �����/�Џ�u�G��۬v��rh��<e�z�5B5u����m�?�Hy�3L�80PZ?��,C`��_�S�Y1h,ĈeU�
����x����IYV!��#	�獢g�> *4�Ipr0���Hհ�{ߡ�v<f��FC�-� q���5�)w�s[5��K�uG?8|7�z�(��<�OS�5�~\�~����i�� \ﱙ%ъ��z������ ��˯�t���fx�F�'_�Pe!��=�����8~e��0]�C�)`��CS�3�o�����ě��ָd��,6-y� �na�<����4�4}	�̻�Ĝ)���T\S	�m��Z���J�2�e�0�h�"Rar
���KJ�y��^C��d�J`��V�	frC��@3�P��ZNL$�ȹ���r��H�?O�Ȣ����=�Gz�ȋK[]�%����do2_��a/!E���<4J���p �cОO@�$���8� j99^g��Ϸ����S�>��ǈ,�+���p���g|� ���,)�U{��=�����<�S[�i��p4���2���"����2�h���`�O6l)�o��	�����z�7�8�t΢�9���`�sg� +0r�˿���بw+�=*F�z8�zB�C[�cٜI�$)�:^�����%wZaL8�RT�5vMB®�8B�-�bu��'�;~[6KسjZ�_Aw�:f���麼R.�-��M!-ɳ*��\2��c�N��<b{iI1��@�kp�Aa�}H{C\g�P����F����C���G5jG|���3�qa�+y�����"S�R��ʬb|� �4�C�b��Ҟ��U�7��zOƿ�AH���^+��f'	&�B�`�⨸I ���J*�&���#4���s���٫�ū$�j���|�a�%$ᵚ��f{���PLoR���N7)��X�b+K0�4tv�*��$�)#�p��H�"h��������тemm�W�Rdc���
P��])�ں�/�	�>��}�1��s[nh��g�'лP�<8U����j��ح�ra�+tM ~#%�#U"A$��k����_R��"}���Ơԩ�Hޯ�'�O	�g�ɭ�a����V���~	����:�)Nc���wd��P���T�,w�ap�kq�N�����ǣ��ݘ]���VO�ݳ�0�}< ����BW='%�R����x�s,ܓv�_����E��۠S����X̘�KMMZ�#��=[�.��>C�ԟ��[|s���4�_�V,��RY�@[IjW
�Q���҆�`�q B��XD�.�#!�*k��qY�
E��|oA"���ֻ�xC��Î��X�TU$Ծ�jZL�j�}��������H���:�aо�'H��\i/�����s�EV�?CL��֒�M����͍]Gй�Y���[�ZE����N�\��d�"ct���Cq���5�dk��C4�Fp�ݠd;Y��[�@fC�岣�l(���b�2V�4j'�KRԬ��Hr���ژ
�K"�9��Գ�J�Y$F��oW�#��@�	�A
V�p�i�m5(�G�����f�2���ĭي���#g�̼�tX�7�l��n��~s���z��9���&B��_eF�VP��u�1�n��,�_M[8!��iS@�m�¬��(ro�ޅ���Ʉѝ}ol��a�$��{���~(���w啮wMو\5(�T���<��k��/j��9���e���  4���,X��5W?�;�'vF|�Z̺P$���$]򂅸���Ь_Bj�҉�٥j��N��X	��r�,��l�����Ve�����r{ɉ��3��9{"�#�����N&���2ط�O��( ����z���=��3�"��H��s�9�lT�n)8Zm���r*�C%=`����� ���������e��ˬ�����삋p���5���� G_������m0�8����+:{�|�f ������o�[K��8l�w�FT�I���ya"}Ig�([�^5w�&&O^~�D7x�g�?B���>j`9#pOSң�ډk��Z9w�+oa������W[ڤd����[/b%�v�r8�������N~PІ!#����N��ښ�26�\NC���9��5�����*cθ]u�F�V�i���*�<�*֒g�	�݃��n�`�J(�pVv�ߛ�P�.����g��!Y��U���ӈ_��7��0�]c��_��YX�q]��a}h�H�7�V����0[~t�Kxw�"���>;b��@���X5�E�ݧ��l�:���-�w�I�͔��Ujz75nE�ŵ~x؏���h��F.:��'r(��?�ݯ�>�i���V({���i����pG*�j��l�����,�B��G�4����7���_@C 7X �Z'��PP�X���nR�q�a���c���ܴ.U��l�(���	� ��f�+l@h'p�1�c�t9s�7T�2�L��J���@<�V��s7qFZڇqe�jT��D1�׻'Y����k_y�t��{���!*8�h�+�*��Ai�v>��B�&EEc.߄�+�@�d���u�����8�<V���w��s�_C��.b:��?��e�y��j�H����q��̀&��w�&z��#Z�3nޜ"����n,���aL���ג��DeV��#�7/b�^�<�8�[��#$���B�ni*ǀ>�l�vI�I��<�o}��I�fNO�NY�F���:�h�^��b�t���$B����k?�� �櫡�x�}���LSU�g1�c�h&�; �k+\����1<�N|���R/j��}�� ?���g��sS������<qG��n�-G�6;���)L� 3��`G����6맊%���6�s�7	%�Q�EU�H��"�,$�i�߳�59	��O�U(����_}��5�<C�U�j ���?E�{��
���L]�DJ;h��ݱ�'���GhǤi�:�"5'��˼�<����H�K�}!�p��IU���?1sQ3���9�"�?��߉h��s�����܉u�rc����*�5~p�i�Ta������[�F�I�{�u��A@��<:�K+k`�K��R�9��-~�I�G����k�DPܒѳ�q��ED�V2u��j�%ǖ-6�D�Qؼ�1��G4�K��p�~]��)�&#������aQ	���D�)W���[i ����^U���y��߉�f���dgW�D}�7��>H<�����B���HK��z�,�t�x���M���ICMh�hY���jɜ��/%�
�Si��N�v���P熚7������_Y�<�ilZ�ّƲZ�6�&�_ҳl#���Z����:���'�T{�Z7��8Q�W�~
w�S�s�X�-�P�h��e[Q2qe�$����V fjg�TP�GHQ]J�T����mf���L�Y���1���ĊCQRwI
,�V�5�2L���s���Hu�&7��3�8�̸z�;���D]ᬬ߾�j��i���R>.Y�"`�<��Fa��H�����i�}�s�E�s����n����9pEϵ��ڶ��t�feqt����b����]PG�Yx�>�󌈐�D2���%�W��p|c�IX�L���Y`�����V�*q��m �1��m���L{�.^�7d���T�<�i.�����%�''�}�����y�ܕ�j��a/��D����&F���b�&$~ZL��a��<��=��s��<fN���tb����j���vCm�A��h���08��|Br}��]S��/v��<M�G��)�3��E�yf��������\���'�p���i��o'_�������^����>f&�����b�Ԟw?�*���!ˡ;����� �F�bHv*"�﬒4<��`G�9NC'ʦ;��	�����|a�N���B(�J�NI(<��/(��8��ӌ��hd�2Ģ�j���uF )��b#J�u�POu&~8J�&е��,�lH�������eq� �4q��e��/�H�* [-�JNd�`�9��V�����<�2���M���4�םů mq��J*���z҅2K�N��N7�9>CM�������]�ƙH�RQ�y�>�8�I7����O�[���-��s����Y%_S?	��ǆF"+LZ��1�U�[+ �F2��n�9;�3��?*����*�� ������|K>�V���؝1����Cy�A�y�Bs�_�Rp������}H(��e���ν����v�GZ����H�4������@.��7�V���e{f�b$	�����n�)E�.�w��d�2�eދ7��v��Zxk0-sq�Uч��e�1�;`���%�%ʔ�︇b�#�^����T�-��?nPU"T��{���� I8���j���r����SZ�?��<Q�F�'�����6;�J5���0����.�nM�x9���}e%�8�k{̲����Ӵ��"`$���H]��X�|㟠j߾���2+���b+��.A6�<��܆�*|�o5E̋M#���?�
xqF����+�7����G����<;3�Ӫ��g�fM�������P�X��\3O���|"��2��0�>$¨��6�h���*�}/�t9ѿ$J�`�A;�;)�8�������̼TG��V�B烆���IfU|GV'^`v趨��UD"����[���u�C4��� ������/���zE�u����-`PL��k������/�#�	������:�V'8�[a�W9�.g���yR&v$�������e�O�� H������&�܊_�kr���)�˶�e���xv���f�lqg�O���m��xI����b~��jE���^�2�,�����8wnFdx���Oٔk��6^;Zw����v.�z0{��J�t�zb�Dw�GN���<�/9�:f���gV��M��D-���	b����^�C|�i2�X�F����"��Vdf� `���=�#�L�s@/��=W~eCq8�1���:��(���8r���*>SH	.�<�ߺ�lm��j�g8?�]�;���Pn���w������g`1W�]l2��,C֕�]�e��ɐTE]oE@5��n}d&�nS���fZY���68��?A�iD<��9=��݉�h턹�8Rf�yˇ�Yq�blU'�-��l�?��ud��"	3,�!��(�Y�ХY�̃'g�Me#���u���8�:�H̜b�`�Yg����!a(����W� \ �����T���Ik)YS�~$�D6b���&oP-`����λ��$m��6�G�����.@�ۥ�]����2��Ǌ��I�^�t��x5ћӃ 7?�'q�"�[(��*��>�e>꜃��W�;lq�K0�'_��	=�AҔ�������R����pl*9�&��TJ5?��q<��b՗UAXB����b(	 ��V��&�G%�Y/㐂����(2	�����:$��V��u����B�|Z4����Q��35�Jzn�/F��;����(���
��Ֆ�&cL*��?)���˭���M�e�J^l�ߏ��z oa�@/􌬂YW��M3�@���.�V�L&�鬪�M�0��_A��8<�l1B#�^��&�3Dm�n j��f/�dM�O��M�$��v��,�xM\R;|]n��2�Ϭ��'����:r�`��,������ī�j�tso�mD�1�p4�� ����=�&gM��%��;��Y��0�s})�6,�*� ��͂�|u�1M}�9��z6��JtQ�i�'��	���+�"���7<& ��Oq?-����/�g�$�YE�n��W� �#Я9z��!._+�����`���T,����uYF4a���mQ�%��~i�u5U<�Ӡ-���SNN��-P�'��rp�3��Z9g��\���z07��aGɚ`ΛL��f�	�N2
[����"�"hY �.��m�%���/��s��'�|��nˢ�n:Մ�U͠�v�?�}����}q%��ei�_A"�A�{��P�ؠ�H���-��'�e�r�|������Va�jo�R�i??@J�;�a�>��F�<���{�"�7���p{ �-��y^�2 ��X�z�<6��/��iY�n�*^|�[3���o��)�	4^SS�1�)�6Y������Т�	I6�L��T���>D����@�A�>����s�!,�q.ذ�h�TJ����D�ޛ��� ǢU@���:�W��R�8w�>�cJ\��U/�6�,������ ��Z*�!Wh��shע[����p���YߠF|~*):W't�����g�kW�e*�E!�����'`��N���P�l
��~`��LJw�����}1��U0f2L���?�zi��ћr�4��S:+�YQR?j$F�RF4r�.%���0_ɒ4b5w�����)����0��mOmN�=����x�s��æ�M��ʃx.��(V�B�����X� ڬ�qwz ������"�A��D�Ρo��J@d;\��.�쐞[�9�j����*�<S=a|��r��sM�fJ����<��5�XU��Tp؎�@�p.+��$9%A�7�׳k���:�̬u|� �t�&�~���fС��ᮋ�����$��4D�KS�u����@;�}<{����rO��w�z��،.G�£��HBĝ�r!Ѱu��J�F���Z�c��j�F��Iad�`�d�R]4C��sѩݽ��.]Gc�"i�X�5}�>�M�5����t�0�9���A�2O�_u�x�d�^��@^O|�"��?
�.B����{6>��6�iO�#��j�����P/����E�@�uO ���w��@:�\�����,�'AK$K۶I떈�ky��s�9 r��F��n܍��{ry���h�K�K$��XM���/�b�y��Ùbc��Q�]���s��˾\j��2v�"���fu2�m��6���i��	�gIM,f�~ �c2��6EPp��m}�(�fkT��[.���yi?M��y�N��
@�]�@��z��8�˗:�Z�%U{�&z��� ��턺�i
�k�{����߸�'�TP���c|_��Ҥ����`�&�F��)3
(� ��k�A�L&5���X�O�G��0�/$;H�쾾�wǇ��D���%1�*ֽѳ�Q���|��h��_Y���-CBC�ʨy"9N�xK���)D�ZZ�d�K�Cνac�'|1��r���uA=��n�+��	N,4/rޜ������Z��8��<u'q��=[!x|4-6+���i�O����9{s�z�ܐ�}D�Vt`����F�����}Y\D14��<�>���3`4�TR�#� 8^EBt���1R���4���Cg{45�~Z� 7�$Sz=��:?�	9T�g뾇�D%��O���F��t�/��!lK�[��ڍ)DS��׳P}p��Ł�\����ZJz �.dsф�ZAuD����P2$�R��Y�M�GV�2�T �o�X��=Fə8mC��	�J�S��vm�}SgIs^\/S偹Y�^�P���ó�щ�oL�vܕCms�{��M��n�u�cM9��ч���#�P�wR*wB���2�����<r|p,��2*p�&/[=�P� 
Qe*n�����ꭚތdNs���]Rk����t��{d�{J�MT}w�V&;dR�d*���f��Vuʝ5�*p|-�W?5�V+��ғ����k�GVA8�%u�]9Nl�4zv����4��#�S����p���4m��u�;��yVv������%'�&�З)��hh��F�+!���B�w��	�p����G��#���xyD��+��N���
z�t����z�l���!��j�1P��T�i���8�y|�{}��0��wN#��+��-�,C�P>C9�Z1�Dh�?��A���V�}0a}�'���0�����y]�z���O�
�B� �C�M��֥��`WD���buH�.*�t\��q���:[���:� �,������I���.�6��}�4��n��^�9a����2m��<�-԰6���3�߳J�u�5"Tr��S��䵬�/e��&�2B�.l��T���]R.����P��K�U;)�"?�)�3����B����?�jWsϚ:���-��3]>�}Z$�y�3k�d .���U,��n��Te��X�F���]0n��y�ڻ�3��\�%fAWt!�� ���К������Q��P  [J6m)��Z����#�
G�)TJ�c${���c��l4�S�@";!;�\���F��:�:�!|�٤�v�u� Qqj+����Թt�H�^yq^�|�/�B0�:�NEg�Q&����}�l�T���/LMY���T)Y^	��y"J��׹_3�3��9�|u&�@Y�?�hE�]�=�8��}����Ѣ/���#�kfxL6���HmW`#,{!���U�yM��̬�m?{���x�c$4�&�|����2�z�M�M�<��͠`���R
_N�������'�O,�A�����W��jj���H��;}d;�a�I���#dz�՘�W�k��ٞ�9[g ���� ��3��J�h�7t��e�*�#s����V3/|uP�d��'���O�>(H
[3�l��_=�t��E�f\�����p5V��c��t���0~�@.tZ��a�NS������E��9S�t��^�;��L��U\�~�J{�p_�q�y�Z]F���ʉ���wFk��>(g�S�h�����3s��F����#�NЌH�Bmcf�l3�����|5^n���!�8RQ�Xg�s-@���F̈Oܰc�/x��p�Ұ)���}�x�v�ی�G���ګ6��Wm1Q�꣍U�ư��
Z��@��A\���G3IU��#E����!�w0gؚ�K����Bm��A�r�Fj���ˋ�f�[fj�R���������X�Wc�����Q�"����3:@�h�����Ik}	y`����y��|���@�CG�!�W�0�N����(��0TNfM��ߞ=c�F¢���,$��3-�sԘ�J3|��ZS���,�Շ�j½RP�?��5�{�Y�'�0@����!�(��ۼ��l3�/�B���M��ɘu�_1�v����׼��1�`�VX���"Z	*r�D:��ws�g=��di��ۛ�����$�`��4[sF�눂2�E��! � �g���݌N���ۢH�L6"��K�y��� ]����nz�L}�r��2��V� �<�F7�w��Ԋt�jU�!����k6��~���c$���ГJ�lk��ʏ�D%C��	mai{��Q�c�B�EM�HA��m,9P̔_ގ�]l�UJ���}G�v&<�i᡺�Sޡ2��A >�nڄ�~�KK!Ӟ��(gco�t�:c��*R7���e������v����*�)Ѷ�#୆<7�ñ��M�H��as�Q'�^ߢl���2�-wQ_��K]�ʂ=�y�׾�&�H/.����[����I����Ȗkq)���J�C��-E<��k-7�#Ų�0%�	��z��m�p�λO&DM���z�� ϲ>=}�I$�D]{0{�5���䣟�d�F�C&�%�OԢ����$��o���DKw�֛��<@���?����c2��E��������*hm#�P���w��]{�&�4<�	�������dD�7*��,<���H��k�
�иy�:�}S�"�B��b��~��,�|o��rE�^�})Xh~5���uN�Q����
��ߞ
z�~�c��p����n��+Nǫ�.lNn%��I6�5��K��u����lf<�\ �t��E_B����8��p�ǽC�"�!��>���B�8Ql�N
���f����,M��RGg�w
�{Jk��w"�h��4P�x����p�kb�%RX˰��j�P�yߣgǫ����zQ��/�Mc���宂�^4� �R����\�Pɦ�v`qiMC���k��} r���!�����<pͩ=�0��iS.�l,�;`�>���y�H�B�H��K��h;[Y\�EYΕ��~�G�k �}�����u�św`�ܘ����6w�V��~[<�C��a(n<!w\X���Lv7�t�̕��A*�R�A39w�6R,L\K�K/�7������TL�p�7�9],Ҩ	=� ��ܼ� i�W#���9���4��~D~G#�u�zvf� �$��e�)g��9��L��:TU�z2"���ラT�3�}�k���i��'�tl��l������h9�O�+w���8M�xTO��Uܙ�d>c�I �s�F��r��du�h�pW���z�.�{w�g���#��Db���k�֮�����>��X(�9�?�e�*����b�����p5,� �B��]���.S�;A\`�I��N�ᱝ�	^ˤ�*��$�\%{�!��ѪJ����`�
<���=�t�U���z����H��zf8�]f�E�9q��]��ZD�*J$���B��U��->�ٛ$�nZ����|��a�r�)Gn6Pjj,����k6�]oj�C@���t���i��k����#���O77������ͩ�^�q,��|p�{��ׯDe1��_ӌ9�L���K}d[��GC�}l�ȓ�	;R�h�� ��IjT���^��K��,���j��]��v<�C��[�q9�ySfA2�| ä?��D����\f���/�0-�^�|&��n~1@wQ�Ƞg2�tl݄	�6�81��pqe�~ex�fF`A������;2颺)�L���R\�yP �&RE��;^f}!wa�W�b#���)->�ǌ�zV]��c<�q�{��&�mLk�p���ՎhQxZ`�����,ü�"�2Օ��O6BIKJ���T�E��䖧fH�5����}��(�$���G
$Y�`�剾
��uձ�ߔ�0' ��㪲 ���썑�@���O-oc���e��T�0O�'�Zw�+�R��_��"^M�*@�����a"�|"�R�&��O�kch���֓�a:�S�|)�P�����g���uO�ˮ�D��l>�D{UK�w��f�/9��^O�z��gJ/��G_'���_t�ɪբ��~䏸w���|91�j>��4;|Ǜ8!�t���f�[ұ�o�P��G�Z� �o-Oy�#S��������//��Ae�K�)���D������A���vAH�~�/v؎jz�d�T8��8���g"��������tR��i�м��k�X/��5B��I4
��R�w�-��S9�����6r�1D4���]�������:�܂O��b8p �06������Ϻ)R��\���L��4�3	X2� ��iPN��OѦWؾ�<dW�\-B1��b&2l�wR��y�t(�@|m&K�+�)k�X'��Ya��O��M������v �p�!RZ4�Ά��ш�_�9���ZY��i�r����M��&
��R;�.�zc�����t1Z�0GPZ
%�����T���+;I	@��:��Ry�k��`�y��L{��Y��$W����\H�w�f��H��S�5��8!
g�!(�K�����<H����ʴ�fDK��|Q�;\90����t	�n�%���r*�D��*�ր����ɮ܏	�vy.B���O^ B�nbny�v0U��t�2�_�h,��頼�o����4D;yU�w�X�2A1¾inA��7�1�n�&	S7ȇ`����P���&rX6�ʙ�L�H���-[&���n�Yxn�э�n�;2ǻy�ޔ�����d�Ŷ#Z�&��k���3R��ѐ��O��$-�Z|�Ns���\&��xp��g�-�n�Ϝ}`��W<F��w�O�m�Z{h��r5)3-�3��;��.��^|�y�6�hr� �
;ڭ:�ƣŴ������#��p�V>�����?�6,�G>a�6�L[B���鳣t+0Ծ�0��9 �Vb�ӊ��oV>�=�6���OԲ�i����~,L���9�	g���$0�l#9��#U<�"d��4�A�45cu`�� �"�/��4�J�0+��m�Qů��;1P":=��'�$��{���_�6ʂ���{=����^[��ad}�tߊ��[�Reu�V���[���dm��1j�	��a�ZYך�U���}����8�d�m�Ҷ�e�b��OqY=�"�h8�
M���������s�ywG(���+��X#��r���F�6�m2W&��Ҹ'7�0|��U��)х���s���H 䑤�e��UFی
���璼�ظ;��fCq��h�������l���\��H:�GC�qf�����:��]�|��X�g�%
\�ػN���U%(�/)b=T	�6<�n}��3�v[���������&�*��l��Ӱ����Y_j$����J\rh}v9J���;>S��3��++��
�%�o��>Ro���<58zb��.'�>-�@�Zg��厼��pѠ�Eg�9/g�����g�m�c,���5�����Z�@�. ���������Yؑ����d�Q����Ӵp��2��@�����2�w2���<g`@�>}��]6*� ��O��3�vE�F*[�]�Zv�f���,��n`����6)��k<�4��?�����(��[�'��@�S4�}���l�SO�o�WǓS.Wھ�e�ĩGa�kfi�c"ʽ�y����.w���P��������	���U���"�
�(|��܇��b�	������4+�f����O_��*'0� �V��|S��4��Oȑ����U�}���Q�K���J=)-m8��q���J�L��>���������g�P�\	�+��'$�ԃ�����	H%�v�Ao�/]޳�3Z�I���V���&��zs\,9o��!|�������
z��d�2��B�N��V�!�{�s@��/$p�h&�"Ԧ�52��c~=�̌s*l�d�P��A#�������2%��B�?ջ�h����,6�M
���oc�â&m�<����9sƟ��6����MP�	�<�s>K�t\������>4�db��	d����/Az��N�j�Nc(~�.���yjW6��?W849����#�z	IRhwm�į��m�zYP4������A��N��>y�W�=)�����s%��]֕�`Eo�U�!PI����O��]�z,�8n�N1�����[]���9��0�&��=����L��ĦP����!�]��n������c�/���� p�����Yb�~
�9��ͳ��Ĩ��<Iw�srhToޒ��%�,x��`6���_�������M˱�Н�b�{0�?�O�y^'3�s��@��cQa~l$�L�\_�2]}�]浍�ԥV�T�&o�ȎIc_��$��J'=]U>G�	/Л�f��÷H�۪6T@��X�#��9obj�n�v=�	�#�=��ˀ3sņ��i�_��)���;S6����������=�������vmҨ.���e���Fذ��Y�3�Ob�v9x��X���,��=�@l�������t�I�3/`i��Eɪ������5��I�ɫ�i֬�q'��F�����B���6�j�����^�(W�ߞ�zD�S�R	�6�
�	���mg�X&S)X�*@L�԰ߒ�T��S�I�d�tm0]�z<�Hws�m����V�$o�E�E>頻i-F��7(�`���߰�{/顦!�3�z5��×�{$Wf{��<��=���?���{��l&p�rz!=˃�c�I�F��% ���`�v�}�m��1�j�3�k�;6�[�O}-9ĸ"����ȗ�{,��PW��$~?��q������I�qb��x�eF���n'7�h��㗹V��q�7��� �m��z� ���G�H��'��.A�7eAS������Y�6��M?�{��u���߮���,u����8��@O���3(D#�� r�E��ٷ뽏0�E���K�!�µ�qĳ�u�O\���������}�� �#	�D�Z�-Kt����x#����DԷ��w������t\<������)8Q�P�,V3�M�a����k迧h��i��z�{�d���Ȭ8��u���c�2ٯY6�+����l�řt��(+�`)�of=IB��C3-
>Į8��F�Z}0�qE��d<�+��g��Eץ���WBc�r�#�9_��q�8`A��� dE.���hF{xѣ�\�n��;À/r�Z��R��. ��V���Q0?���tc��P�}u���,Qav/�7��w_�y~ؐnn�w�gܢ�D�{g>�}�m4g����;r0���i�����T�%b�?_�ON]7�]�)�|��ut�N�1��ʢrlJj�J�JÏ��� �B���'n������5d���cSY#.�t�V���T~B�*������8�����Nb�A�`v�`���L��Tufyo�)>� ��a�A��.��as)g�Cj�ӭAT�(���o�eY�/���� ��Em�˽ޝ3�ٵ�7�m%�\R�旎)&Q�&�0��� o�ID6�P��,��s�

e	J�,�7#Mݘ�B�E|:����\0�Z�yt3�@ؑ��`�~���,m�#��IJN���G�}:Իg��0�w���B�X��M���p鳽���`�,�?����ɘů�2`ր0��٘20�0�[N?i+r�X�3�K�3 >]�h|S� ��km�����J!h+�J���y$4����R'c$����^h��g6Z�aF_��6QJ���X�]�Q�)n�I��h��!L
1|�\�#�h �2Zzh��ɑr-B�MRhWԱ���s�sX�>�5,>Ζw�RZ�+���K�XL�x�V|�ēՌtY_�:I'0����;	J'#j��姁ExlYl��`�����n�9ڷ��>dR�fIn�O[mr
P/&�=�2;������z���9߉�S3�����HB9�����4�nsG3���$/��&\�fE�h�_���UO९�R�����4]ZR�wƣ7m���x�u���6=��y�י^Uݴ��ah�6��n�Pa���J�f	ˣ� �]�� 1T�|��2,*�F�7L��<�`�3���	LECY:́+O���zY���h:���da�C-C�_��Y��G�L�z����\�`R-v;�~O�ґA�d�.�������y�Ӥ+ڋ �H��w��֋���3�x�O���:RE��~��o���A����ь�Wp���6��v� ]�_XyE����U_��hN
AJz�#q}�Y��1�$.XDQ2 q�wU㍤C���ߚ��K�z��&�Id9�9�}�@�F�_Ű�j��e���n2xgS�pw@���A�������'v1�¦7ۓ���8�������ws�$ ��FA����9o_U�^�kN�5��-K|�"�꟢঑�m�s���D��Ć�,nhW��oHrց=�����Q؛�[�}�^y��Q81:��x�������	���S**aN�a������X[�L�����-w� ������?�P���Tػ~��{����l�ZQK�)h��h��$z2A�3 1�q����w�Hy�����6/�l*�;YE��,�GRA:�5�6��:.0a����fJ|�XYp�~/�� 	m�,w0}H�8�Up>6rP'�M�%T��%�[��P�a䯝W��0Ӫ|�J�xj��<f)~�Q��n{V�w�p�d���YW-}G����͢�:sV�\�%��A>:�����-�X<�mŒ�u�A���w� �R�����Z�^ֆu�1tG�~�<<�;d��]�]!Y�t�n_��q5�� 豧�G,�]�b�'"�}�>~	O
�Pda ٸ#��2	ݭO�e����'r�1�8�:�,S�	'����J����7�P�W�?�)�HUG<�/	5>Eg�5���^Ǆ�3����RS��W9]���7Q�ԅc� ���2CL]�
�yN����+������]F�{���g�	�W]�Y����5�,���_�c0�!עXS$��ؚ!���$*+.����sN��s��q�)>��F
z�g�L[��91��#���GR"dN*}M�v��{�� �n�lp��5#�$m�̸m�y������^�ƆlZ�:��֗�U60�z�_�>�9<��'�m��Y�*�$G�WӢ����7( I��X+*�g���0���/�az
:��A��:��	Or��P�,�cu��`��(�0L�Z�4�w� <�
r���M�w��NV�.Z3 ��<b
�ꨒ�I�t���|	��W��QN�Y�!F�m��k#�B���%E�:�P4^��l �VP}�ѐ�j�P�8��p}� �q�}���j-����ن�z���l8�H�ϿV��s�~�ڦ�~E^��H�v�J�H����9l��O῾j��wZ�R8!��$���×��ϐ�:$F�̭�q��7��Kt��=!K�p�4�0-�ĵn�a,�k1/�=# (�i�H�/|�t�
�߸�s�J��yK��&�\�N#����O����%瞰�_(I��^<��W��M~�V�p��l����)5a%�%M�`!k�h�*�K��%5���a�j.3��w����?�p&S�ճ��"ƕ��ȶ�&!^�d�h^8lj ��#����;x!k}�,U�KTzs�P��t���l����<W�w�3���w��N!3�����=�ڪ�gC��Fa���nc�3�X,�r��PSF�62hs1P�ć�(꫍���`+=�­�6o�tD����Ӓ���0K�(�"nOt́<��t�.���,�W<�sC9l��y@U��s@<�`:�����c�^�5�n)_����|���X�F@n���E)���h��r��i�<��z���R(��9�3�T�c����e����o{�������-(jt��]�!d�BiB�V�D�l��O��2m9|��~�v��PpW��Ν��os]r��\$q�ck��\m�N�-Lpab�(_�>7g�u���v��u���a�|+�4yx�<!.ˡ��-�"ER&C�M�,i�Ú/�:���t���:����6alT��V�O�m��4N��EF���t�)9o���5�����T�5�s���J��x�qb1H�r�Ch�kn��4j�t� �q:�����Bp=��✌�w�X(D�N^�C,v��EJr:�)�j�37ڈ���<�1�1h[ƎU�Y?���V'"���4�)ha�L%�*��ug�V�S3g�p�G�Y��@�����L�	�;����^�9b��z����R!ڡ�20D����gy�M���[ ;�M��ui:�%d=|÷�w��Һ!�&�|��25��X�I��M5g�����x-e
���T��F��L�4b䨆fp�%:��K�1s��������(u�ab��.F˙�N�!���pi��� ���E��6���pC�Eg����w5Z-8����!Jy +1֗7��V�_�
o�&�+���ꑠ���C�涔���ܬ>>�^`�q�4+�x>� �m�ׅ�xג*|�s�,�Ґx9	�� Re
(���	����?ky�h��7b��(K2�=��ȥ���&�m��.l�0n�I���*����L�i�TSN���/4&�C�)a��h��G�L�l&�.�S�<�^ �����Q����g&�^������H��SX��ܣ'��Yp龖IƠ���;K���ˀ���n���|,{_gYe�1��Y��)�w�d�K/ �ǴpP~���fQH��8��f���v� �����ʑ_9Yޚ*-��C1\�>�P����a<��ꐗY|β4�) &?�����n-`��sJ�Y(�{V*����z����R�^�ħUv��%���YN]R� .���8d�u��/��:�������#Dy^�G+���2#?�ʚ�i����X�=�GЀq�#dΰp�����Y�G�T�eӑ�����1D�(2���t�s�`�U2l٤��V���P�wՒUpEHE��r�H�|�����IΠ�R�a�����`����y�X��?��D|0A{�Q=u���w[�m��L��
���{(wv;��lZ*��>̐�ɵ�\��r��������W����֠�s�ǅ5�/��p��^�~^=)�e!��?�k�X�5<�&2bb�3ر�����Lk�IG~}�+q!�-o�a�F���xz�
��M�" SCW �dh~�E��V��S��]hOs&PŴS�}�倍�oV�Wy�����d����Rl,܆���&z�9_k�߈�ɵA]J�z��L�U�聶;����7{Z�`�iQ��5���,Heʐз7i��at�� E#�9�X�|ƈ��&�1l�ƿD�܈�%�h9]�l�fm�^�$���Bq��:ei�#6����p:;�p���^��;Cn~�6�� &�Q�~L����:,����?H�ԗ">¢-
��P�us13<�'r4�q��k~�!Y=�0{�^Q0����e
���{cq�ٕ�x$9G<O}n� hܶk\�v:(�F[�t"i�w�� �H�w�>�5���J�A�r�̛�!���z�k�;LQM��̜I2@�g���r�������eey�6�X��Q�;�ƙ�>�����+Z}�o(M�(�sQa�����ު���=>e橘(f�R
hY�Hh�U���b��y�K��g������Z"�;�����vreՍ�g��d� �PT�)���Móe/ �q��)J��.m�~�A�MZ�2������鵝��>#��G�]<����ރ�ju�W�6aL����=i�{�tD���7]���w�G��ɟ�w2R@����j6�/)y@���]2�4�6�P�?փz����+�c�y�� a���z��A����)�p�B	��V��x�`j
k���d�QV��A�;$�فl]��Xxh����0Q��Z�`��.
����6����C	�%���v _Ӡ�d����gj;o���H#Jj�=Z��g��}�Я��T�o4��s��"�4�]�Oq"}���ߓ-�R��~��ѡ��DZ��㛊����O���� d�7n���s��a��lN��2p	^�{2�&�s�����Ma�z�E��� ��|��W�ը��F& #9�������D��kr��g�X�G`4Mt�
�UN��Ƽ���<N�d��I��*8Y�f�����T~�a�?��D��_=0b��Jn�XO���D�_���j�*���Z�D>������1R��EF�;E�q%;Rt���'w0��"�\�M���.t��������^I;�o�b�wT7i%��6����@�o}�tm� �Ͱ��xe|�2p�9���;�N��:����%�[JDF�~�t�ᘞY�} OX�k��>ɚZs	E+�Ĩ��d�*Gn�Ki����͔�	PՈ�E5��$ȍ�Ä޲�4�	�� �o�����O��8��v?��P[�y�30�� x�Q��M�tXs"zd�Z�2�޴����yk ~OS�2\��E�B9������/��D������>	+J����L#�`S�q�b���K���?T8Q��@h��lń�C���q\{��z1�e�\j:���1n�*���8������2�Mb��+���X�{Ht2�g�X�;	"S{L[u��.��]wqB�)�V4]�<[�x�Pc�`���w��!����v�NqG Q�s���c�Ju���ٻ��?�~��nu��犜"D�un_�^7͂�`EP,+��v��+��r�<3�*�E'�zZ�Eʚ��. Mp��φ��z$���������d�%iՄ���m�k�fl�n�\(�Ԡ6�#F)ҩ��l+��������]{sD���=�OI����x̍5��i*j�*�U���l�eT��f5�u�����I���|�LYxgׯl-;\�Y��h=��Dxq
�Tӆ���&!�
�n�8T����T�{�D�J��(��=�$�	�S��xi���`��y#^��&�<�
Ƨ��0t��rZ3�E�g}���x��<�κI��	~@^��-B'�AGx��$�{�2�'� %?���55�P�d^�pp��zF�s2�>��ɲǃDwX��5���JY���xo��ǚ�߆�����ۄ�r&XAʙ��Ю>2I_�w��r��U�x�y<������=ʖŷ�$ltW�&����@1|�Q�J�Q.6����a�d�A٪��s��Q.I�έZ���k����{̕�S�^�W�	KH�\���v�"_�5A�>�r�bye�_��ZD�3�=�iLy�ǆ�Q CuW�S �m�ǝ���Ǘ��N����2y�Y��M֞O�o��Q*c�-f�T��g�:g��/�@I"��73(��cCi��ܐ4���J��B��I�j�*\�%��*j�Fp�'�O�G۷�u+/�����^�U�v	�517���[�=8 sK�3�����s�)N�e�2�@F�	.���GO���K�Gj�Aiy��4�EP3+� s�������ب;7�b��h_�n���@��y�"��P$s�r�����MH����y��F۫ geSc������Ԟ���\�a�|n/[��С@c�kF�c1V�6�F?b,�\��F���|��m����Qw�Za��{�>���r���!���,��������/�.{̖BS��!U>n@+j�:�1��2u/V�r��{��2�aswzq�`�Yr�(�NA����Q���౲����$Tk`��ȵ���t��W��J}KtJ0q�
\6F��o ����9UE�Wln�I��4�]�w�+�ڨӔ��7�%vWM'҂�ʀ�J/���{�d�5ko}�]��wK���f���X���zPɬ���b�H��o����Y��i?G��@�J�qd=��w��F�5/�ȝ*<t�ӷ<E�@㬀�e�h���׹28�m�)[?H9$޵]
����.�T9q]�֥�=�?�Jڼf��Ov0�B� U縘}��{�K�+�e����"3��15���n����!3OM��V�}��+T�=��C��1���0��Ԟj?L�[̰�!R �&�q�@��Q�=�G���T��N�@���y�������j{N����Պ�<.��={�|�+:b�j0��q,��9����T���d����B��S!�"�V=��HNn�0ٳ��c:}��6�e�0#��W�ˠ�G�����'w�C+E�y�l��\uEv���n���:w��������m},�.�o�f�I`���U�7Ҭ�k�j7MŠ��
}�n_��	̋VɓLp˪�Ua6���{ʅUU�в]q�d����:��i�������E}�O(�4F�����26@E��A���Ě�-�VW��qBQ�fJ!Nodլ��-!���k���Ŝ�y����+�Z���v_�>�3HƓ�V�����dڡ$]����Zu�����f��,f�x��w�C����%�!�PHɪ�}�{��]p�r��Pr�D��͢1���?�37�8��̀<q7'9<T]W7���뗾hn8
1�%���U!"� ��c0"DFeL�����mU)�b��N��g���Jz�����ex�+|��ѫM�G֠�|����Ź����Cj)u�@мPL脺�E��Z�~=����=x!�|��u̢i";������~�m�[�!
R����w�@�|'K"�t��%�/�j�l=�D&\�m��=U%!�O��J	��0�z�e ��ȭ;:��&2�����X!̐����IXǩ�aD̡��J����C�Rєz���:�T�n��*vn�D���.��7ahVe���pW���i!�|�=F�'ׄ{������ܲuh��Y0v��~�H1�ڪ0]>7'7$;b*s�Q_�;&	�j<��|�G��AHZ���������[�|V�����e�D���$��� KsUP�m���E�[Q��O�M�HH�V3�AŶ-��WX�}U6p�\W���<��pz*���B?��0+����,��*�	7tG�Ej�@DdRM}=�s˧ ێ�\7��b`Y��S]���˲U���L��Z�BkJ��*�_ݯ���f,�MB`�߉<.)K��^�-�pO�b��x�|�	vg���8�f���t�b�`�^ ά�غ[�K�u������4�3!�]�ҶJJ�@�j�g��7"gDOi�&Vw4�u��+�	UX�gs�Y���ε��K������{X��zoI9�sV��+�g������9�Q)EH�$u3����!&[��`��[+>`�.X������75�bR�$�Lf=tI�QGZ�^��a�S�^������1���#��A���\�{�bkm}���y���U7��_���s�BG�%�]��9�jj���<K}sdv��f�������ﵦ�b!;�F(L�~�b{݋W0���W�,;����1���\] �K�vyutoK 8G��:I�2<u+�)�G�Gpږ�9�������8s�Q [	�iF�,>�,�0oc��%X��a#=�*�O�yj�'��M3���+>�{�%�םcS�X�37�K�J�@R'��u��R����d�^�g�Ǚ^���B�eK��Z�.��W!m\--0!�����!�n�^Mo�GY����8���B3�?���4Q)o7�h $#_c�����[�:�Ճc5��nQĜ�xv�W���C�2
(�Q7q�Xi!Vb�����;����=�A���vk(H�$"{�� d���K��p�i I3!���u��`�Fm��p41�7���d���!��Ǚ��nh��᧌M
��|Ӂ���݅��$����+����$�I�M�S�L�|�ʌ/"R��Qϥ�l�R�}M�p�u���'l(�+���\I��* K�*r����l�rG}2��񣘰BҦ�΅5u����-�x����N��[��壠 \�N}e�О]��f�"vM�پ�᪔�R>uWfv��f�0`/F&#��[@�ڵ,=���F\R�`�O*��X%�x֊=Y	��Y~��Ȼ@1]u�4���s$�"޾�ͥzIv�y�����y�$��ofCi�E)a�1x��\���gĬ�d������Ka������u��v ��C�����	�?�X������M������Y��>��.G0I�` �E(C=7�߷��5��>g���r�`�P�Z�99��i3�_���t�!JF@��\u
Dp��UZ��v��x�{���m�������Xz<�Mr{�O� �����'uaS&Q�:�u<ci��ֻ�"���c:��{�m>�-��9ݎ�KOWo�,x��eF���H�ϗ`���p�y�h+�N5��I�^۲�r��U��9�O9�J��{hӢ��+&�=s�h�ϋrBgF�~�DR�m[�����,�S�G����M��q?��=�����*�Y����a��
<��>aUN�7�&m��n>���އ8dw� �$��H( �y�fl ���gf*.ȎK��3�3��D����/_*9�$Z�hr�È�B�KC-��b,�&��8�̹�Yc{�QIy�2����$)>g�m�r�v7[i�5����y m(��9����Q�O�ۅՋ��"c �Kr���2Rэ�eV"�^�k/��H��ʻ��-���.�Z=[�6��9�N�^�̫Ч�#�H�~$��;��z;�-6��7
J.��!��%jA� �V06��x���@��2�%������*��zk�e-��d!�=b��B f�X'�F�d��S-�r�'����e"2F�LTT��Z���*'q��s#{�����_#����{��Y�-�\��D�`[g����d�XGG+�嶣�����V�$�r(����Uf�⟐=�WC����>1���n�ͮc��s��֖��ID+�}��_"�
���.ZM�Ǘ�_��Y����͖��v4��&�C�?nekĹUۗip�a����f��y��=��Cw��A�M���i�����TpABm(���BU���f�����F��>$��m�HaZJ;3g��'|(�/��p;|�=��~ް��Vc���
n�-�΂��irU*<�e���&'��������Jk>�z�fs_ǥ.�����-ہ��%3IJ�ȩ#�X�X���|GX}b�t��qN1�sӶ$�4ZX>�T6�5�`��~���l��>��!vo�������ǻ=�1݈�c���o;X�)6*+{&���#.
����GF0�7g�(c[����`���~��\3B\;�7�D1��̆Ea-ڣ�z�9���E��b�?�xP�@8�]N�s�,� ���Z���$5F�O���fo�\4`
̋M�ᇶfx��K�s����1�`L��r��-�8N����y��_Z�z�m����8aaڐ�K���7)�	c�aVf@I�W���%YM�E>�S������q��i�]�&s 8=R`���.����Ξ�БW��޽�U5X$+���R�IAw�=�o�إ,�.08������Y��Z��� ^�������1~~ýT�[�[f��W�\�J�{=0(ҋ�2�bMW�E����hX�M�3]�a���g�f���ܛ8%	-?�*&�I:�|ΐ}����33Ep��X����Y{�7���@���clO��Xo�V���]�L���HeՓ��!�jT�e�1��6Hdn���O�i�U�o[��������O/M��iT��jS�j��r)���`;U�������*"�t���B�x^��at��`����4����MK޴���T��\?u(*7�Wߘj��F@�s�v'�O��c��v<N�I_�姄y�7I2�$́}`���R`X�����LF90r�ʹH��i��5*��d�q�hj7��[��1�-!�U=pXd�w��L�ꁛ�ڬ% �� ��R@�������o��0��Lr���

O(D��ӭ��ޓ��ݐ)�*��:1@��R���*T�5��6A�N���c(�X�[�*��t��*�Q���s� w�VYt�nA��n�6�w�j3EX����+�����n����.,��E�vq}?ibfcc���[���z^ 2n�O�8<��>i����Z( �V��<}�V��N���.�#���8߄�
�Fz��f'�1�7�,�V�$�j��;���W�I��3*�P�ԷC ��Ii @\=cEU�Y�$��);��кG-AV�}jۏf�Ϲlǽ�������[}���9�o%��$�b��@$,lc�6�n�	�䪘.?�~'n��/1#|�&�״����X�Frv�2H��-d~����[�)�+FG�Y��xٹ�Z��`�7a��w�}n�ٛ}燅i�J�[�|$:�p{�O��_'P|�@��*@���u�x.G���!������W�oM�t|�	CH�-��Y��\��|�������E����X�ON�����٥������pp�r��Ph�L�Lx9i$�Ӫu��P�O|-g�j���V�x�~9�D�3�GRIT= �� ̍�)��S?�@L�WٿPZ������<���A�T����@��oOݞ.���M�T	�s�=�D������h�Bd�m��o�j#!s��(\�>w?�:�)WT����� ��=�k�^������Tn��m��cZ��\A+����@K� ��,Ȃ`��D�o9�*������g��c�gFV���q��o_]P�+��~�s�v�?�to
�/�����K��X>2�h'(�b�Yb��]v񎨛��[F��Hw�6؊x��^-���3��u�l�ZN�{�+�~�a5�jI��tS7��з��K��ԞRz3HzfZ�]{���S���8ņ?+�7���u�3�*ǿ 8��6����|p��e�}��~��vm�f
�י]�"�rz�V���QoFP���$�1����yh`���0���P �yG�QQܞ�OE�k��d�v�ݿ��R�`��[��U��`%�Xo��l��c������u�D	�h��\2KU'��K:u��b�7F/}���?�g"�ͪ��Z�8�s�D���9_�b?#���7 Zn�>�_���֎�c��:�M*��/y!�y?i%��٬3Z�5�o$mF��%%x9���7��+́<�FGB9��,_~�tNՋ�k������<["�s��,0����=s��C����a��=���[??1y0��7�M9
:���%�5L/I)�o2�����������O_�g���*��=D4΀����>1kV�ݢgd���(f�f�th��xp,<l7��(���}��
�-B{F^����a����ς�	 )`a|F�M��uaj�; ��QE�ܖ�M�9z�w��Cz��9���B Βg��X�����ZV�Lݧ��5I�ER��v�"NJ�q�߫����Lvn�@wSS@���틶v���E��4.�I[/)�z�&bK�}�`er���\��⽨�����5᷆����7�0�+���k�b��>_��ǉK�����h1�F�u�	������$WH��ǱV�@�c�Z�8�� ң&Y�!sR��Ԉe�O�2�VԚ9�P6
���-���~�[���U����EV~6��Gݯ�˫����Q;�o'(OL�L[�BZ]�\}ߑ��WVy�$���#��2TY��?q	���Þ%ڰHo0\ъ΄�H3�_�N:u[�tIo(Qc1��|���'����ez��g����F�:�|��)FR�=��� l���H������N��*ά���G��x��Sk�$G%��H@�yoO���4S'E�i�!i�t-$���Y��\�?T<��9��[(^g��)���5����e�'�vE��������`�#)�*ѹڥ��Z�����Z�yg��1�A#ȖI��-��Nġ3���;�B�z�CeΗ����<x�|���]��
��c�H��WX�)k�8�챶�qA����ɪg*I�/<���im���"m�y	�&���ܫ��V� $K�@˥n���('�AGO[���ۉ��k�.�)O!q��%�3�.�R ����)Qs}�ͽ��X
��ͼGd��R�G	5;��殛¨a���݄Mn �0i_|�(P.�K謬@':��A旊�KE`����@Uk��Q�-E=j�����3Lq-��r#�4�Y��W�٫��&��SI��{n�y���,!����m�"Kr�"�O��B(��5��=�a֨<���*�"y=��� )q�����"P�t�0�8��'F����#��9σ��i��́#	9o6��N�һj�s��s՟�	2H�A|2��E乗Y#� ��B>�QM��w��#�噡�!B����Gq�cM�ƞ=�Z���fv�(�a��ېd� ����n2�y������ڿy�q�����̒ ��(|�[�N�{�zJ\pH�zP�'��a���?	۠/��m<\�-x��#=�$��$���A.e. 3�6��BL�U�wO�8�0�X�X�2~6�<��O��`�э<}�vTU=l#2�W�@@���%���3���i>�L��U��Ԍ�a�z�{�)��'�O����xK��>8����u��#ea����cʢ���J�n���	��đxx�Qq��-��"f��։��t(_�_�L/8����Q,p�!�b���Y��J��Q���umΨK�� ��JjW�F�� (�DJ@���~�i7AI55�N�A&�V�n�A��!&�� p�a��k����Ξ���Chn��.����v"wv�}w�_�=0\$��O|�y���w
�}��W���~ܖ�й�A�(�,����,@�B������l�W�-d��a�Ɨ$5�!���3����w0Cd�?6��l�p��g���P��p۲�}��j4ޫ�Rg C��=q>���SND�
��ƴ���LM�0Ux?
�u0< N��a�1��7GǳW�D�#ޚ�����g���� �g�s�o����j�d���,p6�H}×qb܅W{f6n��x0���g0��S�ť��FB�MG�n*銀eN~)n
�����*!��8:?�ET$ ��.�]XĤ��$���0��/fs-�"�)��B��ј����,�V�1�ݥ����r��?u%i���'5��d�b��/L$hqRH���� ᣐ��@���q=+E{q/��j$_��+n�����ș��swQ��PC9ĠV.РK��=�׍ﲒJ���<=S(Nc��9�]�V!��g�3�6H	���=k�p�K�V~�d�N�_��F�6��cZ7EtD�ݸq��EZw�O���o�k6mя������V�=�8Q�1��	�񴨀PE�\Թ���F5��zT��8�a^hK�v����`��(��}�M4#lBa?[*L]a���?z�G�ݳ4��Z��,���-�@!�u�D>��,�8�F'6]�Ï����>�Nɠ1c����2��$� ;��Tk�aZ���57��6]x�J���xO�����H�NУn��bk���8�|;�I�YT\l!����!�6lސ�QCuk���%����D�/���a�⃬�<mx�c7�́�ӵ�SE�Q��|R��7:��R#�҃��)z�����?���0=fĖ���q���2.�k�B^�	f��fu5b�]e�l�*�O�_'��SD�-��9�Y^1����ɸZ��@s�S��<�3�11�C@�����G/��2Q�/���z��?�*��M51S��#�#�-,م�O�u���ضqu_����_X1�_Y�� �㭋���4aT����$�S��QZ�����FGf�*O�NQLEꂷ��7�Ҕ�������9
�����8j�n��q锖JMdMw��7�	��;�E��L��s�Ж@�������0�P���Y�G�v�^�)�uWRGǎ׷-�]���j�xA��CF5�C+�4hT�)���M��CsIG88�ݎP_�w�*o%�,3��U�ϯ"�D����x� I�lۨ��"��YK��}fD�q/B�P���We�윯����`�V�7��c]�B�!ഛ,'��|i	��������>���WD:^i�˄����$�,m���~�E&l�G�z���/h֤4ɟm�^��ѧ\:��O�'�3kF><r'�gp�T�w�+�)!��C9^G��g7!�]�E���6U�#���nU��~�Q�t�z��G�u�#%��!_��f���ɽ�p���N~�;�c>.�^'�%�D�j�� ��#3@O���j���2j�GK�1������ڻ����qn�����eg�[=V%��"rT�T9�4%�o����)�&��c-�#
�;d$��%f�3a�1����
�u4�z�H ?󑗥�� ���^��ZiB�un�qR�zl�~�04�3��	�3�et��t�v�cB�m�H4�6�5��:~igS��q�>"�o�{
�bf�� Rek�:ރ 8'�1��l������=�3ݵY�.CN�C�&���/���p�^_k`)��Sx	5[�g%�BV����br�Qcj�jTv�c,$��p��e�Ոc�1�u�a�^;Ȕ�)��2�B�bTI�O�T�K2�-U� ����^���b�{�?����^�߯ D��8��^�qU8��_̀5k>�˭�g�0���Щ�����/G����
	��X+�f�Nן� +��/V�5WN�""^*�ѹ@-+G����[p����d}���`��rxo��&٣�C�'��@f�c�[d��p�"���3��b�<���I��ڜ���kV��_���ަ�ض4#puM#��;�L<�B���C���X�Ozn�2r�y�(���a��=�p�nW�[�@ڞ(Z�������?Z����Q�0һ���	6GL�͘g��7oo$������rlvzG]=�aC�I�w�'wU$��di�"}N��^�@�m�<�\�M$�U� ���G���f��ڛR��ʑ��M���ъ&��p�b~a��n��D �`_?}]�;���u��:~ܫSqd�*�4�9�M^)H���; ��Y�48
��>�uّR� %�UZ,413?@���e�k�q��X�������"��ԥ�]~�Qj����Ҝ�i?d�0���g��_+~c��f�ε�\I�?�}�ɞ�T�Mc�| ^;>i�3\����8��I �����z����r^E������o��N֟���i��5��É�TN=fS��9�3�5�dg����\:� �6��n��
�ȳ�/,V��HVwȸ��	\�^�"�ن>๯G�׷e>�s��
Z=�3]�X� 0�э5}��[Jk�W����95�K�"��0�c?I��$�����a��y)�G����/5��$ӹ��?a�u�>O��d�ׄ�����B�)�2:��s*ߕ _A���9R�m���)���y|9�N(�@��N�~�e2AF��� ���Q�����#�p�nND�B{DL����D�ok�͌�j�;w�=�s:�=7�/>9
��o�M���Ǣ�l���]�&��
� ���S�?�AV��m�$v�D�&�|��v�;�Ne;�Y$�X�0h��ބ_����_7b6$By��,�~�$�ކ��sΛ~�c!(�M�he�ӛɵs��H�;;���:i�&�H�T��*ޜ���L��U�����.��P��œ���z�O�p�1�Z0[`�,����S���Q�����g��L�Yʍ�pشR��6��|���]��}0�"|T�R�� :ӌ,���1�JU��ް����a���v�܃��q`y�g�����#�b��y��l[R��q=|t�&�+��DN_u�?���脻�K0s����V�6��Y�����+��_H�a4��BƉ.I�i����ט����|�y��mʱ��]p9�S�:d��J=��G���,����-�	v;���X�
�(�A�	��C��,E����4�v��{špBǉ A��m�P'��R�G���	tp�����hE;�V<t���'6�üm�O��/�g��%Q����M���G&�:p���(_���v��X$�u!,[� �{��3ej�J��+T�a!eB����?���j����|���� ����|	���e�#�o%W��;���ON�c�7}!gד}PD��"���V*@,�/i0�6{�jV�d���ɢ\��X�̰O�(]ƌ�Ě��dY0ƈku�"��% h����u���!��M&,�ͷu���`NHmw��������G��c�8�?�͵��?��g��~������cn�iV�F�˸:ѻyx�C1 �@HN��X��Hw�U��cyf$�M�IȠ����`M�8�ˤ^�C�(' ��|����0V\���G�m��|W�3��8!.

�Zإ���o���Ho�+��5^�bM��c18���_��A)�c�,J�7����͝l��E����Z�2U1�v�<��z:Ѯ G���Ѓ�x10e�����9�~x�����[��)B�,{�GR Y�_^������N�;L54��YB]�̌�$�!��"�:�q$�;M��Ĝk��]����8���˿G{�v�+����e.
.@v߶�u�Y�K�F��YXL�d'�?����,�i�R@0+4�\�yy��S/^���)\,~�;7y�B&~|�.?1x]:����V�v�y0������=m�LW˫K�j�dF�+(�d<�����/X�VR?����Ahd�>S1�'HL@�ʬ��\*D�j>�C������$��Cp��8BM�D'��kqb����N#�x���	�����w9z��˨jTu�ycD�<?u���C��(�4uz0�0IGG�)g1}��ZgJ�O������s�)�3���ұ�5��*�8u̥f��E:!�9F}lYH�AҞ��V���w3�^_5���~�D�܁J��fb9�`���" ��m��YHeܥ��ណ.��)d�t�"������H"^WiDa�`>��5��Q�Ŗ�4�2�̉~sɁ9k-�� s��'-k�s�y>��:+����X�&�]_��8����vrq0n�|�z*���4�)�E�0�F�ǅ����K�6� T������)+�afI�1�{��&�W���_���=SRҖI�����d����å'��MoN������-�>�E�w�s٭����~�-D1xt'�2-cm�cT>�T1�C�P&kA(��������}�O�fJ?/�%n}���[�s�Z�8p(���\�p��7GxfY�	:M�#Y��hb�?|84���s���J$������#ήs�s�Y�7�	f��'�iV�I��x}��	s�JI�XIc�F�>��lU��쨚r�l�elэ���t�q-S�*N�u�F��b�g++.��w���!�.,p~y��`-5��]�^7lxF��t��a(�C��ddaۀ���)I��.�[_`��Z�!�-����wl)Z$�̒j�]X�F�6Ihf����l=�PG4��2	�v!�8x���Zf�I2[c�-b��Zd��*��4=z����?�ؤH �t�n)Eg)إ桅U�bUeǎ�����ǧ���w��+1M�o���1��D�[�ٿ����s�&K=B,R�6Q_ի��=3��O��cIK.~���~��w�H���tN�H�p���=��f����f��<��cl�����|Cǳ��5�][�V�6v�B�*���Z��S�D-�r貔�	ս��l��.±�I�y"B�r'c�����# �:ׯ�12���/����H��u5ɥ��2�?J��G�nIbh��l�^8C�Ή�4vBW�s@�:�i,�G��$p<4Br����)➰����;D(��j���#<lE�z!=J�p�����/7�#QG�3������|l#ˡP�u�Pk�*rѥ9��b����H�`g�-F��j��4�襀�}���tt[@�*4޵�W� p�Ӌ_E��[c�_X�� dF��We!0iuD�ݵ�+���c��T8NcjX���3]���Fwn�[�3��S7֌;T�!� '�+��"�ʑ��x�1H/��{���[�!��aiL� j���B��ђu�
�O�$C��XĖѐ@�bn,�Rկ<14�<��%��ǭ��y��_�qE�El�N����΅��/̕����
�0��^�RkP��+�WL�&�0)��j �}�_ C�/�{ �<�`��]����J��.K�+�%a����q���֬�.�KCΒ���Jo�U���)�c?��i��|y�E��iه��$�O��[*��D����W{˓wv���g������@��-���<���=��0���i9�-Yn��2f���iR�ڄ�]sC?�6m�o���ϔ?�~ˌ�s)�\${�[�}fI��/.x�۫U�ZƄ���v�7�j����%M��T8>5K�][��Χ�H�c���@�e� �����7�֏!�0���?o��l\Vդ#@�彂(#X�����
����Sc�v6��%T��;O��M�A�É.f��6�����t���@[Q=lP�b)�@�C�\�N�C�ݢ�6���o�mC��S���'��F�����z�U�)�����MZj��<��@A�`G�PY��p���������%{茾�G��̫�T(ڪP$jx�z��:睚�����hdv�o���OL��r��Z٦(gX���sߺ=w�X��|~���q�7f�������V΃��N�h��v`���O8��s5T��@�����3�q��j�v�p�x��hd�
qr����y��lW�� ��!o�0�#U��lk�?��dV�>��|�l��!�{J�{�Ϊ��R�U+j�p�8�*.�����`�@u�����Z�� �dN���o�g�ª
�f�R/�ÞM���U��dO�"�
���~��!eHK��O'��D6^OZ��Ժ�ﶃhh5X]�~|ؿD��F��},=���<�ANǔ��I��
:dG���,S�Z0p��� s���$�ڵ��1�)Kٜ%�Ё�sAΙ��_����,�m�#��s(p@�cf����A4�sO��a���{f��I�s�Y0֖��Q����^u+���F�Q0���%���B��\�Zj��e�XQ]#���bD&E�YI5�H`��,%����j����\o���u��}纷�s����E�*��2*�^�VQơ?� �a�6�����_QRm]���XL��gPL�#� ��J�J*F�z�I���7��#�jh�:���?Q�w팯�
<g9� �H�Q�ĕ?���`���.TwK�4 �k:�7�]�Bf�����g5���{b�|sU��Z5wIc.�ȟ*�#�Ipg�0VR �I;!�C8�)W��/�Ô@���7�In���D_%m���s͟�e�h�h��<_8�0K�We����Ktl�0��'��M�$b��ڥ!��1�����j�`/b��akh~����͉w����V�	�ƽI;�76ȓ�k���s��W�X���þ���x�"�����G)tV�
��!�Kh qX/�JKa�,�=����&�)��7VA�����|
(�Z[(da��n�����d���(,\bvo�8����w����ĭ�+��aQf���l�uF�sMů8��ȡf+�nkYT�߫�JOz�OJ��C�.¢�R�z��qs�Z"�y��7R/��-<�ݚ�e��4О.����N�nU9Z�����XΘ`W�T��0����^t�H`F��$�Cl�D�8"�aA��8۲r�0ɶ����r�����>�t��<l ��S��ͺ-�mKj�g�m�Z���h�ơ+�����R��bO�$n�S���~��L;�2��D@�漊�ܕ��}]���.^�Nb˶�U�2.�Ƕ�A6�����M���9�2�P�������0!P(�3Q���629(@�� ��=�e��˗����|�Xl�O�W܊M{��H�Z�y�� ��w7#�O���3�B	�
·9�h����>v�,	w������rq�4k� �+���۰�-�����-a���ۺ�Wn`CW�#ú��-AUwէί��}z�-�¡j�ҮPDg�e!�B�W�L�G�1�Qذ�F�#�?��QeTzZ�ˊ%U���ߠٝ��i���;ӌ����W�FO4|=��9\Y wq�
�_+cE�0���w^nr�\+��n�'lW�t���G��A�$9_%تgѭY�0,Cl��^k�n��L��P+޸�������E�o9����'! �J?F���M����.�����8y�4�m��nŶ�����&�7��|an6�sT Ӧu�q�tm�[WǓ�&{���X�nȫ C��-�5�Hݮ��`ǹ�3]��+V��]��DO���*��=�)�üna��ƕ���Q��F�mu���DW� �����'5˵���v��!�]+�
�)Pb.���$ep]�j.���}��K����>ΐ7��x�QR�moi�q���odG��`�m��^�a��%�M��a� �L% ��K 8p��+�I��(� D���A�=^�mN@��� F�Q�@I�ʎ�ώ�5*E<�~ybr����7��cr]{?B�_T#?3W69D��-z��ǳ֟5!�
Ǥ!wB@,Yw��J�������ɎSVp��r���9��o7����Ti��	��'��K܈�wQ͌���]��X��;����
X�ĵ
om��D���x2l�zt�`R[�ar�]j*�\S ̭Z�v�T�Ƚ�H*�z��5���W�1w�1�ǡ�0bl�h�3��t'�>m�����հv���%Q�r���McNC�=n_M��Q���PD&�RmƄ��0�H�"Z�p�N�#���6Q�%��{	��^�)�%�'�WJ+�#��Bb��8��7��m�󧬧�^�.K�#�#'�$��]��"6d���;uA���j����$sǛv�T�
'߀�H©͗.���u6alv�+����eUp	�\�NX=�1�l:�=.�F>�a<���<1Kp����s+���7��W�)@���+�Z�%4��h�側{ٓ��FpD���BH�b� [�C��?��-��+t�3Ͳ޸$��yO!�(餒�Z�a�n��,�Ƚ�����0,]K6��Υ����Xcm����_�b/e��'�L�2��
Mq�fh%ҽ	YJ_<'F�i�$
��ܞdd�zƴ�DL
��k8?z�'�\��A��ͮr<$l�i�|����޳֢��.5�5*�L�澢{���c���͠2��Әbǵ�m�H�v�:���5��	u�J�~8j�HC�t|� �A��I�֡��B�VG�X�1�.��N�W=V�����f1)�6t��ʎ�y y�][Cߙ!p:�<)��Kx�����3��V��א ���/O�(��]`~�
���b}�  }�p}J:��1������%f�F�uC]!�I�ʙ�ѽ�̃�R�v��Kꫧ���o�[&�Sy=Ǻ�+#f5�Zj�nR%d�΅�FY5&��C��wN4Z�>����!f��e�w^��p�XnB1��D�j�N�e��}��@��^m�Y1`!�_�!�'���'a�����3�
�P��ޏI�痕�/cp���H7 .]E�cQ����|��Zx\]��o'��jHF����.R��W�-S�"Y�&�@F�w�J�����
�C�J�:�fq�w_�P��5�s(�O�ҭ���(�����}�r�o=I����q+`jw���t��{q�?<������0<�T� ��t�4
����H�̂�W�;�ܘq7�Y��H�Ŋ�2�ōA�ʅ���]z��R/��]u��+�VWO���4���K��r;���RC�68=��֌���"U�i�fg	cw� � z��P{M{@�R`��8�7Iҟ@���������t��n���y-
��]����
�<�G�\u��B(�-�T9��T&1�v����!�ЧU��Ǚ��>צ�Ļ��u�����>�ްOT�ɟ�|^���A݆ps`cj-2Ϋ-˻���d
i���B̅���0��*��tZ���`f�Ŋ��y�*��|b�l]�a�{O�˩Ex�,��W��\��5���h�G�������l`N��`I8�3�P��2���6x�'�!��T[�ʫy�K@c���Q.OL��K�薇���UCqp,pp:�;�>o�'U\H<20-��oi`�UCb��C3����?%�bF��|d�B�Ɣ��'��d|�g!��a�9�&ˤ�i;SM����5���YS�}�;O���4�ҀwaB�3c��no`��pĨ��Ѣ�{բI�z�]��ƣOd��n�n��!z�Ƕ�΄fNؠ(��L*Hd9�Z��F���������/�3m��W���\�am�=|��&J��.}T^��Js��lZ%ǵ@��A�쏱A��.Т�M�V���L#��Jq{h��'���h���^m�3��ı��V&+�������Ϣ;�;QY���©�F�1�Σ�?�;��E�<KP�B�I��e�(���%7�7�s]7?�&v�YjF��%#n����y�T�:F����+ЮT�-�)�dZ��cI�P��~�|,�^��S��#�V��Y��J#�@Վ����N�I��S,�YsW�\�i.��!�� 9��9�1|}����R]s_��K���aFq�:X�p���ɟA�T����2U�$R��b���
H[a�,���Xô1���ާjyl=�q/��bh��2_����t;�C��R�3J���͐f�l(�q@�viɈ�f�U���I�j�����v!1��29]�w �nJY �ؽt�����P*��H	�^a��_�4 S$�4����N%���.�)p���:��KKnK���)��d#0�᩸��C*O�̋�H'Hu�m4�3��oNML�qyיK�����*66���]�#@N~�rh��o�B��Z�7�7���|F.��q����6"���%����6��$YN�3���*�q���\|ե�TVEc��s�V
R2�t�#C��)��%C����{���j��L�qGQD�|�װ&�l�n�Ͼq�tà���9�3<f�!B��x������#Y������ض�7%�&)A�L��ʢ�^��q�����Jޒr]���gw}��ܗ2�%������y:�-��'[Qq�Ŵ8:��|�#�AI��>r���*�H���2�u~!�㔐 ��.
i�$Y��(WN�p����nl�d�Jd��N�cE';I��OL���_C�w0zCHΥJS3me�E�1^�V����� b2J�h��Y��:'+7�������Õ>�j��U|֒=ٟ�,���g.Q��t�b��_�^I|�L3�~��z��Y>�C�0�.�6�I���+g��#�K=I93� DC�Y���� ���F���
���{�����9������X16�Aj���Y���~��GO�<�p�7':aUb�_#�5b�,�0�n�B�gϥ;_�{������T �E�L��P�97����Nm9���؇��1
�eo�a�v�8���ʙ7�r��h����Ea���<z��I�bY&��7-3���|�I��P#2�͑�ssS<�IqƳ0�R�����%څ,��*��" pd������2]o����%��l�͖y����%d>����,~Am��/��v-��F\W�@Oܮ??`4nAO�>����m�:9_۴�wk���z)?K�𦢭�_ѹp �%�d�*co
���ں3�,�^`���s�Z�"QD���RCRq(/�$aB4��9Se���O�3�ǴDs���/��Y����,-x�ϛ���\V>uI��dJ�5[���n�h�LS�@�����W,C)�����`�Y�^�ɠb߳%�.�`�����3n��	te) L?�[l���^�3q7XF
���G%��iԝ��x�+v�����xy���Ig:�b�>����c��W*�M8<�e�Q�ď���=���Ǽr���;��,"Hؠ(){yҋ(s������?{�6��5eԽ���p��=��0���}55�5���^�h��ʋ�\Q��`�s�WС�#,1���t�Suh�eɌ6�y_.)�̈́&���}�����:��X��H����<�x����4%��¡��;�G��6��x<�Ѳ�(_�t�xȟ����]�\�S\��bS	���)��0ۉ_Y*D� �ݯ�hᆆ��1`H���`�M���t�w�F4p9�.pxϐ��1��� PV��"����^MM��:=2���4�m�=�\D���y��y���lc˰��_�؀@��B���	}u���5�����Ҭt�jÚ�`=/���_b�R��2�W�殍EN�,�W�]_fk`$��^F�+��]H�=dߵ��m������ڇ���b7���$�D402i���Q���a�=kT>فf�)�j�0
���3q���;rSk�<��)��|&I_[m�Z>��ӒҲS~#�e�LT��Ov�+91����+��l�S�rN\?��AFK�y���]t�`Q��k-4p���L�+2"�����c+L�4��]%$�&��Г"�#+��:ټ���0�'X��U�8{e _?�H�Z����48W�,yz������ףyx��+����K}è%+)���|�VpݽHJ����W���Z"��ہ��	+�0}(2@�~ʬ4�r��	�S����q�b�� �Դ�����C2����l�z�'��ʥ�/�������=�;��1�Nha�hZ�r��^9���J�i��Q.���j>�����A-�G�m�H(g��]����>mb(漮���x���w��-w�Ч�:0���OKJ|~�FBP���\Q5��V��ô\�P�T�S�����0�HUAi��6���e�< �>|�8Dg7u1ܛa,r���m�������2�(B\�����rc7���4�y�����j@�l�����v�uU���{{�O���4���d�����t�����|�9s$� "L��01mc�t�i�VW7ğ���}��Zr�X��tr�*@���]������:��su �LĂNs��RY��k����p)�rk�c�L�������D<ګ7y!��瓉�#.2���w6b)�*�,�&�Rȹ'5�3.�,�P�	PޯK�i�6�  �]f6�G;H2�Rv���H|��"�~��1N4i<��[TB���σ���yM���%���>ꤒPC
s[����q��<�ו:���z�(q�`��g�)��|��N�j'F�g�����F�zvv%z!�1���*)z���@�)��{��o/�^R��jw�Oߌi{S��z!#��@�(</���Y��W"p�L?w�����>��� �H���g}. ��7��B��"�;�~i!�9���o�_��(�G�[�S�N����kJ��%3 j,�p�i$��������s\
Źu'��r~�[4�x�1=��3o��B�\��T��D�mn���Y}��h�Q����Ak�X�r�\�R0��?�;+�����Bn��$���Q�ఇ�BL�l�W��
�[��BL��T	�;��IG����GÞ��x�@�'3N��'Y^�t�YA��}�{�r��"JI7���*oc��U��J'\��i���|
p�R/f�\�vd���Y�	b3^�Ć@/m����rV'�>�AM�dn?O�5ؾd���b-35��ki��t�)T�A�Z"�l�bEs�ܕn�?�j��G�VVx"�$c��f(�<QH���=s���o~����ߪoݫ^|t�E �����j�-��4�B�ޱ��x��ށdU��2d����{��~h�*ǁe�!�&\�|�X(��@��	.c�R��	ӎ�[�.�O�5b�%��ۤv }71Ft␪���yU�����S����f�����6]�E��k�*f�	��4*e��M��T�,؀67AY��'���B1-��'�(��g�]�,*�3�M�a��&���@0J⍮k_�̤��B�sԯm���I��Qϝ2'{TSaYl�R��ZX��?�����~��� �H{��Ok�^� �x�^�^�*��+��U;�����e4���9ζ�B���R!=ɧ3G��~8�F�^����"I�������KP�G�������v.|n��j�]c��$�\�x�q��C?�/������M�F�AF��	!F�:G�x^�+�-$ٌ{W�	�k��YK�
��fݦ|�PS�0"k1qx��
,a� p���V+�5}��Qt����uG��8��$J����z�9$g�����M���aWKE������A��e���,�'��nM�i����J :���.'h��l>��M�xXzU�,�V���s��ǈ�VՀ�n��(N�z�b�VQ1ȎL�ɡ�(v�TzZ܎j�b�P�u���U7��
���4�1u���Hz�ԸЀ������Zܵn�����̚Ȑ�6I���������~B����H��j�\����뼤��=�W&/O��"�(o��pr���װ���<p�TL�ʯ��&��!B`n�/�e@�����;�o��T���R8�����{�n8�J~ x��@��j�2�-*�A5�ܢ�._qV�DIؒS}�@������2��.<��)�>�+2�@_-R�r񵆍�/B�TB)�U��e�3?��rX'�ָ�ԁ�K��~�dl{'�͊�h\d�@5��lP����б�=�`Y^k|����ٷoC����lKc����p@��blUS��T�1�}I�pt ��;	7?�dXo��]�J3f$>���c������� �*��<~��)�$>���B�h��d�d%y1H=/W>�[�2�y�_��Ø�s��� &<EV�a���UK�ZXP ��h~eĥY�(�5io^�������4��6� �TCD����� `��Ƭ�(Ѵ�p�a����hu�vնx�I�L��O�ϻ��P��O���w5��j��H(��@�Ať����фc��hL<&=��.co���R
M#
�����������U��;�ぢ���������׸���L]�y��o���>��HX��μG���M����[}aϭsz
v/V�x�:T��?e�77J�0�iE���@~����U�0�?����czI���K�q�o��=B)�C���	��}*^WB����E�8�Z�N�L����%����V�еtw�(W�����,��:���1������hg�9)w�^ˢ��%��_��q�//��{e7��p �(�8:�<�A���g�d�,�g�l$�b��7]M�&x�'�bV�`B3�w}!�7�^	}+&bWr�	��,/xG�V������71��Ҩ(�Ew9��q<Cv�5��_�N��z�3�Dyk�����p'��6�[�a��@������Mӹ����q-�&>x!�FͰ�A�f��6��s��:�\|�v�hM���u�=C�!�����Ik��/دC|j��7rE�����FǄU6�v ����xbN�U�"!e�:E�����Z.�U]._��J�^/���=�/��
��I����g���zѣ��� X��>"$�|�+���'�I^�JL(��H��ul������1��g�*�~,�9�ȕ,���}qMvC�[Ŝ���:�#������/F"�M�:��:,b`�Tt�ʾ+�?� �R��S��?�)�ڡ�{w0xټ���_�����=���OL���<ͫ�;�2��er]
)� ��Ay݆q()�;�����U�S����S���Vs-��6)kA��$d<&���V6~U)⬒��{�rP�r�"�vW�����j�hډ�Z��0�Áq��GӤ���@!��R��M竹�ɨZ��7?��H�cO�� φ4lh�;�e�+[~+���~�`��A����Ԭ��p�,�X5�[������@΂�w-8�Cj�Jo�E��q=�=�$_���`�4���дne���X
����ŋ� 
	<�W�E᳻O�ý�
"�+V��0��|�u�E{��t7�ps�γ���=�z�����lSޒo'�p�,SIU���0%�frX��	��Ãg�s" *Ӻ��� �C�) �W)sa�~!�:5K�gZ���YqI��/Y�I��8Ԛ��ҳ�9���7��悪5����"	`��~������(5)9���}�F c��)ե��7)�Lt�iČc���� y���).�8�T��s];��s�^G�l�����M�0C|��у�
�΅�q[IRxn�F��qZ�E�|��@��e����2����E`�2���߼~]-��K%��2����A�]7$W��3�#bP��#Շӈ�؆��mw��_ݾNS��I�Tf��ؐ5
�'Nh����#0�(p���m`EGqG��=�Lv���=�55��;�a7:+rg�q��B��n��0KJs-{X�|B''�9`gW� =�E.�f׆!ՠ��jo��D�x�Qn"X>��w���Z+ufK:5�{.��b%B�������C��D��>)�f�d�ٯ�U�.2�u�R�Mr$ul͏���0�����C��8ꊳ�:�Jݧ%����V��Ĺ��Tޖ)���Q�/�;E�����f,�m���p��ݸ�>�5ݒ�z(�w��}�����=�'y�Ͻ�b15�2��8z!l�"[����vN�̷Mz'U'`2��D8�����h���|��xe�C��e@��+��G_ca���sϽTuA��������g����$���N�!Y�{d|g]���MV��D�)�Qu��F��~��&g=n���!`��� `w$ k	g�f;��6�p��ŨZ���S����$��^�f���fmQ"�0q�{�]q)!Jv�G�>����O享$wp�<+fvYϛєsX.s����{���3Vw��i8/H�yOX���E�G�IF�� �� M9���}E��3a���7���Y^�NH��6"�dY�ǭX���7��M~��0r���d�8�&���.'i��<N�}�镻
"�mz!�@7�GU(���O1 �k��,�.�]_�r|�"4w�&�a�Z"� �d��	��ТS��BU��Ⅵ��5zXgph�	��]5IXf��@S��ƣl͒��������E��j�i����z���}��O�����d���M���g%4P��۹b��]f�/V
�)�T��-V͒���`��氍zQ��r=�U��1�Q��jC	���P�`C���NrԆu瓎�������Ͻ����W�bf�b
��._uq%�ngs!-�U�"�h|��z�.�r�T鿌}������G�G�A��ꬩ5�FnU��5����'����[�:�a�V�cѡ��G��君w��T��t����ț�X{=:>�K��3�O��~���zfފ!�O.}V!���V�s��eS#>$ͧQ���QTP�%j;��s�b�QĔ8��{�D�F��T?��Og��\1#">9k�NxyO.�/�]o�HfA�Y�<��"${L%](B�u��R��	�I$��>�_��֮A�w���;�ν�lr�F��T�(�|����d��qo��Kl2qVc+�]�J�|�m�(�*�<Rk�d|T�5;*�o�ed��3$j)�1�D�'N�%z�7xً~�]�>'K� X1�ބ��
���!# ))N���2B�o{Z:��(!�b��Zs{�iS���Ř�d\��8�bO��o$�E�-F�(��f�Ϲ�N�탫����G�.|�	�5��V��� �8����FDd�2�b�i�.�����C���o�p���`y�3^^��@�tPW�(1*_~c�BNl�p}Am%�� �_��< ���T�H:�L��:�%�E������b^f�n0_�:�=D�"~%fɄ��V�8�������İO�[Q�_����\Ȍ9Z�p���(�=�\��D���|5����>iC�����hbd�j�R6�z��+=V�]�������?b����܁���m>�? ߹���	�_Xawy���(E.��A%�`P��ҧ	�g7��9s4��t�)s�_�w?�����Ο���}���2u)Oެ��u2�'���n-�y���	�X��QO�9�~�y��YD\*�<��X��2�� 1�;v�2A���Iֻ��ϲ�6�L��!�."�v�
�p��B1lTzPm=cgtRG�P�Xu��ClIty��ӶST����G�����
��@�NZ�6��ޘ�Ԩ���N�}P���Q� �:ЂE�@�䓁������Y��$(�Z��QW��D��?F�E��F:�iFsv�e�oGN0`0n@#[�*�Q*Xŗ��h�,9p�:GN޹�c�B�A�D�Q��q��h��F�� ��'��|t���$���'X�`�ֹ���0��k�?��U�T�ӼF����t�6|����pԉC���Y������E�����Q䂱Ou��0ͬiA��T�2�D��\�&�c"0^���40��9w԰A�{ݤ���K��|ڑ	M�u^^2P!gU��e����'(�$����;%�0���y�4����S�xy���>SD�T����SN�֣P��J~�����~��í��Ku|뫭�j�*��j��i��D�1�ex�N~������� i�&���Z�u�U�����.��h�y�YI�U�z�m巰�@;=Ah;nv��Þk_��c*���x���4��� �%!-�@Z3XT��k�?h�@�2�"2��*f�&ob(��X�S�\E��5�5�E�I�&ȉ�+���������N[a��i*��"FkN���L����?�Û܎����%��2�({c�LF�0����{ڈi�?;�Ck��[�	�$K���ƫ�0���'��h�k��x�'X�z	vz8��sMjN�9�nB�9��c��g�J}�&�#6ʀ3�:M荾���ds��-���Oع̌#�P�}W�P�����4���ͣ�#�+�ᵠs���Ƨ����N������]φ�d�k�8�gc0�� Ŵ�P�%k"�	�&��	Q����W� }��'���b�R�ʂ��Ծ@����'~,�&4��Cp1S@��X�Rk4:�n^�	���z�$�v/34m� �˺l��Dm	�:��)���ꎎ����(�V)�xDlVmj�C'�+Ɋ�=>.���}������(3%��~"�+"�*uy`����	���d�Z�<���DF�B��Lw0���R����&Soh��Gկ��+=g+�/v7Bg3�D�Ok< }��x+}W�.�ATC������5�)�m௽O6�0��դ�7#��D8��0PQ����>hA���%�������$K��M�;&4/�Z�0�f��փk� 	����ru:��U`o!��(�����(�ki
����`��0�����H�+���ȝ��pwÕ�{����΀�8E�Z	|+�*�C������Y�~�������� �_��,���P�	J0���x��8Y+�٪_8�z�Z��yh0V��#��\9>6�]��7������\���Fmf�1���~J�J�\A+��xH( ?�98�A)�'�ưB��^����X�q�<eA2p�u]�Xqj��q�u� ��f�Ba\z����u�����i^�㹺��V(Z'f�)�tDVE�M��\��4��U8e�]�]J=�fdp��l�<�Q�I��O��2-��b`jcn��_Z�@��+�0;��]�����S��<�a�0'Q� �UD�_���)�KC��YFh�o7�(�|>�$���d#D�b㵳������!J�g A% Ը.���8E���ztz��)wJi�����	<yڹ�� ʈ|׬�.�Hf{͝�p�?���<��,$�ɞQ'���(���:%ࡾ���3���;F�&��oyr��9��Q4���?G9����2evu��xȉ�W۔��<�)�d��;D��2+�F �'�f��L)�S�Q���w�Lχς��\����A���� �y��h�e;�{D§���~�Vo�%����H��P�4D�-N�}�b'��^�4�C��+���*	�س�KP���n�v����)盳S_�d���PL�
3�|!ݹ��A�d��/v���<��#*����L�t/L��p:"s߿�vr�]s��B��~��LqP�LF�kR���.���^\[6%eM
�O�(��8�>K2tt����K4~��(����Rc���ؒ��n��{fSd]��*���W ���~�Gaa��s��F��:��d�e}��?�������@��p����2�������p�w��GI_���릒�(P^��{2� 73�A 6�@ bF;E}Cu(��FJ����}Ohg��b6l!I�:��Q0l�I
���͠-u����]	؝��1w4����89r2�v�_��O�,��e�Ϸ3?�R���u6���5/SDn�$e�:MY��v;�9�)f�NБ`��}QF"��ь�w��=8��/�	��`�y��TH�@��=`��wJ����),�kJ�#6ܵw��)��D�{�f��˞p�����S�X�v�%@8�Eݫ��gK>���A�N�R�H�J���&�}�"Z�)^��0;e�RP�.��bм��Y�G z'O�q�r�o"�6y�3�U|L�*��C�6y(=�V����CG���� P���r�nDA(�Kܛ6b���a�U�d�a�M�~@�)�$�M���3C�����s��	,�hq&V#E�̗V���f��u����a�	�:��xU���E���ܼ��펄�+�����%HXN���#3�;�o�M�^hL�i�c�X' S����휐�/O��e�$>=n/-w�[�>����M+q1 Yy��ְ��e�}���a�3��`�݊y��n��{ނ ��
H�ޗ�9�	a��>f:��;A�,p=�[As�?�c��f�q@X�������K�i��0̻�ub�hxE��w�ٝ�b�h*~�lw��������*���v���W,�[B��PDS*��$z�8^	�^�$a�f���,��!;+��ض�:�� ��j�&��U�`��Ql���(F��1N�s��Q�&w��V
�ؿ]��K��49��F@qȣW��K�b�rN�A�-!��ʣ��5�F|���qb*�z�������93\-y@�c>\�ޟ{Fg`F+jCS�S��[a�E���g���U�F��1�^�!v�kW|R&�u��ͤ���&�eQ���=�]�|d�!F,�Ip5x5���M��G[�GB�m��O�Z�h�����S8��x��A���Rd�3ta�e ��,[f����X�K�<mQ�2���&>���%S0�`��j'^�5�=�1S-(��$����]�T�$1ĩR�|Ly=Ƿ��j�����7����J�n0w��"ڏ�r8%|j�D\������G�I��<�����И$�](*�q]?M�k���Q�3�
�l�\�045��T���Y��ʠl$-�lZSmu��,[�1���M�� $n�������?�P�p������|��9n�N���{�M��H|T��Y��D,y��YGr�$H/�4�΁�w~�'�%.�o�Z�3�5TE�^g�3�u;�K��3�vtu���+c��3���춒��阺b��pi�H�����pI4�>�E��_7r����԰%�C3^�o?}�CRĜ:���
�幮��Ḙ9T���Ny�*
��.G�s*�lxh=L�؍(�-����1����w��[b�kܒS�� �Fí��:g"���~�y�g�����W�'Y�+`��\�B�{dS���+����A��G�>��T+��F���H�����_;
¼,M6��,�{��C3w-Q�w��:Ϭ�"�&�)�,y�\U�婣Lt�z�7��O�Su�p�#`��P�_�j��q\٨����}�p�uo�Pθ%ݖJ\a�e���$Yf@��9<<n�T����Y�4��l�S�=���;�gk���r����R�ԝ�}(��1O�T�K�'"���Ǵ���/&�5_�^)����7�1S�Q������>�pw��660;�X�00�z Q�����1���Z�����| % ��͢`����`J��� m���Y�2�>���2y�������+�^���5\݆���3�!E+Px�=2��*��^؛G�%1�B�kM��[��aņ��΁�Z���������ˌ��4��`��lc>��{���l 82x���{��bn}�5���������M�h��>��1��|M � �bƴ�T�e|�VH$�y�ik��8��-���>��en�S��\JQM;�mǻ���v�_�l�j�ph�N󯜻�2$JsbO9�BF<;ظ�`磩iu��@�4J �v�G1w���)�]�E4�s�^�����OFtE�-�o���B����Q���Bx�@��W��*;��j/+p�؇D*��5�0�F�R3���E��TQF��z>@�A|H��*���K��lR�8� Ց�l���(Ҟ�?�G<������=���EAy�`��"S' ��7�~���*O�dI��QN�Ƞ���CmI�晞m��1E�H���h���J͒R�!����jb�����r��6���8'��������qM��N���u<��mb_\�~kލ4	S΃�[��m	����H%�g?���z��?�M�JH-�8�G�!�
o�lP)����d8=}�`�����N�Gn\4h�1�I�E��5�~�`o��11I��Ꙕ��Pcq�/������IY����\"��J�B��򯜦6���0��r�+�������Bܰzz�>��	�{9�����v~�3�r<��Y6���@���d��2���{�Ҹ=�0�?�ec��u���ZL�!��X��M^%yh�A��{�o-��.�	y�I*����V�$��~
�Q�:�ͅ�k�ly���rՕ��.qK =6zCU����A8U8���-bs�A�٨�Qs3�+~c��\�N��gImS(�d�# �A�Cs���'W�|6I�G0�@�E��y�� ?�w\��V��� ژ��{�$(^��!��CN�{9Oݹ>b���\g?�c
ZM���<��U#�?K��?�!*��Q�U�f���ޟ����J��<��󷗣�Dl��T����.��0=&�G��m��m�`?,�x{U��@�x��c���Qy1{Ǔ�g]�5
m��c�O�����< F���f��l�nhL�C��&{r��J��\�(�� a�Ө	���p{��m*�V�Nu�ߝ⩚�_N���1;�����1��Y�9��v�,�]����<��B?���m:��Ġ��uTd�!q�ѫ�=`�g�i��B���ʛ����[_�D`GG�e�^z\�p4�9Կ�/��ؖ=@�;��.aC��ө-����V�G��S٪C�S}��~<X�����L���@�v[>��}�UwI|)�+�h�Ҕ��NU,�T���{�w`��x)���F���&Pq9�l��"��!V������(����qoYX��w���W��v������)������A��?V�?գ�a޶���d��U�Jd$�(otJ��/ᦆ��6D��;k%��US3��K�7������ȮT�}�I�d�JFZ)���Ӛ'�&���<�dw���E��@�f���%.A�5� �f�|]m�Y���yW� ,�q5=�Ti�����pP:�������̪.s���4�VE}�Ɂ-��Ʀ���5�!�Pd#ۡI��~_��Ŏ�6+�}
�2-_��vy��,/>�}XX,ڨ�D�DItF�5��'[9����+=�-�+O��ʃ ]��F�q,�e�ܽ%�w *$C7��'�ܸ|;����ik�#9�q7~�{MQՊз�g8@�BTs���0]�� p��P��3�C�}�a��HZ�<����T;\5b	l�Xg0ҟSG�֭�3o��㴃����� \2�(����$�x`� J�V6W�M�ۦQ@�����
����^��-�s�M{酧�Q�VXu��Pc�C2�(;`�& ��,G"u:u3�{ �=�S�P~��]��P�	T����Q�M�7e�{��>&")���5�S�0\��hۖ����[�9�����9���h]�T�l��	�尖�%:(�g4m_*�
���I��Q��<����xW��e�q�Ҷ��Z�m�n	��M�z�|�����>ί��P��
9{��h9 ;�(��~P-߷TP#�\�w�J��oT/�8���e�.B�("�1u=��˧L[���KȺ�D���/l�7^r܀5:��A��'�nuҪ��4���\��U��ʼn]+iN9�B:��
.�����f(%�F�_D�y�R��kKJ'Vy�tN��`��[�F9�Dw�)�EH�-�lՌڝ�et�5�� ��{�х^p5����Q�i'P�",�����p�Z���ƍS��sT50q ���\u�
-SP�)p�U!��쀋`?�5n(��j�HR�"k¬o�����:��h.�'�.������ �WHa��� �v��^�N�XfX��x�#>��)�C�]p�[\sI��U���J��K�m9��L�c�@-*"�Kl�W�a+8u���$\�.0[}��0�nY0�������uvd���l�G+��Q����*����?�+O)W��������;ƍ�=BQ��^�<��~�2���h�A��*�;�e�����}���"=bT4��^�R�P-�$�ı���W#G�CQJN�Så)�3�!�/��{�i'g���j�w�ś��2K��5��Ǽf���3�t0���|�c�������;>�#' �	��� ��Jmt�+�+1T�j��i�CGl~q�5/��!�����'ek���k1�la�-4l���0ɫ�28��6�Qr�<��GK�|�AV:��-�WP�{x~T8F$I�"� Lg-�����e~�e_��ɉ�$h���5�٫L)�i������f��S�
wg[Bx���7�Z�O�t�Ѣ$������ޭr�oH�/��0�G��t`��#�`8�Fۛ_��9�N�mL	����-BCmL���'��Q�D([��P��9:Z��8�|&2M̓H�wTIG��������>N`�u�+=i���Z:	�����/>wj*Ce+!��>���k�ҹ�2�h�޽��D��J:�'�`��U0��}W�L� )f��m4��1���	��x��J�|E�V�����f��/F�k�b�5���K������{bnE��.v|�5����0�����z�F?�s&W:��(�:F��i�q4@���Nr�|%�4�:��v�+m&l�s�m�ձ�S<S�[�P��u,VMx���%��ύ Fm�c'�ژ	��<}Un�[j�}�`��")��b�2h6���LV!�.������q����7_'�A2�s/r��"�3D`�)�l�Q�
�f�g���z��<�
	��D~Tp�@¼l<Ɔ��Ǝ�����v�����I@�e��<���}k�'���Bj���|^��������7�}�-�C&Y�nO[��s�d��\�ga�1>�:�V��k˃����[&�TK%r3�{t���G��W�Jh���ұ?b4y�U�ܵ��3�n��1�D4�/N�8�#B���;���<�8D��5�@uO��F���?	5���=�ZG��a	��ĶΡ��&6�9面w&��0gH�n�mY��';���7J��D#��Z}��}匱�	����s3Ϩ`�[�亝�D�	��Ѝ�?��o���4AY���S���PE�1��w����l�W�;�$���T�Rr��0|4k ������*�<P�!�5�A��������1�X��P9韀��uJ�~�ف�|���Z&��Cbq���������ja,�A�J_3��C�s,+U�>�"��x1��~��MH܌�Df#��[r�ـ��}���Le�d��z'o�d.�=�J�?��s���Z	q0�_�|f
�u˯Ůt({SBF��6�.C%�iJp�M�^`��8���;�!�<��������b�,�2����r��I)��.�$u�0���2��؊.����m/���Q��r�H�cL F�s����L��(>��p?g�ր$j���[�S�;�-�7��jc��9sk=s�!"�̺��|E�'b�F�.��ᛳi�Qr~p������4�ڤ�@U`q���U>��.�Zy�,���m8���e�X��&qG%��&E�뵾�zJt*�[p�;��sB(�g��MI(�:.���cA�����L����4.�5B�?*���)��2�x�.�8�V�~$�)���^�A�#Cȑ4�!-��rc܇�)i��,��S�����2Ŵg4�Ů���)fZ�㜈)�c��갮�`�O�k y�'�/�E��!	8�j��׸�� �'�ג�H�S����$�mF��&8!�U?�[�� �)�Q��ǫ�\�6��!O���\a8����#_�'_��Id</��h��2���a=0-�]Z�� ����4m���o��bj/Gfj�f#��80m=P�L�p�{��.�ɿ��i��.>.�+��m��/�I�=��7����4��IqD�3Z`aK�S{�����s�O����=h%/�:Ϟ��QY#�@�r�:�W TҩA��c'�h�Ӿ����4�9L�UO_Ri�rF6��!
3�|_��ۼKo ��\HF_^�]O�8��L^W=~�p�=���I�����?R*)=e�������\�4���q�ՙ��f���� ^�a,�K��1DpZt�P��T��fL%����ƶ\��Q�7je��M�S̳�C<��P!�3r,�Sy h�1x!�E�ZϏ�|�V�'`���|.�3�z�E��x��r�∍)�84_���H(ʰ*����g]O����L�ꖘ,����ܸ<|�(���k���V��QF�z3',˷�ڹ����Eѷ����g$�˪��������C�=?�Ԛ{���1�ހ�e[�a�\��I��}����w�TFMXq���~@؋Gx�ԧ���`;,L�]�=mv�����;�< K	�sr��m���v+�]���@
�[��}Q>6�eڤa(�g�����o�����$r�)#L+��l;��4bf� y��T]�[���IR��}��	�����ۆK~���x��u������Z �q��q�yhv���]V���\K�����"ȧ�V��T�SЪ��$2W��LR��؞ks�^���+���#��ȃ����>}ꙏ�,�+	P�6�p�.`(2�b�n~~Y亼'cI^���D�\�F�9<E��GDN�N������SEIn���C�6_2N�w��hg+�3���;�`uD�'\�ˊ���?B����Vk�����ݍ<ar���1�2�haBJN*�ۡ��Ks6�acrN��8|�(�:C3ޭ9^�%���>�Ta`X�����rԷUT����"Փ�������� �G�.h����������"+�s��n�l�s��%�臧�Aԓfn>��|8�#���|��w�mB��
�-��zYT����|���c�����co�8V!ՇM�1?�凌�����gV�vbj%%���uD�c�Y�z%���u�W�\5�]�9�j!�r�i�V���?�\��
U�<��P_w����Aq��.�hm�d8�D�!�q��M�.r�Ңi��6w�t6kF��Ohӏ.�^|l'��X���5�
��h������xH����ي����������P�= o?�.�d�*`� X���s}��Nّ�"�T)�+��.I�cr��i$��%�^��6*N��B���1^�����,;��L��%2����<����%�[�:���ʏ�Z�~�in��O"Փ+P�����ְt�h��nAk?7+�N�t9ݦª\9禠J8���j��[|�]�]��+�}�m�as�!|o2��/&���/PI��~���-za�?�x�5D�G���Mո����� O�A���*�k���R(v�b�y�I�TS�*!������M��s9_r�p����&���*v�d��2�ӧa�\Fv
�ɓklۯ\L9��ǝez�����i�A:��[T|������o��M�<ٝm��I����+@�l5��~��dn�Ak� ю�7sxP����@!��߉��,r��·�8���ab��ִ��O�D:2�޳��?�ú��<t��i)gI^���,>+��n����_�_�����2$9'�rt��6up(Ma5��"y��ʻ�OCg�"�����ք���փ���C�s�ӿ:�!��˼�lW��شm��*s��G�X���tٿ��2����JbXb�2�1?���a��b�w���K�OH��`�Z}�q��wB�A9��d�:�e��ٟ��'
;V��X6������H�FY�G��q��؍�#ˠj%EP��#}������Sp�ϾD\E�z����ښ_:�b���
�{ O	Z�1��<.�A�������d�*;(�=�"���v�b��@�97�vaEj��XI�����;p_Gz��B��?��o���X��n/�B�M���2�Ix��!�B�z� S���`LkC��7��VaHz�ԟD}-���4�Q��~0E���Q��3�x�[���$�����ֳ�0��^��-�h� �# �=i�@D�r��������T�^�q��T�Ǡ�.�{Gy�n�i���:�I�4={B̥D�.�1����X�㑌J���F�⟙*�,ްOfM�!���O^��ci[ ����Q����1��yř
����Gg��<?|2��)vN��f�<�)��D��h��
ϕ~Йi�)w*�,��s�-e;Y��u��E����v�_^.!� �Q���o���f�����ѣ7����i/�N��=�����jW�
n�����st�$e�∙��gVY�����t��u��~���G�hFS�ʫ�cb���+��d��>��r%M�ٝ�k���춊���y�^����܋���֓)\\_Om���F��H&��qSCa�;h?%c��ٖo@��]I�*_Hɛ*�,�cEY���[r��7�^�`�uz��th���w�#	�2�b�FT�pKsZ'���GH{J��܏��
�[�No��D����8*?� ��GJ������g�ɩћ�>S�~�lDj
r#ב[��/�#���$��+���Y~o���¡iZn��zF��K�򫰍���|�i�Շy�����?�)dާ`�~Ϩ4����/x��#<�MPdD�b�ew���h�nZ-[��xB�m����*X�O`±y*9]۹���@��[�K����2	��b�Ǵ�=��(�ÿ�g��$Y�-�.�����b�W��Œ����������L~fY���X a��R�e�mf�7oY�H�-��s���]X����!{�elW�o���o1_��'�:��� ����	#_3f/�8�)�>�~��Ip�}I�&^��60��*��R��FՎ9�����Pm'�C%"���:j��&�D�/ƚ'
�Ն���0��'n& ��L�R����UӸGXpG�k�����J
�:�����{;�I��A��LSɯ`��|6�B�d����1��-0�����fy�O>vlIx���Hcyh��}qC��н;G�l��d��D���3���Q�)X�'�W�h�=y��٦�V(Eܞ���p,�s�}}(5Z�WQǙþh٥B,��G�]V�% 7jV�
q5�Q�לj^n�=]U=�߲�M4-�{4a�$�퐼$�4�Vԩq�y��>91�J�����������g�5�jҘ��Sn�F�4aw2J�0%*���K��������%_zQ�1�7�'�~���	�Ǳ�p04	���zOɆ�qTe�˱�K%)��>"�7�\�:r~��;��PX��s47��k�	��J7�����m
˾@���Ͱ-(qFy	�f|��{�z���:�vğ�Ɲ���I���J���?�ZAXHBX][��ˊ=�pZ���[�|'� ��1�Y�1K���5e��g��^���g�,�ReM�B7"Gh��֨F�;n�d�D���7#��i�����`O��ʁ�L�e��Ф�����Z��A�~���
��'v��R&��wg�R�޹/��<�s���kl*q���k�og'��-JK��jmzJV��3�WJ�Q(��c�����0�V�S��b��cJ�g~�՜��f�-�=ܖ�r�J�V�:7#>�w��HSſ�!�n�k/k�4_"<w�V�q72\r5�ZFX�,X�	Mӣ��B<�t�11���n��;7��I��1�"$�o�
��>��N�i���P����K�f�8�H���]��n�?�`J��KAG ,*����~�o�f�ӫ�8�2(X;��3X��[�ߎ�^���2!sUϧ�[�Y��Zp9n�x�M�ʵe�� ��$!�-�_�Eɨ P�$�����-�L�{�cސ������T�t�$v����0��Q#�_��;���<ӤmW����W�m������2������r��|vi�ʭ@�����:�W����3
���|�<47�j�2�������-���V����öega�`�	�8O��h���6�ֲ�R��<�Lc�FY7Ф�����f$x-�D�J$�I��ĶjK����*#s�o5z2���`OG ,���ϕI0�V}]EQǌ5D��V/*W#a��1͑�Or�׺L���_2�!��./�p7B��-q� �HID��_�F0��#2V+3���B�NC�	��rY����'7�r�3���-�.!�Ĳ�9���!�*Ta�)�}�cz��}�ߚ��O	:OO��$��ٟ��T��Rf�_���i �8�;�ҫa*���%w�'����J�Y�[�y�$I�����%nd��$,��0��j>�.-!�J�~_���3�韱U��ſAň(3�oP~�Q�y)�����4�F����KL�A~S��o@��Gs�ع��5{�
cU�R�~�7a���rD4�������^$��ko�c�S4���^��w}���(3擗i.$u��8V]H��lV�]0+�Q������g �v?~��4]�[F�,k�B�o�}�<���+CN.�'�ԮG�;J[�}1@�y*kǥI�F11��	�ڪ��Ŕ��χJ	�֌qa[�^2o���v�۴y�/$�p|�pF�k\P56mHPO�����u��y�
��_����d��a�.����3���'�_��-~��ǌM����F2_�Az�5�%�M����kzg{��?�)��K`aW��䒵!\���2�G��h,��\�q,���l8h+"q��7�u�a����QGpp�	}f́?V~\���}�� ���z���h�u�_�� l��fv3��C��h-mW�O���P �C��`��=n���Q���W�f9�Bsk��=��up`W����+�K�`]k:X=����x,u���SȰ>�%^�@�?��Ϫ���*��O��i=D���7ۊ�Fg��l�"�=�Y�(E$�����5}=hז=,3�e?���5�gx�km����9�2�&�6~��ؾ}��@�P�2p<��il$��gT��6�Li���#��&�\�����_?���蔘Rֺ̤���ۅ�W��N���vT;
��ح��bk�Y��B�5$��֕�7*�f}z�Z��1���񻔖�k�d�H3�9�k4��7 �����D��?2(L&�ߊq}��{cLGF����F��K�P��q�8��5M��0	�2W�0��"�0���}���!�Ev��o|v�%��<¼�D�I���}r�ãk|U&}~C���y�Og�� ��8�B�-�!�ನ%O��W�m�� ;
$�h
����r0�6���hv�#��(2/-C2m�KK)5����bH��L�Pű�zgcIv*4o�����u�^9���N ��i��e�CQ�U��ݷ�H��U*�G-� skfr�����N�jm�FM1��{�v"i&4��v�L��Q>d�W�=�)��_Ã5�C�C(h�+��ֱ}te�_�,�]��H\�5w|?R���)��yv��I���W�&�(�6of2z�gR��4G��@2Ex��a� �ĬpT��f═������9�!��<�[� vK��:e�,ـ���d�	*�?���ů��	xB�N����X �����^�q$�j�3l��̼r��u+pN��[����Jb)�M�Wn�B����������kN������&��(���|588�By�6b׳(�NReGVo�r�c
dҤih��MY`�S�fd>3��Ɍ��>t��앫����9�U�04�2����<��x�N�Q�*Sn����%���N�,Ə.�_���?�� ����aAK�Xư$�<���������8���'W/���4��{$�͏���߶u��ٶ��N��p u���l~8�rg��&���cM)�4�!!�����y��S� �+�{����a���cVl���m�ҭ$q�	?c��x�;���Q$�c>�Bww���;�]ǔ�w�T�d�����|Cu���;�-��đ�A�j�˸��^�N�J��V~@��V��H���D}�'EKd�@p}�U����58tC�ϭ*�	{�	B������rq3����}N�!�b�0QdF��d�c(�{�Teɝ���\���_�_�J^
�]��$��T�EH����2QO�U�%��#����A}��W�%��E���\�V�Vy��1�4�ć���Ճp�9ŝ�a���$��\wB+��V1�x/&3��S�B��l���.�ۜT�ݦrL�*PL����ďIW2��_�������u�t[���UQ�
�m��@��b߀����ΰ�(�Ͽ�d}��\��G����K���@�z�o�Y&V�$���Ӭ��s�&P8���P`�_�K-�v�w,�m3�~G�$�,cTB|S*+Ro؍rN� �\F|E�/�z�������/2�默���Ҷ���fT�7I��Isu�����������{-����
]�ӔN���,�[pT/kk�wp�{�(�P~k�V� rEF��n)N^vymܤI�#h8������sh�-�d��<1�yf9O唖9l��I�B��ޔH�>�f"���`��`#�\CBz�3c�c��T���CGzR���F�0�bW�N�h�����`����SZJ����醱����v��j���E|+۽l6��(
�ڦK�ⲎQ �M���q'�Ŷo�J���e�?<���+F��g�X�)�+�����T!׬.d%J̛�࿌���*�٥?z������b?<!>9]��e@.���HB190W�̠{]?��{�F���rZɜN�a�|�x��c��!ٚt�_��_�9��[V�R(����VA�z�b��� =�������xQ�L,����cP
ݛǶo�>U&��^��
JR�i����0�	�Ҿ�_r�AW������˥��}IYI=����XI��yHn+�
�Z�@Wt�jPO�:�}kk0�5��r��<�WE�Y�q
�a��cA�Qp��"g[��w��Y�Ȝ�$D09���GZCQ!1��-h��6���R����Y�"f�Yi�+�3�Ms�Xh�ָ�Q��0���>��΀55�h��r�"�r�~%*\�#�!��t����۱Y
�^� l�6l�#�3q;go`���J6ҡ�Q@/�Amqcy�u�t?ɖ_;K$�p�R�@���?9|&�;�ي�gls�I_�q�4��������Iӎ�W���*HAP�\�&v&���s����%_2n�> -z�|0@0�F��B0(s~��R�AZ����\a��X�(�^q�<�/o��9Xi@'C���c`i����1j�B�����9�{�iD����'���̩�ʵ��������ZL,6����c���>S���T���=�o���Is0V�ћ�&B�������Nb���]q$bF��&
��7�Q�Uob�^���E�A�!�������A���9��]8]��"�h=�{�Đؙ�C�?�<G@��L�Z��	䚜��4I��6��լ�W�9���k�UksF�l�-:-����`���6�s|	�Otܞy��2U���{�\���uWG^׺�!ڻ��֪0\�W .�so�
%��P��Yl��J���C{v+����|G����RRQڦ�ҕ<���"�,��j���x�u-{�*?\���gW���m����;f�'Ɋl�����0�x):迈~�Z:���R&A�``N�0$�`]_���2��+J#WK�̗�{ν>E�N����F�C@N�	y�^��8���.�����Qċ�����\� ��v�7��4yPϏ�S�wA��pW(�q���Z�ֶ�1�T���S�EyrE�QB�$�'z�q��K2��2b�� �aK��$�;0L���iRH��ͭ�xvt˥���q��㩄¡�~�~3��\#==�g���L$������;+��q�)����5Rs Bႌ�W�s���/�aJ��ų�RL����ӛ$>�hf��O|�dbh��>Њ�}_���DV�?�f�d}�}�ɡ������Y����7#����0����Yji�}ֆ��u�XK����^���Ww�v�=�����(ŀ[����S� \�Fވ{�vc�P ��E�M��/�篱��(a��ch,=���'�X-=N�	�2���r�����?��$O0��`N��wU8�B?Mqu���d_.G�db��� �0�}��7�	��;����o����|�9�\�hV��b�[j��W���N}��C[�9o�ʳ�UŎ�b)��?ɒԳ[k�����q�L+��W�j��ȣ&n�[����a$|+|�F@��p՞sX�B|��ERƐ�ρ�@��D>�e��������������ãHGU��*P$1r�ʱ����|P�a�`ƆQ����J���E�N��ce���	.�u�l�=��ot�2ӟ>o�V.�&�_���&�笲�J8ǵTە�B+��í^^(]��E�#CV2��j�&��Dm�Muk~����Ԭ�}�-	J�C�oF�$��e�\�?��M����,�r�/����(]�JH2����
[��kCke��ܮ˕5����	���a��<̧�}�
̃^�j;&�4��ň��tϘ���Q�2��	�M�|�}Y�!�p�k��u�߅�+�6�K����B�j��KY;:�	�ı�x8�˪gfE��Q� O0�˰��l^��93�����;����8��UD���^�Rz=W@�9���$���J@�䢒��'�?z�܀�]����DSw����-�"�Wr��R�zjF2j���T/�T��F�F�̺g�$�9s����HNވq��'9��Bj#�5Y��&�?0�ޯ�[������	�pU
�vG��+�/o,10\ܲK,:0]��e�,a��m�iV��"��̀�� :����gۆjR<���f�vj�A���z�&�9j���]�}.�'NN��Q���f��+�%�H��H���	��ie����(������j��T��>J=
��v�L��z��#CHe�˦������BvHж/�����%ڍ��:
�x����ZqV��G�М��	�_��a
�1.�k����1;j`Ob�c(\OS�����P��(Q�r�sU��)l���*]���F��&�CE'�9�	�����s�Nhƀ$�{��g
{�ў%�bR��qg,���-����%����1�:�B�]߰d0������>�����k���@`�����Fr�8F�g5�[F��W�@�d�
s��E�-���r��ݺ�Л�R{��=)�t�`qy�X�;:�V[�x,�Ά��Xϒ=�`�e�>���+�v��BX[�;�]�j�x���.�~�{��%���k�O ���?[�JXJ�x�r��A��o,�kʌ�+���;�3�hb	)w���6���e�͟���k����ˁ6%BtǙ(t��|��_�ꁚ��l8P�T�D����ʍ9�
�)���S�}���l�+�x��{�u�.�y[AQ��^���`Z�8�Ӛ±Y�j�z�k&��hG�O�],��#C��D�s�޾���*���j�RS���<�Ib�� Cj���&z��ɮ����K��x*
b��A�F���:L{{��(0$�E1JO�x����.��y�`����/�Z�G2�]��)O��^?":����ѭ�r�Mݚwg(�fg�s�P��3���$6��lf:�0O�Hm>�wz���_?4e���^���J���P?S���A
Ȩ0ֈr,ޣv,�k	0+%�.�W�8F2Lz��MIF���&�1����V_�����>0l��{��È<��p�W=Aû�y̇�fT���M�̺XX�`���vT�4�suJg�a�]�͐�����Z�k���{�ql�.�����D��q���-4�ù���Uu��z)�z�ç��K�r���XZ�+��S��4R� ,�
���u3N����]Z�	�[��d��<����V������Ϲ��Zc����X�/ *M��LÏ�%B��w�����S�'�l@�\ ���i6rb�.S_`g\�`稻����M����M��V��'�k�K �P2�?/���?�����������f?|	FVc�4����my����L^�<���$��5�\p�&�ܛ���yB�pp��^ș�������Wݣ� *�v�l3�yl�B����T�x�^���4�Mn����+�Q82;�_k��1T���g����c�wl2B�	�����h��%�4���s��t�ɑZ����:�����t����V�tgP�C�df�.?r����gk��4&��VxK��e�A�\�(��X�=�\��1�<~+�<��=`�(���AQ2����go��, >�`�UZ:2~��b6%�(:-}��"�t�.W�ְϘn�LJl�jf�1�ٷɟ% 5�Z)-�e�h�l���Ջ[a"*����>&����t�#q_�|Ş�B�=7�`�`6���g��1�w!��&��wd�$�+�FR�MK���i���U6%���c�jw�#9Hg��mG7lJF��t�}euh�N�u��I�"��%%�i0N���� [	+���w���|fú��錱�$�k�g4>��_I���za] ���ڈ%.�Jd��I�#�xJ�6L�9�?����卵�|�J���{�U��E�T���+��z��?�`!��~�"�l�;������$?ۆ��GX��LM	9��VA
>VY7�6r��h�1���n��.E���@�}Zp;��sPU�Y���%�@
��J�!C(*�}����w�Gż����Ʉ�:��X4��ж�
`�h�X�b3jTF.۶����L���y�&��|�
��No���H?Z���}C�p��z�B�#o��~����p��y'N]7(��b�}9{Kq L̂����o������A�  ȡ6�H2~:�Q�(��Շ�g������W���pIg�Ǒ-|�W&Ĉ��2(�uF�����(Z���1Ҳ	���L#�����|������gȱij�|�1PZE��o�9u+S����WK�H$v
LPR�gGЇ�v�l�����j|�@�:8�pU�u��rL�?��?_Ƿ��8�;~X�L/�
'	X���]M��T��ce(���
)�8{��S�L5��СӺ�7�%���K��Ǧ�H],�\�H�w�7�s L^��f�֒�t �?�Բ�ε�n_�|�m��s�U�l@WIte�;��L�}�lж�V���"vN6��}�f��N��7	4���(>C-0J�?��J���,��H��w�b�aw���+��Ԕ	&��s}z.z��g=Pr���Fsw�;�?{���p�]�T�8��U=Qcs�q��U���׳�5��yZ��1��#y�A�S�;	���/��gb�rƗ%ʫ�`I'��j�u�g�O	O*�c��3�.������\�0�ߒJvQRܟ<y���f����=���kvZ��R���o��h5��=������,m��?� j@�r?;m[�R��,꿛@}��1��܎ϳ�5�h[m�<��I��>�'}]�_`"����,���d��\k'�H$r�h��w\�w�[E�D�uHw�@�����[,��/���ךO�	�<��>�T�u����^��[�.vٴx9Z�vR�й��LY��6�T�{���\����`\��E�P{4Z�"��MCV��n���x�pח�6�T�#������ڪ��R=�c�6S��Z��$����R�E�X@��@[��-X"���o�HO�Me�«��0?�GQ����gr�^q�F��dgl�X�Q�/��?/j@iM什��(J�.2��gǹ���Yf�Sk�����u�M�8���qqK�h�8�F[f�����Q^�i�k0����������r��n��{{`��|�\�f5�?���;�px>f��g�ɇ��h����	��1sZ��ك<
I���[����#��&u<�r�fz���x��-�(?��6�s)���Tt�)������5}�^j�#�]rV�	��cs'�%8@���r�g��ͽ�bsz`�!��n(/}�Sg՟�J��g�#o���::0���n"��!�*��Q#��J��N��dmt1�����ޭ�so�~�6���%ƨ�4�=	d+{: ���R1E�`��}�������gE�iտ�[�_B��j<`s���	��儩��,��:��U�On���a|��i���(̀�ݕ����h��~ݎ%J�&u/�`]��uQ,��������]�I���=��U��8����C�{�A�����5��םq{��v�}��S��Z���p/���삈��:��� ;�%UT�-I���m�ŶL��%@��D#��Ż�Vgo-�H�+zpϔ�A�	��&z]����)��SY	s)L�"���K��5�iF��M^<3�ԋJ�3�?���S���G�b�$&��_�� � �nW�]ٺ7^B�ҶA��M.�:�����j�2���4���Z�A�`t/��z�K�k�E[��?��5�,�
Fn�_mC�=�|�g�g�WQ,�%Q.G����j�_�F+d�Tԧk���B|��1clgy×���ط��	h�y��'t�d����a[��C����Q���
;��3dd�ӛ �ų�؆��ċְ��н
��<쇗��z�~	�`�\"���~���K;G��o�7�NSB���؟mq�El]ʲ���^�B���X�s�ƶ�\������&��R�X�P�9�V
�6��Vl�(��m,�H����u��>g|�s?�9��_��!	�7�Rh���;H��g0k���	�;a4���f�D=�Jkt��ߏGM~��� �i)ؠ�<�t�ʨy�F�≽)Ţ�N;��a.�_A��)x;$N��';c�\~Q����ǰ�y~����8��07+�ޒ�ݏw��M����uO�Q�-#����:*V�xU��M:�;�.�G`L=<�ڸ+G��<J٨�B��3Jf���rr��(�)W�I��3o�a��4W�7��w�\���v6c�d �۷��W���k��['�=X;l��3!Q�A%�\#q�1�o�t&}���ZU59z_b2N�����!(�_?pA4V�ixY9��q4|A�d�����
��x��?`5�T��Ba���L	-f��Mp��J��2��W֫�.���}��z	�nƬU���Ū;�}��c.�L6ok; ]��@P��EJ�5��z�Q_���GN��j�� �Z<�Oi�����k8�8_��ϸ���.��;�UG/0�dFw������&E!�����̊��g]_��/7�{D���,xmSB�Qߨ�XTï�W������스j(:hCW] ����^}Ycҟ؇������Pܦ��œ��#�GX+Y�����%%)_a�fOQA��8 ^"^�ZR��E`3��X~(���/؈�OB�s��)anQJ6�U�)1A`.%�G�D�e����#����i4D��޴��Wl/��S�'���V����q�*c�K��D�TX�����-]7��I�#q��G��x\]��o�j��`j8���a�M͹���jl�-قm��saM�}�SX�M�S����S%�R�w��E͆�`�l39�"*����)��|��y9(�� ��눥T�ݸp���Xc��҅Ĵ����Z�$�y��(�xY��Mit�����]�KΉ+�t˴�W��X8Q`�5U�}�nK@w���5��G4Q.��#p�i̜�՞7p�,/��gE�a���'�T�Ɔ`?Lh�SL'��mj�VPR�'<�M=��)�\�@,�ͪ@^���C�Ro^�1g�fiW8�A�7�X��QH ^7��S��W>.�b��{Z|�h��Ir?�`�fb�R$�GN%�i��z�6W��ǌeh�_��u�?28	t����7�Ƕ�~UW\��A�aZ���J_MR�+C5W�<2�I��j�l���ů�
��h�N��x�ne���������t������k���=%����i��:�SU ���-��n�z� ���O�Hn�f�\����8HC�Ǥ�)�hMlQڟ����(4�0��.�|�LF3���@纅����tOS�"��\Z��|A$�*Ħ�˞հyt�������1Es4Jn*>;�bʅ�:IѴ���sp�:%a�{�uۭ�ݜH�|-���_�)�ʱ�!UvP>��ĉ���z�)�E��~��XlV�%@�M{���X����T�f��{į�^����ϙ�<a$�����ț:#x�!��E5�����b�̓�O��a��.'2��m/c�ŉ�7)d�:�����ݴcK/��i�
��Ԭs�c�3�M�s�3�}�W.k���b܆�=�L#���\심�]Q���h�[6��TU|�pX�ar���1��<:��#�}�Wڜ����U+��I%�]b����|#Ϙ�i��}��Ck�tr@Z!Gf�϶�N���C�����Q���v#?}:!�d�p#�v�p۹����}&Up�K����ʋ���,> !/����WTtY��_@��$V����%���$_$���M���@�r2�"�>��Xhʵ6]$��������B|�
m'�T�;i����BM�zE� VoQ�^�5)ٓ��XG�<1:����^�U�<m���bY/�*�H<�|��
�	́z�4ټ�"����}����w�֙��5�5d��1�'8��Y�CV�z����7�j��3����s�60Ց"!�^��=��-�Q�J^�}<����;�l�O=�C��o��	���u�^���|B�N_\=y�t��BU��S�X�ia2�5zd�ch�s��]��� �mߌĭa���)o^.��aaby�W��F�H���>ʕ�&̫�W0J�s��e�	�^l�=�{<�ր��d�����]�취:�\1|��ӹ$2���~
��n\wAK��p,@G+��
Ī%��\���%���#�mҞ�&m��E[�������Dv�O�YdXJ)��ݠu'$�}����e��R�˓R���d����sXe?�UE%>�J2D
�J.`�{t�2�Q,���W��^���W�{g�f���� ����z�� nY�C,��a
��_�;�/�+O���qB�B6��V�zp�/������ƈD�k�$�7�Y��Y�����&��%����� л�7P�h_G��!+xEƅ���U�$vIty'���1G�뚫��K�t�e��OI�3z�wdf$2����>DcE���_l�h�u��$��q��׈�Uӣ����ٖ�/zs� u4�y~ycKK����D��"'rx�)�ʙK���\�1�Z���jֲe�4+g��p��x�U����,�G��Ӣ��6�19�ғSh�f/����H�r��x��qE�b�~��-���F��V�A����6