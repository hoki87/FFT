��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#���������l��U�~�׏O����j9�PY���`T���x���s����uí������P��"��b%>�1eτy�<�gܰ�N�Y�	� {��I�ɍL�ݫ�G�R�k��Q�!E	�5E��.��:�͂2��y�m�-�.E��i�����YS�
��@�H�ۼ��nD��Y�l"BU�.TԊ�=�-�����q���Ǹ��j��ԋ����tr�a�ٵ�]�b	��%�ɔe�)rYOjX5;V��R�������M\�	D��ҏ����9c=�Vͼu��Ro�P�Jf�tRvsY��c�"n�XO��	3g���Q���^�Bʹ�7gQ+Г���$�-��t�8�����A���<����l-��*�|d�n����j���E��oּ�O1�m�̭���L�`�<�a�uYV�����>�=�y�m%3��.�������Hj���(�����@�y��_�?�4�}�j�����^m��.�U��$u�&��U��� �.�3�0h��#̻���Ȁ��l�����n�('��t?+p�}J.4ѝt֒��?�7���t(dwF�����j�Ԋ)�ZKnem!Y����tW�E�СȢj?L����z�.O�	�I@�q*����qf߱���k�]�(���7�	�Y
%��ANɉ!e� ��Ab�F���}M8�Sf�G�R���0�Y �,֎?�D~M�ԩ��gJ���y��2��{��@�Yۯ�E���ԏW8���*�����V�6r�i��D�N��s�I��z�b���P�T�T{@��֬a��g��q����Y8%�y���R�޻�e����we�IҲǳ]�ǆ����L5�)h
�3NX]���@��������s͋&��{{\*X�k�M�>l0��+l"�������pC���iuB��L���v���a�g��g���q�2��S��˭;¦�!#����5ۡ�Z�?�E��Y�n��& �L�
�)���9�a���J�^!�Y�����q��<���9��Ć)J��;���w�*:+�s�����	��T�G�곐_���z\D-����BToVD���}�H2��Y�������^�Ì]��H��d�i"�'Rw卬F�R8��&���t-d�V%�n�e��
:r����:��VKύ�@�{gv���ƙ�2�|���i��G�G�F��5%_å�8�q��dO� ���̢\Y�й��1y��
��Em���w��*-���Q!\>	��)�7v��0nU�P��D��D�>�hX�&Dٶ�u_6�"{�Q�6'kI�(7ڟ�B��ʒ��wdh���>,s����ꊸ&�n�8#��>�*m�qӛO�ET��'�kqzvs!#���yݷ�I�'�P3e���Y�g|)���֢����2��\
��)*�u>m�^X����{�pm]��=��K)�K���OT��`����s����m����m��r�OR����]�-J^��J���w��Q�m*A+E��>�J����qAl� ��3��e���A�Y����De!���Hs̨?��nO����d~%���a�0��[J�D���<h�G^���s�w�B�^�wzd��	c���ݿ�������kz�]����-�����Yt�#���+1�x������E�J���%C���� .DGo�ȎBʣ(W5�D�)�&u5/-iV S%V@��!	A���q��m��Yq�l�F�{�ڥ��P1�<]y<�f�Y��<D�l��V�d�|F�s�&W+�0M�G� ���n����5Vk�J�c��M1γ��ˏ�K�_���>�.g	��oz�s�����|�4%i6���E?!��?{	^�a�N��Bz9���I8SK#��]���yFd����XZ�����r1	�n~�'�dv(C��̕��&ٔځ|����X�AO�] YP�!D�F���B�f).�Sz��^%
��������|[L�h7��d8�]@ĉ������ѳ
Xv�Z��<P�M��+�����[��9>���X��[ϰ1��ڕksB�$�Jk_vy�N��$��bh����{��H�/�j5p��nB�f�ۏ���<1�螱Z�%�����z
VE����oXr
�[�(k�v��6�e*�5��3�>t���j�� �f�e4�%������y�E8����芽����C�j�6�b��#Q/G�e�
]{�Պ�6Y3��>o}ޙۡ�ч��f����h*,|6��w�l���#F>�̣��^3w��T�2�pҞ[���{�Ȗ���v`|6�W�!�)�6I 8��p1H� DQ�#� �������Q�R1=!�-�G��9��聠�����+�L6]�J���A���W��L&	B��O^�u|�g���m6i;�Y�mKJ ��m�l��{�ZU0��.�|0G�K|�tj��ElZG)?ݏ��%`d�I�;O����JP������2�	���]C������o��U�~:X�&��p3l�d�}�E��_�>�憤?ZN��V�(+�@�չ#ڽ~����A!�p\J���;��_��b��
'@qf3��H�f)��͡��UR�9���&a�Vv)0̗wdT������u�I�Εb���|�b�B��j__R�kS�G��l�Dn�ஷ�+��H�^nz�	���@��Qd��\�����/��=��,m�pF��o���Q�h�f4�g�y�{�)�M8�~��Y&=���V�Fmf�h�kt���gb>����I������Wm��桐�t_�N����G��>V���<[��vE$?M�s]��@�B������U[Üu�6/���(�(���r�1��� �^�
�{'��qVÆ���p����ů�{�b*�(2P�y�a]��؝�F�Fd���PK�Q����N�
!����q�dUi9H�R��6��4T\��T���p�w3�� yOo~>A��۹�)�c"&�^�s��i*�n�{�N�-<
���ƥ�$���{�g7WW>v!@�#I��xAS�;f#��F/w�~�V��o���]L􁫡�!���;mc�f�kІ^O�E~78vmڠ�Q'�(����x�]�����h��L�b4�dU�s55`@��Q6�k��B�UW� �i�O�u�Ժ��ɑ$�$�9�8q���@qv�6=��-� ��9.M��4*����F��QD4�LZ<t���^�#5��J�nd��p�[���=��#�Ƴ$����P��0��h��(pu���cc����T�ĭ[~��|�x����ٙ5�����2M���s�z��_��>��ݢ�n�O0�W5��1{e��v֧��WUm���ek�h��z�?�K7�v�F�J���)�*h��o2���uF%'�����V��đ���1 =�3�:�-�6��bk~���2o��-#˘LO͜�ҭZe��Uǵ�{��3��7�t����W4
�Jɍs���<����/�[����ML0��W�n�m��1�%c3�)��Z'9�E녯 �_�����w\r���^���:	�B�tr<|>E��GK�$#j�E\�CF��p�&W��qoGв�p(�J,�e~A[T�Gݱ��^��"�R�(��4�H�;̓O,zpQ��b�g���u���2%�6Z�b��\uŃ!��qGJ�G�n���C�� e��r���j�>}�����_�O�No+�*12\}�p��W�F��g��T�.y��lF!�����s��$�[&�z�W�O�`P�	���\9���}e��K�h��K8���1�+�d8��!�~g����l�]���ɝ�Ϥ�Q'�c�+b/���'�.~mdEy?/ P�M$̝�3-Rꉗ��+F�pENC�V���]�UQwK��ɀ)��nC�H-�� )��\��;����5�v����O�~����7t���0�0i3�������Aq���1�V3b ��B��[���� �AD>�QyT�n��}�BaN�0��2�@�t�.���Y:����i\��kF��c��f17�jM�U��#WaMR�*�Bʻ|&�p�����d`�`���$��K������Dd�q,f��V���;�Geľ�	�[2��(.��U�C�V�QQl��Pm��q&��~�s�OtA�::>迬�x�S,���@�Y��D�]���M�*��`�Ռ`��7޼sY;Il�Hi���\7�ʠ���� {��6�|bWM�Fi�8$S	7�N0�y4�8=�,�O>6:qh~z�.Fe�笇�;�� o��VQ�>q���	� %���)2��w�"�%�P��Z�?�ñ2������n{e���z��X�y��˫�oWm5��tg�����/��hB�o�����+m�O������Zj�H�q���(�[�W5G��S����!�'��mMV�-Sܴ��8��]��:��ǆ�7��4Ⱥ+M�U3ȵ�\��3�F��b��Xq2����I�l*��_'1��ީ�ր����f��� xi�z�� H�Ǿ_9{m���O�S�)�g�"�J�2g�U^�GJ����\|��0��c�݄Ú0�.�����X[�����!���KF+i?��+�<D*/��U�w?��R�IQ��_M%�Zѽ������n��̽?�]Zpe��s8o��������~p�,�
��N	~�'q=s>[iK0��.��35`a;0��5��P���b�5 l�� :�`y4n(%ν��S���$�GDf���>�\J�}j�_�j\#�2HS���M[#�c#nH*Bk7i$�P�s #u���,|���;����e�\Ͳ�jӤ�+
��ݠ�����q��3�!1ܶ����6�^���^��9�[	N�=����@�Ar�`�X�D<�qڃ����H�[�"���G\�6�#
����;��P���g;oT���&`#44�-��g�|�SQ]�?]�A��V����I��w��q�p#�%e�s,��y���ïR%����i�H�m��'b�ID��vdA�Mg|�.�#�-<��u#�ǟ7�>��v�/��㌳����e�����9h��X@�X.�f��O�i6�o<��ʗo��}�*�Z��J>h����Rs�d5�V�>�6��ٸ��X���f�ڜ.��#+9b<�.u�&�u�pd$��l�S��=��c0�\W��1⤆p	k��n���I���O-���M���5	r�>���V���q��w^d��﴾����j��UCF�Gf�+��0l��»(�F�5/���!�n7L�Z�`
|Q�Ly�dP�l� ppv��qXK��ޱ屺�+sHA?\W6�~�䐋�7��[��{��=�_�����Wt��÷֪��q#�T���T��j���~��~��Li�!M���HW���(�y(��9in*��8n2IC�BH�9���t�����4WQ�3n*��0ڑv���M���n����|Dy�:�;N3Q'fC(�CAU�֎��t[���*��Zt��+��.�o���q���T%Z@��ֿ�k���CIV��Tw�8-�Ӕ)�iܭ�J�b���Q@�����F��[F[
�����U��IG ���܃��*�
�����ʴ����=����sN��ut��@h�mBs��Fi�t�2�M�(,�#l\"+rʫ]�����R��G$hH�V�q�*�Q�N��6��AE�6�b��Q۷����\Np�,�ǻ�D�Eb���F��"]�m���E��a8q _dg�o3�^aU�5��������a��\v駄�+�D bI���I^=��"��X5���=�N^�aB=&J�$�'DEw�?����'�t��J���;$�V\7/̧z��zh�<��?�z[���(���E��dr��F'>���� r������]L��a�N�룉{�:GOa)�Ѵg�Lo�b��d�@)�"�(�	�`b�e{�[׆�MzXc��$���.���L�T�Ϩ���L*��7�O`ML���A+�����z��Q���f�<�H(����|�mFL9��̨��%`Ɵ4�|�n�F���������n�@8(}�����F����PԾ^5�@[CivHj6Ғ��^��V�d3����t#���!w֔�����=qV�,������B��9� �C<Q��g~ҟ�¦��'�J
��k�~�l%�z-����q��a"��h��K��s%L��01C�b�Lv�����ʢ�~�22����� =F��w-$������eQϼ�M�;���"52��)S)h��@�h��	u￁�"���te| �z�W�6��Tp��9亃V�{CkG���l;�-c�kJ����T`������EVG���s����&Ϫ���nY�k���jr>������t����M�cl��m�'P��(�>؛�듆$���oK�S/2�8�w�L��t���U���[UD+��K�_�"Ir�V�՞��<O�u�z��J�����8@L>�^���gHmtp�g�*,dm�2�H��655m�W�ڌ�������v�j��^9�|����_��ܙ(&�HK\{��Q����*�Ӯg�1Z�0<�7~1�8�b�����z��_�dR�d�����Hő&�[,(���_m��:J+	u���f��k�x4j��� /B6�Ǿ�_��\XD8b<���t^7���&���,|�-B��`��{���͚\
nI�{X��"��j�o�u�y2`iH�nr��uU�{;N��L\�Ӟt���9 �i;emX1]�/�U���鑭��	Y؂S�J^\V��th�HK ��K�Ż�2nm\_�y`45M��W�Y$`��^5�D�[A��#���D���r��StaF�%�O��`���xk�:p t
�`6�#\e�WH����t��~�!KFӸo%�%Ny� ��"��#�}���L���E��f0�����p^�D����d�8������>#����Fxf��p���'����٢���k�<SQT�$�c�����1������s&&��g�ŧ�=�3���x�B(�"�fc�>J���la�����5|���� ,󬲱lhPU<�ӈ��E��<JУ�u7���`��
cI�����D���������F|��)�0|"�ԕ������p�\2�:)��b�3����ܒ�(���-�u�=d���2ˊֱй��){��������E�B�n����ܤ���MfY��ݐ�06zq����\�t"����'�cdI��	;w��~Ì�/_�^<��6y��5ǌ�����	� (�E�)��_�@ţ����@�M��t�]�;T��+���q�_9���nYt{ԝ󋽢�s=D���?��g�VP��f����ve�!
Y��o"N�
Ysӡ�!����s�7��8��̂X|y5".����Mc�{��K��	#�!?=~���4�b:�d�螲鮣�,�NmW���جO=I]�%F7�%kq�Fj���Է�(,O�uyl�-�.�SvY�ֺt�y;��Zs�P�?$I��Tdn�����\\˽���W��bl��ϴ�?��9��΅Ӡ��+�NƷz�y��(��y��z�k�QMM�l�hv���]݀��>ǹ?%���i�rLU�a��9�<L{�!Պߘ�ML5b����x�0����?�}Bo��p��D�_�w͝Co���HM��}e;?p���'�d��#�3/�O�J�l��C�P��F�$a�,l4e�^ 
C廙��7F{jK�k�W��h��������/�s��zY��g���j��Q��j�j���;Q�ɂ����jf���E��\��q6��Au���sbS�@E���5���c�2_��$a8�0|�ʡa�� �B�����0��/)�{�(!����uE�~�M絈�^�z�#W]���>��sɛ$�k����z���Ӛ���0���`\���ԏ��L��H��$C�{�*)'C!�g?����wI�#JY�����x>�}jf�x����bċ�6,��nM@0���J����&OY	��ַ��䲊���������x���4��rҷ���ŖFQ�٤��6��H��N�\!��,�����H?�$��s�]�:<0Ϻ���/��5\Z��}	�Y�&��'Q<qU�O�^�)NKC�4����Z�O�)^�i"x|.Hm��XB�p\�d�N:�/�+�Q��Ւ�D�F��c�8�0��r�?V�� �̅�6� FWK�SS�e����Vmt��ߡ�<n}��<Q�+i�R=����!z9תũ�b��&�+�`�1痫_�Opj"�r��Y�ә#�[>n����$"�?�GӼ�/YtЍO�r/�:�%j����n�X��r���t����0�\i�N~��"8��1��M�ߣ;��n?�������䠤�6 �#�?=(�H�r�h�O- �(Pr�X�-�;�II�p�&]�~��2x��KvR@����9��kWDMJnc��������PE�� {�s����ع�3OT�Jȉ��5?R�z�s<�3-�TAT�P�r܄`^	�K���a�ss����$���z��#��/�ǰ�U
�⟘]&�{:f)��C��6��@����i�W#j�������@��#�L����U/��`�C�of�V�Ue���Ё��_++��c˺�4X9&U�d�Tx��*���Z�LpR��
� ��Gk����Ǔ��fܽ\a9��ے@}&��Ȇ3ݛ��2���Hď"�G�3��'��>�8�7�1e���v���a�G�1�5�{O��(�Lir��ī:��bu��B�K-�ܝ_7�Q~t�c�����y�+�,t��C�W+�㶙�R�a
��R�:V����M�l�q�L��������&��Ċ)K��k�n=���e�A	�g��m��D��@���%�SbL���W�\1�������Xo�)�a0TBӍq��$"�u{M @OŅB0����`B�Өvm�Hp�����F�{7�:�Y�@��{s��~n�h����]FϱZD���1�or�c�xn�<�:�w���|���|M\�-N�X�b�'�X���na���yp;=�!��¯�6ޘ��g"����ؐ����&���՞[:(!Em���<�N�|�3I��1(۸�P���fc��U�#I�R���Vǒ,(gG|A�T��8��K��mW��^��nDu/G}>1���K�8}���	#T˯==:씡K��uA�!����)�!ݵ�ޫv����Y �}��^@1A�MGq-����j*�����M�v�"�1{�e�O^q�u��+B�߭�?�kfN�˝GY����Zc�wøȘ��Ҍɉ���gm
qA��%	���|�\���i�|�9�(��)�k�?�7x�zV\U�#�oK�;��B�l�,wٖ��z=VY�;����S4힚��y�gd ˩��y��=>O-y;Ls��_~�Bn;'E���E��RU�+��I���B6��tO�4Rȷ�.izQ�^�8�2�yNk��CC>+L,��g�oU��m��K;8�"R�4.�	�Y�����J*����Y���� /��V�$VA�p@�V_��>���Q/{��CbPk@(a��=�R������?�8���цd$FG��m�$��VZ�U (� J6��c��!UM�iӰID���_��|��ߝ\P�v���v��A-_�!G,{��uTn�,�N&���l(&Dt�]��i��F��ۍs�{�@�\-�e��k���+~w}���@ϱ����_�Vտ�Y�/.�t�J1ch%^d�!������}i�U��M!fd��뉍���pik�zy�A�L��D�����Q���M@u�v�-d�Yb�k�j.���3f��5�}��5����q>����%�0�/�E���Y���/N��5B�O��L-
�s���Yq7���M�S˨���'��\ug�#�=��ds��"��nŵo�?IT[�ͿаD�N���x~����us\��O���D�{C������X�^d�A�-e����Yp�"���5d�!���6�|���m^G����+q��R^В��Y�w(��"�\"$��Yw��k�E�$ .�?A
���l5N'�%�7���uk�ffk������Ϸ�|�
U�l��0�In��m��{-���]#9|\� *�%��ޒ-����~��U��O,#3�"[�V^�O��i��$��2_(/wi,�A�~�T3!:.�c^�*�� G���g�x����L�[��Ϗv��� q�0�f?^��`#(���v���^v'R	�It�X��
{�.d�E<�m�&Jf'����S�[գ]��|W�:QG���\�m���
r����au��O�!h�R�EX�~�$�(i�xX������tT�M��&|��;��qO|�w5�n�m(�W"j�!5lw����E�ՠ<�fɚv�B=;&%�����H�B��RF����3U��BZ��ocDr2iz"�1-"lĐ4��t��m�6	<�f���w�'45[)�?f|�z�t�N�}���a�5���9Ou7HӺ��w@C��4e�<�y�Y��(ΠZq�L�?�5���
�x;L�<���6:��[־��DdW�.��zm��@6�<rdv��0��������Aw��{���x���4]]��,���.�KyK̴M�f�>٣���y�S->�y[(!7Q�q� yau�Y�5�uA���|�LO�Z,����֟U�;�Dp�����T6��������@�\�!*� �lQ��t����Ur⫔OI*�S��)�D9QY�k�n�b�%~�&h��d��G���C8p#����ɘc��sk
d����m���/M���*�7���.Ú<�e�3QW�(�CH��BA�v�x��܀h-<�z够/�L�Ͷ-���)<W͹'���?��m�G$�(	�9�t�jqO��>0�
���S݈IU�6CbTt)� �P��}~U*V� u���G��Z��}v���������^ec��;n���У�p�I�\�e����瘪����	X�x��>��J\��UOv��eN2?K����&����M��"���3���Te��bw�;����~������{aJtR.��OY>y�;�Z��$&�R\�D&F�e�+�ٖT '�3&8�r��:P��ѐKqS�~��{R�� �[U�������=B��\'_@|��!T7�eS4��\<��^l�}�6_
v��{�%$AҸ�bߵ6�.�j\Ϧe_8� ��y�`~����w��8�Q�Ԙ}����4�f�jۭ�z��������Z�ԃ�����s�s@�=�wN1� �Yִ�������j;\��-�J������XB����7�:�(��1�v)��C�.%�����M_H��%K>|-���V�Lޕ���SvH��i�>"�yK�d4.�lD�h^]�"��YѬ6���8��`d���-S�-��e�`-���^�êZBk?����QZ��F��q�{���П�t~N����7��Ƣ�>%�Y/$��&��d��g��	�D b��>�>n9j�ݍ߈��_���?��c�tI���u�_�)PSu��!�����]B)�l��ސ�?�r�O%}�$
�?�q��CV��������PF��kҭ#�q=/<�1d������a��`>]t�!Uc��80R���qd�b��n���g�K�l�9�:3���psAˈ	��.��d��B_hD
p�9|�� �~a�ѻ��zKBG�P(]���~N�5m+�����!6�
�W���ĕ8�BG���z��὞��,�L�{���FU6�egsN��N����g�����o�'0OL�ȥ	��������Aa�\��߰�V��o�/��������@� ����|��K�s��ی��J/��z@�3��|(��x'�x@I���K���%������g���g���6>J��Eo2 �v��i:��B�cc�eLڌ��!�i��x�g�fw1k~޷���<a�VR_�H�%��c	����I6�"R��9�>��^ǣ���5h���FL='��������y�\�,J�&�kZ^#@� �k�wa �6L�H����R-?�f-��������鈸�I߮�&�o�����M��0��I�e���W���F�K �̭���~��b2�����)��(Z#�{"��1�1��]��AD�+��J�e?�a(�L!L~]ʒ�,n:�LF;��s�7X�p�Ա���@jK�rZB�:����3�R�s:��BT�� ������֝j�9E%�<���8Le��;�˫$�(ӿ�R�u��l��A�X�����\fߤ(d�|�I���]Ո7N@����Fh�q�������*�H�Zꇑ�wG�H
��2+��wX�uo[�ƨ��c����S�C�Na�tyN{�{��-�Z�՜LE�*ɜ�R������p�B�I9 ��m=^z��֝��˗&���;'���g�=�w¶`�н�(X�+�fS|�xo�Y��EN۞������^�o&7�����W�7B����ѓU :6%�cQ�K_�Yi0���
�V�O�{48�K獻��v����e����f?�/���a�Cf�Q�s�b���: ?��.��e�_���ye�W��w��33�$�r��P�q����a��y~Άc�7��R=U�� ҄�_$gs���1�[j&�������zL��i[���R����Q>l}<��fX��ݝ�E9�{��)���#Χ�"�+C����[\�e� �G�(��\�8��Io�!�Ci	��F,;��78�3�����oV��g��{#�f�2	���2�%WޑU�����V�V�^HUȈ�?Z��6�5ہee��&5$k.�I�aV
R��܊�дG"l�c9��i���e���$$�iA3U���1�d��A?Sˠ���Jvc�:��Tߍ��u��G;�C�[XIJ�˜�F��zd��C g��0�Y�ʚE$�������2��7�/������N���q�u�
���ڛ7.�݅�oHZf�������]W�uo�>�<��k�5"&��f��<I��&P��+�e�.�&�������d�|n�:Ӎ�3R��5S��R�Aʛ�76�����Nx��p>	�1�K*��e�"ŮΗ̵F�]���%��GD��m�����/��:�ELm���Ϻ�%�C��L���2�$+���;*��p�R;Os�Wއ�)4���l6��~b��再�Y'�^���J���!4F�QYׂ(��H�� �}-��1w�Fv��Pt�Ȥ&=6�9h���i�-��O1���S_�rn�qy�ȳo����������F�!Rp���x�?�x��r�C>p����dQs@O����)<��a�{Y������bF��b�!nǵ���{��G��J͉_ 	)<K��zv�͍^������5�h�[ҟ�ԅW����C�ɟ)hj^���� ���xҡSL@�Y�@̫Hя��� mtH���?�.4����WⲬ�����85���\�e	C������`���ki�6F���5�*nA�&�TՀ�A���,YEq�5��6��1�c���4�6����!J��(��� �׀��9��PB3~���� hF�
��18�.�s����F_��;Q�e���8�A}���`j<ߧ����;�5@fJ���$8��'�*d�����~�5��`�sf?��>�����E;ۦ����̲�@�JU��<���e��g�9F�F8��U��� Θ���[��6Sƃ+U�l��@Ӛ�i�6e�By�j�3���í&�)��ׄ8c�v�"_�t�j��-z�O`���<!T|��812Ғu�_���c�k�n�-��Y9��1p|�5L��rz����m� DR��� p�<ڮ���vB����C|&@R𦔔5��T��5uj�0B�ډ�<���Y�������=�сBj��t��[��;*/���k������0�.b�f2��D�qKk3x���S���fN8��G�Yr�Z�4$�e�nW]��8���dٖ�O3}<��R|)���Mꋞ5T*��]g��s(�p����� +,��[C���i/�LP1�ԘG���A��/p����L�����vvh܍�c���9�"�m��s0��	��)p����q������y)�𭍻?Z��u���-��:�[�oKI���C\�@���M�c&{�NVJ'"�]�]���9q4�pT��%g�>F�nv��d�wM�jܜ��\���V�B%�"&�+��-�f0��2Y=��ܴ@�_��<���ԟ������8�S���ț[[M0j83�f��Î�[F:'i�RkW�����^{]3�;��nL�|~�Bo#|�֣*�Z=qｬ�^�y�D�}�E�������ڦO&X��	�ZHg:�G��.�Ǯ����� \o�q#�y\ �ͪ�Ȳ�,�^�*�/�7+��_�Ӳi��>V�5Y̤Ӣ��[��������2�~���8'�31��?Qi`wk�|ڕ�F��3�'$s����юS�;�E}��1"~��r�D/Ho4R��5i���G!�z9��kz�K��G�O�st'�q �³��uv�<���-|�Ն�W��wlҼS��͊��;����&B~���0V�"6&�c�w'ݗc��@�&��S�a�S��0Z����_�Sd�5hiY�d9%JN_�����WW���yF��6ZJ�{�U��q�6&�2��'zq�g���}Ԕ���W�O>�G�%����G�v�͢4�1M��Dxr'!�'9�\�N�4�~��(Q%`sO1ٙ��?[Tl�5@ ��/6]����W>.w��������A0���f�pNwM4oг��j,�yBM����S���A�����>>�؛��]	�Q:��!U�����ʲ6P�i����`�����0ՙ�������_6�)�����;��!�S�����Y~<>@ͯG�Lԃ�ۈH�Yžôj(�����D�i���[*{nGI:"�]�kX��!H& �cZ_o]�zw�"���5�(x��/- �֋���ݴ�� ��ft�-���� �cڛ�#�s��Q|p�Xy���B]
�P�th�a�%3S��%M|�9�:����
���z`D T�4�l�૳ER�<��Z��~�����lBsz�Ԃu�S�͖2��=��T��M�z��]�e�/����-���f���{�����H��wFk �U8�rT �_|��2&pI��l�Xc�a�s�Σ�S`���)-[\u����_���y���q�s���٧	 z��	���\���K�՜B��}�y}���,�Xf�+��0�v����ڮٖ�.7���<��LQ����!
U~�X���c-x��C'D�U�'�4P�Jп����h�|쮷y#r˷�Ӓ�؟�z"�x��\E�^|ʞEd�;M"j$S7l�G'��Y���a�>z�QS�Q���Ո�%���0�Y23���8څ�.���hh��1��]�x>�Q':��|��СUq1`	�F��/!���_)HC~��m]X���i�B��fIŨ����D4����(�dC�73��bQTza�"�Bg�o��s�=a`��ʋ΂l� ����)8��b��:+�v��F8����*�Y]j�"Xd.�\Y$��B�`2w ���,RS�>J�6WL?@X��D��eJ�ƈFk �Z�=��0w6�_��|7��ئx�;Ӭ�9���[�k�������iY��p�'������]����_��4ԍ�� ~�
�
����
�y�+�nO[D��h���q'�k
��D���<���M�m���%<Y��"?h�V_>�ay���Ȥ(�L6�Y��L%]꿙�2�NR�B�����$!��GFbx��y*=��r�CkB��Q��`l�4�`l��&����L!)�th��������ڒv�Kn�W�^��Zǅ�Bd��Y�5��u�gaT��qV�,�Q@��Q������[���*{y�R%�m��*~�RF�m#�'A^Tu؄�ԉo=1�_8��i�ٳ��u�,�P+��O�߿�6;R�m�J Yb���T�4ۀ��6+�7���cYӥM� s�<��#cQ��+���N�ڑ��]ZI�����9�#�pi>U�n���(�]�,&o;�-�_�HQ�����k��Rog<��=?�92VM���``�;kb�I��r� qN��ƨ�y㩫> Od��(��p_���7�G�ްn�!;�B%v*��[��sAL��Aö�� Ǻ�A���u�*y'�������G��n���0N�Ԯ ������z��'Gu����J����>�"6Lb����>�Wע��i^���~�����G>�7�rTԱZbyPy�q� �֥o*m��wT��-��p_�eKJ��t,*@e2�V���)&�]4OVLƵ��`�c%%r����r�4����~�yۻj�Vơϖr`e7GG��ₕ�Vv8ނQ�w�Ha!�����f���Tꯍ���c[��X3̣y����/ڐ�o�:H� tO�!V]w�Ps�G#	����u���kL�]�6���I���?dm�KՔb�S���X̣?�ƺ=����\Ճ��	�y3#�*��Ѽg�������W�"����ia����?���JvYJ"^tKJ��+��3]�dkA�o+k~���z�PLW�<�<�0?�l4��N7�����~�����*����gw����Ƥt�1���3���$��'�0�� ��������5Ѥj��$.�L�mF�JM��2/�vY��gH������#ط>D�#6پ�Yi^	�#7��������xj���$�E/�m뾒�R�g���ۭG����_�R��� ���_ ���x�O�=��`o���ԈD=�ۛRD�BT8�I�x}A$�GZ�q\AQ#!9[B����l�ӎ�z`����q�=*�0�\�Kc\�0y6�����[[+�[v�.��t�n�
F�/��b򐘌�E#� N�8{Y<�r�h��an<m����� M-'��C����2��0Lֻ��!�.<���$��^%�Q6Rh����)�g]׆�Am�,6Kū|�j���ƍr��ez:��k��'a�*Z~��uBf�3`���bq}�@�7������^�qgh���j>g�k��C#꫕hvJ���Y��F1	�و!�A��A���3��	udyq�3�.��z��&������2��x��h���_̧����7�8�{�,�*S���M��]9�ߧj>l��("e��~��&�+��k}�E���Ց�2�E��U��ʤ�`A�������ڱ�666}�
�v|��"#3o�#R��#8ar~ͅ�"�f�c����-�M��@8k�H���C����)��W��!�V*Ze���B�4����?d�(�+%��?��훴�FJ%G��!��[�M���+,���i�܏{�	~W��.6��$�vӇ����w���`W/N��l2�->V� �o� I.�����R�����L��NV� ��<�&K��8��&g~] ����Q]�W�EkT�W��o�XŅ"���f�u��k�.g���U�X���|��tO����f=m�>w�5�=��pt�+ZVem�R�ͯ��^�J*��˩���@�kV��]�/��pݽ�;����M.���_rmqr�:�o�i����㗥�v�%�dNq��h:
5�o%����T�"���5<�]n��\�K��n�;���;�HS9jn��>��
��lq�_�0Bl�+(�ܡg}]�g���Ah%��6�DC%i�;���e74�S�����׆�@��Y|C���c��ن֟e9e7�9�b��c����z�\Ž���-'�H*�˘���4�~���8�k�a'�\|S�a�>��	�6���S����X���"x�Lb��g�,=�G���z�5hMn�X�����0�	����>7'��N�}P����ۨu�N��,���*�q
�fu޶��7������V��N���y�|+9�l;ނ��b��*-&��V{��'^f�O��|��#9��(t�{O���yi��d�I�R_�℣%0�ΧypR��kg�7��|�k$��+O3�!,�*��@������~$�j�|@c�Y����PC�Zb��6,���Xn��v���O�x�T���O�(m*��JO�c(j'���U������w��i�kA;У�#�C���P�	BF�|��C�E��s�� �S��s����yЍ}��.W�^]Ζ>������׌pA���u/y������oݙ���*�94��UlI����H��ىeFo	�l�c�0�y�~�w�{ɦOu*>nod�tq�f��>���w�6&���ǎ�W�m]�{:��JiU��O\��oQ�}��;Os��w�ߝ���ibz����NQ�����⒑�:a5�q,5ͣ
�"�{��!� �z��#[�c>�;n���;���#�+�X]]tE��h<�в���X[�.ٹ�lxZ�F��Ey:-R�-�K��[�4՝�Ι��~ uVp����~�Ý�hH��͠JC���!�+㸭4���`G��z�/l]�5��A1[q���󏣽�7��J B�o&ֻW�(Pc_RJ4(}T<y&B'D����i7��0�����9�Gم9��+�:��M (��(BwbG�ƕ8 �ѡ���}R��Y�Cvg����}��)z3\���ӟm��q��+"��z�҃gH$��l<�S�w؏.�?��S�Y�*J�!͌g?@�HeD�zhƮ��}��dqSɅ��&�<N�Um#�]b_&�9��ahM����lGzHZU�V�C�c�-�D��d��E�Z��D�o�ӹ�~�eqk��$�
>����=w~YfK��1�&�[�w�]���,7Ff)7yw9O� �ݧ\�R��UN����}ϕ�D�~�-�m��J��w\��&!�������a�o0�7"��a����>"����u�j-R�9.a��@qg6�o�GO�*��ySi�_�'4����D!�`5UhU�#�u���-��9Y��7Y]9�:.@A���fS��A�}@j��;��PNR&�`O�=z�-Lp��^q��G��_,�#�v� �$�$yw�����f�=�n��Jӗ���[�8�OV����a��im�ZQ���ER�j���)JV�����N*�U,�ٌ����+��p���O�[���l��on��ׂ������v�
�k�H69m�w%��//~m����|�� �R����Sl�A&[�Wn���˚e�}�54-C<����0#ݧ�`��*KUox��#�8�5WrmJ��m�0H���*���Tz�!����v�WS]|�1�� ���Љ %� �ʷ���Y��@Pz����;��}��+��̏1�!;���ʈ���	���G�\�Q0L��N�]��1��s�L6�D�ce�<c
��d�/z��<�����ք�K�Pa\���k8�-O9�X�#�>�C��r����W��݋�"Ll���FVCiTy�[�͊׶ʰp;*����k�9�$��[V[�#Ď����{� J���H;Zy�F��%�ώ�U]��I�&$��R#��̄������[�lH�����>&xO������y����Z$s��(S�%٨sg-y���cd�����n�!����vX<�p26pr߭�˩I>@3n���DY����G��<��n@[�C�sA�8o>i��಑�{i���"��C�-�秘�E��{T6K� ���>��>��)$��`m��K�d�`Ml��4�4{N� !���W�����u\`[������@:f�x����Y��8��� P�$w�u�#m�o�W>�s8�SbG!��x�@\$C~-����*�	]Ĕf�Z#�������Yy�� �Ă䳖��Qf�ơ]�3�k5\�o���-��i��oty:�L�<#�s�Se �ڟ:E�<��7��=óq%l |�A6��,���u���}�J��?����z���)�%��u����/]�45��4����@񣍧`�	��ErX{�q��ԭǴ����IV3*�-��(��GT~־/�X7�*>���mkrvÙ`˷Ktn5���#2���M�G���%U3�5v;�F�:oN���Kcc��a�m8����mڤ�?�*���,V�P_ɐ���BaC�K#�by�sMf/r�:�&�imQC����c��<3��*���Benӗ~�3�stj7"6�O�����/��>��輇U�x	dJ���N���	��E@�G�)�<�T(���@cI3I�-��Q�$"H�Rb���â���T��[4�L'�Ƕ����o��:¼K@K��E�����l�gY# ʿ!��p�� =��^1�I��{6��J
ȣł�{���>4y�p��G��:��g�n��*<�p�6���a����݋~��J��-�<n�M�)J1�O�$�x��sT��:v���;�Sy�y�ԩ��p9��ɱ��jBe��+�=��L(���'��QO�S�^@�M���aׁ��!��~y�5����2�ٻ�TW�Iq�m@��%_{����וҵ�I���Dd�әƲ�.�)r�d�V��yT����~�z*{w��ٲ\�E���]�/�J7|j�+�������?��cX����mv /pM�nw��u���؊�|����h�BA�vt-aC��GK��W��ƭ��}��t��!��g�;���;��}�|@��b{yP�����	Qº1���û�z%���Wb��5
|�����p�^�O0����HJB �uhR���Ϫ��O�%WC��S��qZ4ҝՋ��#V�Xڍ��J�٘T{����=�l�"����0˩S�DAcA\<��ug��	�ͮq�/a���
xu�������}��qw!�������qf)!��E��*�
9P� �Q �f^����mlY��TOrڞ���S�2���̼����)F2�o�y�S��b��>p�5M#���D�4U�]�;]�Ԑ(��������J�#HH�rv�Pp� �&�}7���O,��(֢A��,�ȅ��M���<����-��?��5iV]p^���+���p��i��=f���� T,�^p\1��T�<�CK')�5q���tq,�lh?�֒�Lţ��bn�c}�:��(�X���U��6�n���fQ���ɾf�D��d����\�o�S���'|�.�!���ӎø�Y+�j����b��+PA���	�g��D�|3g9��ݔ��{���DCT!=R��\�#�[��MXU_��݊}>�-�̮,�@�]�h�0�8t7�8��@��%�A���XO[���|�·�Mx���p
<���~9��u)�IFk[�UN
���qհ��]��o����#�kH�nݥհp���;��K �&���ӄ�t�,a�1�.'�p��m�x� <�L�&��PP�����L��.;�}ũq����p;����m�2�^�2E���ԟ,P[�g'1���� U�hx�-n~�l�-�T'5h�9=.2���6�98T"�G���t-ѵ2��[��*@�Q�Έz�G?fऽ�g�E�.�)k�i�ix]���5��J�gO�c�"�3q�RT�I�+j-LO� "�P�2��z��q�#��x����t�V��e"���������$�#����b�{�H���n���[0dF��V1Į���$��;6H�2�:���>���(��7���̇x��� L�d-�S��ɇ�l����e��hr�Z�6��C΃y

��Nh$/r�.2�L���1�B��*�z곒�~8����L]���W��[�C
>�wf/"�_4G˺PI���4�w�(B�\�g����tUe�4������H�_��}�����*�=�.n�R�FS��1g֫����6׿. b�k�ɏa�B��1+$3q�^;JU���������y�؀��8��8H%G��"�R+;��� 6�iKݡ>+�	���6@Z_���2�ÈD`�gR��M[ E|�U�{��Ͳa3�f�E��كP�%x�ڊT�{oY�71�$Asv���b�N"��uIq���x��7z!at�ܖ���LZ�o���_Hu/��	�T~�s���]�~���6��VtL�B�!�D5ۆ�Z̈2D��O���<5/�L4N\�0�~9+:Zr�bq?���:��O�[ң{��}���B(?���jG�ĕ}��\kLf�����ï�(-?=37-�y��=��Zw�d.��3�v�x�ﲌm��Y�n�VD�?
�e1��������[)�ά���rj�yy�[���C�\�U�7\��+KVBOuΈ�a��
/a=�ݙ�����=���vw���5\�b@_kg�?dovwL<R��Ȧ����}7Q�C����4��Vp�S�+o�n�J�Y�=��{dX8���9F�a��r���25�T�B{a�����u�h�H"]6�[���+���� ������%Tˣ�e�,I��*d\�b�J^<Y�nP�	���R�o8��G��R��4��h�q� ��{l����S�#J��\�Z��R�[����qCst�����Sg ���h�Da�����\����e8uS��6�C��	��������A�֩k����{N ���~�A`�9{7�<�B�,��Y�Bk(o�����Q:7����0��?�W���0���(�Ț�ZǺzI5q�^�o�f�ѐz��Aʮ����:�8"p��|1��)_2�{��m���'����fT[{D�Щ�Ի��,��4��.�mQ���5��[���R�%W�˱ӳ*=$ι4CM��W�p��2�e�F�#����w���	�3�s�nc���،�1T��V��>�b�c�xfd���$iԾB\cɕx$ �C���[ƅ���[�4��.��K��mP.��.{J9+0�����^}�,�v�����r���:����o��
h�x�E��� !+��
�T�����cR�I
��F�֌�y�ފ#{
r����!8'��\$�m	����v�DT�G�!�}<M�]_�X��K F<ߜ��{��9�c���|�.��*��/i�N��\��̝��QR��$�d��J�w����܌C�0��,�{8�Y���n��$fP����'�~�lŔ4L8�;�d���3�,�3u�.���rT�e��\(ZۯI����ѿM�s��3� ��D��X0���F����껗F��)��mB�#�����J�K��\,���"yq�!���4'U~ڨ���r���6M$g���w�Bxq���E�[��-j,=7q��X�\��R|���z���vrڭ�"�n��
��Y��7��[�������Z���h%�o�jZ�7�ofr���`�I�l��0���EOc��Kc����N���q�?�-.q+�Cb��p��nO�("���� ce*���]�m˃��_�$�0�w��G/���y��f��+e#�q:�Ń�e;A�+F�o����<r�� `,��N�3x��)F-���v�~��HΊժO�^��>�	z8�a��g	�o�����:�J���*�N� YC+v��5���j��3��֥kP?�T�1J �՘��I%���t��Wݮ�D��(����T�Ư_JN�KO���r�Zq���Ro���`������Rf77U���]ٕ��ү���>d�BeP*I �l�u0JtYAL������½�뱴�m;�����ƣ�K���S֖�~C�ᛚ�SS�zϩ���1.��~�U����1�i�6�z�P�C2���d�������~G'4�<��F�۔DNyÜ�X�Ӧ'�_5�I=�D��7��5!�c/�d�A,���w�]|���^����Z�=iF�����6ܫ�t���4�v �
忤^3�P ������z�C���;+'3GT�f������?�e�u���Y4�B. K�Bʱ�˘$�D�����o�kn��%|��(��QܩS��f���2��n����k��z�;N���`�����7�4��4�ShX�9�O��T("�dF�q�2΀|p�rf���z��8�)Y�hUV�pE�(#���J�W���JB��aHFiO�#���]�Ɠ�&k�"5�Q'Jm�@�؍<)G�w��\2��Ŧd������"2N��� ploq��g(e�����*vg>����1�y�R��l�K�⌲,%v�3��3m�RY@���z]�}J:��44��ū�RCP�����^�&8�W��9f�@w�,�E]�`����l�����^�v��h\ъ� �8N��u]+��f<V��GCdP���9F.w[S������c��Y�U_<�}�ׇ�����<T�Ν�e�O5���d3]EL��[d���%6�B�1� ���a^;j���^��៊��J��Ri�~���y��ǫ�&�̇�|�ڷ�T�X5�>�e��"�d��4�D����G��o�,�%WbG����J�hM2��h7���w|��QN�"
�#s�`��D��7��IN�i�A35=P�;��h>� .��}��Ǻ��_�3"��L�x���N.��g��_m���v2u��7}ip��э�����S�D@`pq�R'��0\�%�Ѭn�}����э(�Э�Ed��X�l��~t���E�]p4ٗ���X�"�!7�h��S~� E$�&�s<>K�ư����d�����p���J���~W�8ҝ&��$�{S�V�-ב(�0�j�,�����O����n��uy�F2�i>&����햠��C���r�3�h����^�Dx�f=j$��TNaH������pDH��i�n��1�s�3�T��2�R`���W�`dd�pSHWl`�X�3��II���Ӧ� ��;>��U�ݐ���)>�R�4�pS�xĻ4�Z�D�*I�-���]7y�����֠��!K��rH�d�'�PĞr���/�I,˯��#�2�����"�GL�"V�u��7O����$�{CO��ɑ�;�b����!�0�.�l��� F����z�@���]"w��o<�����)�s�ۅ�\�7W��o��.��g��9����1�D}e_E���k:�)�-�<(��B���Eo:F�ƭ���;���ʋ�PTw#�:�6:)_��l8�����AB�i���Ϩ�!tڳ���,x5�x����U,Taǌ�	>9�g27*����I �P׎�w�%�ȍ���L�7'���_!�Vk;|\�'&tw�!�b}D���S+g���rJ��'�%0|A�
N���yΜ>��qV��0MZ�*ڊ��pC��.�؋��'twVT���O��$�K�jcټN'쟢�^�D�}p��YC]��T��9.��*;�.(и���މ��'�5L�s[�M3��V^�vW!�鿍>����}�;.���>�ƿX�yF2W�~0&@��Ψ�V���߳q�f��{k";�.�}+$r,�5���(7���=�'�X��Ee#WfԢ����,^�C�=�Su1 �R���i�b%.E��6�\m/��Í:�|���p�$D�Lm�x�F��ͣ|By����Ɋ>w�	��l]��m'��/{��eD�z��t����"v1z[���"��*Q����xe=������P�,揔�4�es��֙h���^P���?����iP�i�f񜍡���f3��� �T�&�+r�\�ٰ�=Dl�.�ȩ�1w八5���I���'9�F���Ǎ�|��R�(�������w�ʨ���Hjc�;�3���[��4��w}���h��<j��F��$�\����q���d�٬�����ޡ��	�j�g��bk(\Eo�e9.):%�~a��k��[�©H%�<Y9+��{�&�u	��Ԇ�ɂ�@.�(y�V z�1��y ���e�\	DP:~ Wp�8"�w��P%7�$����I��9O�s^[ͱki"h���g[�
�v��ƜF�<ƈ{�R
.{}����Q�<�r����nh�tC�F��
�ւG��)\a�ʾ�4<>tDGlf%M�T����a>�IX�o�!䮸�>��	��췔�{y�MU��:k>?�*��3@��ʞ�u��A����T�/��چ�1nE���Q����e� ϥ>�pKwl��^�Ktv�ѳ� p����:� D`���=�%��n�ΐ��T�FA��ʆ\�%��-��3��c����Vy���s6���{�IUpb����s?�7亼�.��S��=��`���a��*i0��z�L� ׀�ޟ�@���b
b�Kg\W5n)���IBaevp�������v�ѝ��w�r� �>H��� !P!Q9ӕ���?��w�%��w0��$p��1(�ĢK��M���ө���~�M�9��c�r�'y��^���Rn0b��X.����-�U�Q_�(.5qmI��g�0������qPL�Ϻ��8���aƨ)��_�sA�.�s��!��M�>yQVbT�6]tB� ��Wk$SX\_�5D� ����K�Qj��l[��Y�H�������e�1M֘/���:��4�$��%B&8��[v��@e��4ރ��MD�����e�YS���4?#��B�M-<�O��Q#2�u��'��|�:cބ���J��0�/�ANH��~}i��(�iE�C�@�ݤ6�����p)�eW}��8�t:x����5�m���R&?^h�EϽ��C��z�S�)�+�{U�3�\4yWzh�t�}�+��et�횹c�Ŭ�f���m�^$���F$ 0�vji���0~] ��ÉS�h����w�8@w&�rTl<C"{�l/������Rw,ωP�|�#9��7����e`-���zL��oUc���m)��Z������u�HCi�nX�ͽ��6��DRK�^�q�4-Կ�d�_u�}%cYeU���U��	y�U�ň߸�t{lF�:NC��n�<_�{JJ�Vg��-�������f}���(X"��	�z���o[C�I���la��!�k1!�X��R�rފ��om���֢vm��=�S������-��1���YgM4����>\�����5��A6G��F�"�˨1�ے�0��n"W�+��̰y�%��\qg"�WU�= Y�g/pe\�v��;]��J����a��]/{�le�.�j0�;~��V�O�Y�a�q]t��Dݼ���L��o���� �Na�=���2���X��:�T �W����P77-�2�5�� l��F�{Bnz����@�n`E��|������#�q���UJ�8�a���8�������`7JPi�lP����.�[��������~!��	0��ļ.��LC(������A)0��F=0� i?�0st!b�vY(慒myO4/[�λ���I���e�-�2Nj�dtg����G�IQ�gmx��=I�E��/�P��o�$�Z/�/X�M�!cZiN��9*x�*��\�U�	Ì6��Mᘠ���3�j#끺I�?G����WAd�_F4Ux�]���K��\��_�J1�����u�ͷ]V����Ns�ۂT��b[��܇���5BkJ;�+����
BMwi`~��&4��Mx_��P���g���p��綞�����!��`{��[�nn��7� eؐMy�2$�����n�v��
сFAf�@���j��ڴ�����������x�ӕټ����#���+}uрM��K�N�Q������r���Y_=�Z�UI�������*�����sP�a`��`�&�.��Q�Qr#[�=� #�,M�C?#�|�ڙmLCxWPo�/�M(�H0͛�C.�#�j����?ct��?����q�a3_����qCoY溁b�W�$Y�ngٵ!Vľϝx�T�]ܙ��t�z�]?h�5F��~VU~|��z-��=�n��r���8E���d}�5ϔ�y���[���N29y�Z{���z֙����w�@T���2wE���Rr�������s�#.�tP��.
���4i�z�fyq�ߴ,�#����pJ�ҿ��U�d%b��t7S���x_�fm��E�+���������^��t�	D���8^�9�W�����x�ɒ����r͍Y��K��!�B��I��|3ۘ�l�{��>֥���[I��(��v�M:h~����>�l�$�I���� av�R'�6�V�9�I�&H���x� S@[ݩ���\]�q^b�D1/E1!ig�������5l� {�q��Zz����SIC���e�Χ,o��i�}�/J'�d+PB�L&����BT:K���9���pP��&���^�J�+(�M���]�Q�Q�S����׆��]���Qh���X�01n`�ߕ����V"�U�xU���0q�����iR8�x,��G�������N����e)���g!�����Q�r�e��SN�n���Q"��̀g��NN�t�*qU��ͼ�n��|0S���e_}�����˛��2��n Jx�;�gn�0�B��c�f6�XA"Z �o�T�W�Zu�˔љ̖i0"�#S:��w�\,<���p�,��=bH]}?��@#efT���0�1���in� i�\�!�^e��9�[�]Lm�IC�<�̰��pٿ+�s��kد�k(k
w��a"5�)��F���X[=Rj�Na����7��w�y�#yF5�)x��#%s���uP���+xd����\l��յ�?�,�>qǎ��Zw��h�jW�-u�8���k��-�&C�e��(�q�e?��ú�=D5���!�%_��L+[m����3ZM{3rЯ�m��x	��'�����m��]%.��˝0�t������z���5m���Sxt��^}�{��"s�/����8|䈆=}�8��S�&QO�Q�$0U]���g����p��D�iK�?�1�!cgτ�w��y'� $���Y�DkO��♪����s@U��@`q�R&}�!q2��T�BA�=�<�b�͡�B�[��P��z���Tk<�_*��ܱ	sC/K���U�6�N�v<;Dt�l@�b��L���oR47�G��u�-Vm5��H�/�q��,�~=HA`�m4�y��]S-;eS�����2K�D�"B1I7�.*�˸ܬ�p���l�P�QH���(�Ӳ�g	�h��Xq��}�5L��J!�h@�r������WӬ�ǁ���:��p����(C�x�C�d�5�tz4DI�%��_���7�F[���A��s\-f�;Ŀ���I��	(���r�+��ii	{�8�I��Z �1��s!]��Μ-��0L�ED��T���
]���vԨG�@wP5a�lb� ^�����.������4um�HA�.q���)ч5�񕐻ȳO=HYм�\�|/U�a.J`�{�T]��G"��$Ћd>9H����5�c\^�] ��\M�����a�5>�7���w�x���'�����t��s��~�&�B-���ds�,غ;s���]1Jz�4Jv=�u*����<(%jj�c�Q�x���r���}�Ii��v�tI�1@�`f�R��:MZ��d�*�[�/�����X3����E���x�9�����ie�\�d/uU��⬌����!NC^�?�)4E3^�{"�����TV�?N�#�ܻ�0�P��:�2�Ǵ�P����)g�"���A�w�	�@���sw�Ճ�ԬM�d��DwL�0Yx�}���kX�(�v�l���1��'+
���/$:�K�:�̋�Z��#ͱ��K~�a-k�>�~9tj��p$'z�l)�e����)d�5�.�I���#j�>��g��@`���Ww���<xrE>P	n�n�2���G�4�|\s�1%;��_���6.�1�O�,�,�+jM��e�PoT7)��P��~�����+V"ץ����ķs�nw�5��Q����)B�S���[VT�q �"+��-
�-&a�����w�oVf�=�����=W-W>�z�v�?kkޘ�8�K��X����_��
'�k}MyOJ�~U��<��*x��8��P�~&�����N�g��G� ų��I��/���Igd^!�LD�f��D�.��Tx�D@�4���<ǽ,�7is���J�^]�+B&�v�T�^��L�[�� d�iԨ����}xq���q�VAl��D�M`W�#�V�e �0�Aib�_�YrַcSm]��AC�]��'.x�د�D,*��&����i��{�W9��ɥ�x0�&Y�I��Av������X�2o,��Q��W������(o�lB!�l�i�kp��5y9��� �{���]����P�DV����n3����Z�%�o�B#�'`��������Z��+Qqo�T==)���c2�ݿ_�*H�L��z���d�w��NՁ�D� ���-"�$|x	F��_�ڙ��֖�S��X0��77yC�>���t���\��i����1�m�oP����TUR%�h�'پ��B��S�����E��V��䏃�y�z��4M�%�T�oZQFx�Sh��(��o���0%ٰ���,����?��krD�_ы�&�`�=�F��w)]�ٖR�s���� /�1�;��k���������%<���d���Rx�*�1�S�4�4>��F��0:pw�	߀n�E�g��?�HL��V� R_ʹ��`��]@��B�/�DmG�.�7*�"W��ST�4� �.~�p�.���l/lv���p���]��X���?\�J��}����s��r� ���p��O��P�&�po˫����!�{��6i���B����Pég�J�[����΃`�o������д%ř�~oc���*�����VƐ�&�cB�&
;��E����	[*-�\��3�l�}u��#K�s|VOi\�!����I+_z�J�T8�?�mi�y��q��9�jd��]�����w�@���2�����}÷e�o(.ػ��s�m�ݝ��8�Bm�5���o�ܘ 
.f$ٝ�I�Q�c�1����e���f8�����|0���G����4MSp�^�gc�|�C�k���/�M"�N��Əz{t���>U�j�*`f������5c9t�ҿ�#�l=�S�r*��Z���N��{hiᮣ���S��%\�e����nFEo@�}�)��� 4�R��7*������TQ��d��3�)�.����c7�j)^_#�Amrx�z�Zlj��"?zm�yg\,��w�+����z)��x �~!��{����e�Rv�:��&/��5V�2c_�oQ�m�Ձu%�H?�iܠ���:��n����P/�p3`H��|�#����~�7Fu��)�a�q�d�R��5��ybl�'ϼ��9e
4n>!{>����.lҹ����uf3�:E�l1J+��#��))e�2���%3v�����	�o��q\ϖ2���o��):6���5��(M �[V�n/>��>V����R�&�	~�x�\pÜ���Tuu�[�	i]X���كczM%96�y%�9�[��˕ �G򾌢䄧�)��W���-�ϛm�A�FR��0o��� [+��咻[�<��nUr|AE����e�q����Gf�<���b�)����ߵ�4�������5�ЯW*�C��ܭ��=L���Ň���݇�"��t^�b���!��0���p�Whu_}�g���S���K��%�X��̸=A��+�dL�w�y3�ď��L7aڿE����#���a��W����VNp��i
�����Y[����>3t�^��KGp>�Ʊ��9��w��չ2`�m��R��(�F�\��*����~¿�/b	V��x,-��U�@�f ��s�~�cG�oׅ�"]X
��짏�0٩]w�9����R����$���;�vN0��f+�0V.VJs�&x�p�܆��v.~�Ќ`M�S��t�m�U)ۙ��xs�
�8��y�(�÷7��zE|@���U�ʲ�V�x1_�ۺ,<������&�^�ȟ/�i�2�����
�Gf�Aml$I�y�"?���!�#���<�7��������Q���z�:��z�(��f��y��J�Q�e��o�>����@��� ɫ��C��E��޹D��ձ�i���p�.�ks������yd���|�;X�(躥rQ���HM۫$ۖZ.k ��C��\tyt�� �E
�����9?�j��8n9*���:���A��?y��,�i���+�6�_~t�|������3�(zk�a�! ��`���{�@*��x�[��ʁ��;�w�/�	�c���t�xN7�"W&��Yȱ�q�4�m\p�/UGh�9.]��Ы��˝Z�1���&�W(�����Q~@T�#v>0?؝7���"�[2��Y��ǩ{���lPMv���EK�iy�<�!W����X���f�&d�m3��/W�I2��݋:�蚽��B���Mf��{���/"�<
�ׅ�*欢
A+���Ȋ��2����_u��^TĤ+�k^b���ܰ�a�fc�'��DO;�yaȯP����?-�}�r԰'t�'�ȆV�%���KJZ��t��z=$����?R�X��?3Y��!|�x@Xf��c�'�O���2�U#�����xfc���]M^b�Y��A���a�oxk�L��/�F�S/p�ʭ��ۆ��Ja}�7�		/_��䎷�u� �KB�;��@c��5�15��C[�Z���'�w/'4��:'0�n{ B�N���05�*�8���!9_��1�O�xN�)��%�~�=�=�Ը˸3\��v�=�Q�5�
�ű:���3$�`�h���ɘ���c�?�a콯^xL�|�g�~^�V\��G�<��[��"�JA�-��_�����>���gh$ǧ��+�\���Sϫ���Ϊ�l�^�ѩ�@��4˥�ya�"�iY���z�3Y��<�a��jx-!�h��DR�׉���Ms�l�o���K�hW����Lջ��2%�UBM��������u��^L~�,��)�X$<��XUPp~ws�ۺ_���Cy"�U(n�+� )��P�~�<\{b	q��b�g�/C���$TM����Ӳz����B�����๹�aZ1�b{xu���dʿ?��l�B,�;����]bl5�v���`ۂ�b�?7psG�'��:{�RZZ��\61�>17j�>Q��%��)G�U�r0WDxTo���K&�,����m�
laH2��k�*�FH%���m�u0r��됡w%}#��j�!�Y�2|��?�uz¹p�'��#�p=@�Rg'馑�`�2�4�Ig�n�Q,L��i���[DK�N�7?U�_�Ϛ&1ر�s������S��(�w��Tw1���(�\��^��
a,R�~#cE���ےZ�0"is��p��OԼ��
Ձ���l>��#'r�(ӧt����My��)�<ES#O���n;9ݿO�,ه��ba���'��F�f�aq!���DbF��qGO�D�{�"�Y1G��\S���_�t��ͮ�WPݵ�"�SF�hG�D����5�1k0leFI��C(���E�i�M�Zo�BaON�*��K�c��җ_K���RU8��k� �#�	3Uۨ�'5�A�D�=]���H���e'� k�'��Z�Y�M|�x-s��U�a�n����ɱ�ʠ)r���I��]���hfE�_��t�n�xGtw}�yN�3�Y�ru/��ܮ�)��Q�}X������,��	_����ؤ����4��L [.��Oj�N7� �Q�ca�e��v��'�O�1����ۀo�l�7�(�J�@��>,}KL��E~&Π�I��NV�=sa�tT���ן
} �Ā [E�"�ɳd���W��j, �Z�wfրOBF&uE�z�<�ٲ,|V#���P{��N���|��8�/�$�w�s<T��,kc��([э)X�P��c�<ʲ�5�H��y%R��2ͥ�T����?H
���/����BEV�
�)|�f�U�#��E)r���6���&a�C�����'g�×n��Od`�9��J�q��y�J�-R)�/2���ԍ�ɛ1����
�)�����UB����O� �eP8��<��?<��%1p�(uk!V�79Yt5����h��|�3��}`v��*4����0��u8���Ŋ_���	X��S��!����C��iPկ��~C��(i4t����fM�M����a���z'[���ڔL��L�Ds���S��a��=0�V�oS�~�A�{��w�]�?M)lV�Vz{eq��h&���}$��T±����[Vg([��g�W{�;c��xd����=�\K��>���}��sn��A�n��%����`@�����`(Mމ��Y�2��Y�a́Q6��<4 ��N`���dn����'s&��䔣�S�%G	�1�vo��=��`o���e�湩9m��Mjr��%k��y�r���3��%��N�����{�e�����E	��0������j����^j�����6�Y����t�ϱ_��i5�n}����c۳G+��x�],Z� �o�d�e�H��Ƚ�@a�y�K��^2�s�>�s��YPۭ 
~\���Y��h`��Oy\�*����>�n©2� 2eTG�1������H�!�������1���3������k�r��g�_�S7����������Q���T\��c����77uY=+9����i��ɨ`���#қ�0?=�?	����N��JXthh��t���@�J��R�u��;u�=CO*}�)���;e.����)�Ⱦ��!z}���A.����� �Oy%���ā���4ͥ�����B#��)nvcm���ёy�0�p !��=fO�\�	�� c-'5�w���e^D���(��Ob�ա��ǰ�}�d���g`^�p?��u��k��Mz�WeV�VX)������ �~ݥ�/ '�o�t�	��[�����z#�we9�ar��}k�,]:��p��;s��N!����/������2��i����=w����E��N�2������UoL�}�Yl���0��	�}���ֈ	g� ������п�ROag�}��͢R�oV%�p�1�2�F_��R5�V07Jp*��n.����ѣ|�B�닡���جZJ��C)�
e�	 ��)�Ӱe��M7݄��<?�Q�i�>߇��%H�ە��J��Q	c�W��l[�&(G�G�^�#�������BE-�dd���#v���JI��{N&[��ϼJ�H	���+�f5t��>��/�5�cRA��$(��E�gXOw��x�9z��n�Jͧ%ъK����XBJ�j�}V��o50�퓆�d��U2�I�) �QRHtv"�,��"(�Mh�DU�QrY|�<l��:�#����Y�W�.��t�p���0_�K��w���UzC�+�S0U��ȗM�C�k�:7����g�1�	s��H�/��S��m˳������j
;��,�����͒�Effq˹LLKE�A��r!?����{���Dzl5r���U(����_�H���6+׆9��L��7�)ȿe�h�ůom�8{g-Α�N�@B��,�(.H�.����v�.)����P߱��O��B��St'4�'1W��~eƓ
5��7����� a�ܳz�U��y�덃u+~c�q>IQk�l�E�|�d�Ry�-f`�Y�rC��tl}1v�D��Ľ }Vn�x��	�Ѻ�u�xM����k,����(�֯���X��O߳�hA��V��,?���z�Xh0�@�vN���C�@���5�#���{ ���W�z��#�æi��]Y���JwV�X���;��x����W�*��6����-�CRQOY�[�Ŭ0���+��o�L1��Z�kOqN�v&.��"J�}��̥&k~v�;�\K��/�uDvȋ �-!��ti`�:�z�>g�Wȕ;0�R���a��9�2�>+x�C�V�UC<}�t���^�v��c,���q��HT�Z$'��i�MR%�|׎�P�y�8�q�	���>`�psp������b/��N�T=��pb��`6�$�*y���?�U����^�o���҉Ï�'�y8����܋�`����T*�����#2.}1��~x�Б��� �Vыa-��2�;�%�Ȋ>�&&s��e�J1<�N�I��<��:��֎���=-d��i�v�:4"	��"��Ӿg޽���,�u��pǙ��8�� ��5�]����-�؈��c�t�u�����k�,h��yjbl��Z�C�U�� p�n�8��H�R��%�O��������$�z48�s��t�C��ճp��u�+8S��:��sP���+�F"�vm�!���{�U-4�$�5�]�T���k'��K�`Z`9���y����2]�s_���m�?;�jMpۻgo���S�����ӂ���U*�[�4�$����r_3Kڶ\~��pio婜q5��ڜ��U#��f(i3�0J,�ސJ[��U}�k�� ���Vq+��r��c����F!�L�f6�t�A���$}M����p$U�/Nt%g^�@��]���;t�x��̦dP�IpDJn��Lܚ'���U`��@qkA�+�74��F!`�� ��2����A�=�������k�WB�N� S;�����sJ�-h�1�l�C�`����4_1c�&ܯ~�C}��G���� �[�������^'{�pN�h9�y��lL|�aB��n%Y* �I�?��̳3$(�9�V��
���~���9 8;8H��6.v���sk��C�S�
�}3��m�g3<�6&FP�,<\�CK���$x��~U���*�c���������}jb���g_���B�WC�
ߋ�m����'�c�������6x>2~C?x�<̟Jg��awT;486<n�P/^K{� I�h������z�?t��n��i��ď��M �B��Ь�1���VZ��G����5�}^DQ`�bJK�`��¤�1q��Rdy�LB����Y��kh�(x�햌�͚���3�G���Kd,�E�>�trK�g�ne�_�G�R���0zU����~�"�a�天[�X	�y�Vc�H�5��`��Ѣ��n����g���Z�RF}�{2���[>�,�M�I� �o�A�3iqf���PGכ��A_��8��=���/��c����@L�ڕ	,p�?� �b���oѷV�z�r�*�I��A�Nٮܴ�Y
x�����`ֆq��@��|1KH��]I_i���&��h�(@����pt_ֈ*E�Hå��Z��ON\�7O�$��4�g��XW�*c����X�ǹ��P�[�O4����L>ca+�ϥԵ�5��Wh�	s7T�#\G�X�N����*����QW˻��b
���w�c��e�.Ƌ�r�Z��kgfd"Ѳd]�ؾ��5v
�V���hOF�F���������q�Ymm����}�n��C�?��}�
�_;�<:��lȰmx�_D����;�Cb|}�h�H�7W�4�,4:�@H�h�d���uB�y�i��1�qK����XkB�
���I`$�Xz�����r��ӻ�-Pd��4�6"�sՄz�!����;-4�Qe_�a�u+R�EFs��ߟr�w�9O��<��&n)�L潷ZA[̦ɞ=��V���?�|ZM,C�w� Cad���0�Nx�D����|�j��-k}T�ؚ��^75k�7G���Ęd�6���0�ӿ���P�m釳E8�Sp#����N+l��@.�(�°, �\"!bC��<�{�}t��ɦ�V�����a�z�Eb���'}pl΀�l��%<���]�Gq>�~���˷�	l���%�J)C=������ft%�0�u������j��v�p�v��Tv���,��Q��_ʶTY@�
ˊvy��u���'�D2U�� X%�����L��c/���tXk	����x>��bJ�>{���3�\8�lq�ν��G�a �V֊�Q�qe�K6u�n��$N�� �w��!�@/L�{�^�A��״Ў!��t��8 3�M��P���f�uK�jdOE<3,�h��G����t\lȻRz��4�[Ee7-��p����y8���-����)o���oj��펮p�7j��˿�9,����%�l����4�� t8"߉�7ʚ�,M̚lQy�n_�x��L2-�г�����}ݗGa^���p�bO��z���`>U3����G�.����c��W:NcGCq*�Oe,�a�K�fS��H�i��~a.4��f�Xv�?]�D���N؍%�5����	�g�ʊ�X&�'�qyq���8��v7����g��|�+ dm��O�~��S"�jQ V2�D�8�Ͳ���4[��8ey��tҿ��#�__	�*�Y;��c|Q�%M(}%��FB�9��\��E8Ǣ�j�D:�F��Df�}�����yկ�%�����Ygi�t��bKӟ�	�b(E/;5ݥl7�++�xP�<���D"6�M����W�➲���I��	�$����W��X��1#���V���}D���nN}M]��߄�a��ev��50�0�����nx�#���3_����:�(�j|�+C�Ʃ��o�۞|��Ե�tZ*v~��6U4�t�I���dGJ��} ���} 
I��
ʾn0����u�Rxl�KF��OF�A�'�G�s�]�歐\�C�g��l�|h��3R�G��xj�LSs��9�[��/s�P#�M��l���k:�sJ���YdI,xغӝ�����lQ��G�� �>�2fԠ� �C$t�c���7CX��l��	����Z)��ӣX 0�<�W�^F�p��h|����+o��Q�b����K4����9�ҁJ'R�ؘ���ky��a�I�z���/W<�Z-I���w��:��x9�6�HD�/�Y8PG\z��%�E���tJ�}(�eXM���!k(� >�5�����b�'eD��oǆ��Ð���у6��qd�ui�JGY�DE%�o1^������	�&K�Ά�]����R�*�c���z�����,i����}��U�`.Q���"����ռ:[�O�4.�?�t�0}����C�h���z;5�6ץDծ}�`�wz�<��u���}�\�ʴ���|�z��}?EI	�{>Y=<������,y�B�79��,.)����瓰h�5�'�q4�0h�Yܷ���?Ŏ�n��M?���ŧUK���v��=����o����g�[A����q8p|��,\�����U��% �����S&r|� ���9ʙ�i��`E�f�o18����?���c ��	#��g(�D�$8`��5�k�p2NSr��0ab��A+�b!�!�|��W2�.�~`�t�Ƚ^��p��6:tAt������O�����ɿw>'/y�+��NăEԜ�93@P'��2KV㐏O>��Rt�3;�1�>�'Vm��Ns������@�sl���7KFp-���͌�f�ٽ����|$�eE�Zv�3������L���4!r��X�3�����Xs�v��ϋ9-um!im=3���|���y��$t�-�r��֔!O���7�<�`�����>�3C��.��+Y8�����X�;gA�3z[F+.DB
(�U:y�z�J�l� _� �hD���ć}z#��{�n�����Z�Y��9�;��KX�ё��U%�kA���0$��vC�^��I��>mn�pp32�t5��-�h�ظI��!�����O�Κj��اB��Ci�`��-��m���]�m�w��Q4�ӈo��H���p�I��AJr������}.�? �ٌ�]��OZV�'�����/:�S�A�p�����h���F	��n�O����~F��?�\�H�����^�+4ًA�̉M�k%n�v�r6�ۮ��c��f�럄{�4��%�����(��4R��v�p9�ʔ&�d@Åi�{"�u��П�A빆�T-�n!4|O_,^�����]/��Ş��8%�n�fPNSQt�����QI��k�e���urDC�ӝ[�$^����G���4]��c���X��O՞�{�&�~~x2�k�� ��y�F�@_�XE�)H�<r�$
�����.���c� K�m���}K�0��ְɷM5'��������̈�ԒbxM��`�h�D��mF���ӊ���6�����b���W����a���<����͙ٰ�Hb�k{F!�:�{Js�u�[��:oCEkA=աU}2��L�%���:����*���K�Pi�5��jO��CT�N'~�;�yR����D&��NRh�~��LQ��_v�����5�XeɈ����,(��So���j���L���VYI�s�Y߆�4q�)!��t��D��!�4�̀��r$�ځ��$�o���Ӓ}��@Y��aq�0�0�����)[2mo�d2�&��7�A����9 �(Aư3��p�?ܜ��:B�e��C�&���O��X�~ъL�?�3�r- �	n�V��.j}Ye���v�l�c�&�J���!��:z;y�B�>��{"پťGr�Օg�G�~��Kn�=����C�����c��@F�9��E�5�Z���d�;�v�p'�F���2I�v9��o�M]�������Pӫ��P�X�@4��S�����.���IC�\���~�m=^Ό)l�t�'���M���K�LL�Wg�`@{Ӈ&A�/%�h}m���/F��-���A�)i^��o�u�~�{؄uM� ���Hざ��_�5���A;���w�rz���0#���k̉���L�Z��}MR[�-h�gԎ na��Xg�`��+-���\��9*+���i�4|����E�p��C�]R���	�+���U�`mdp+5��Y�
E(n�T��\������i��'+0`��l��Oq�j��k$O�TP�1%5S�j�T�J�B�h�$��ؽt�v&�]�O�)���Z(�q���r�!j�P���5�?�0����A-�Un["�P����7|�ƫ݁I���w��!x#DyC��ꝣz�ll@LH���r��bU�Û^��`/�Z��K�!���m���s�����z��Wt2��ƎE�����P7cţ3u�W��1;0�@L-bլ���X�3M���t< �[� 9�%ػ��u#��`�֛ܖ�S�[�`��*�zsi`����H�.���;��տ�jZ�os�%�g84_o�d��;K�����윤�C���U�nS�5��Y�$����L&u�7�rCN�A����,�.p�����s�>�����)����ַR)��r�Y.��o�����t�T"y����V*zytO�����]�����D����9���\�S��Y�W���Cd��}��o&� W;a�D.Q�s��ڑ{��6OT���L^s�7{��,�������Q@1r��X��@i�	���`���U�yqw!�|1�w��0��̐��ً�]1\�6�$�z�����ҡ�[]ߖ�3���<U�}8��������M�4�f�/T�n͘3tR_��w�،V� �Ue�S���B�;����a�]e>+W\��`�]�أ�|1,b����E�Y\�yI���Ԓ��񗴚�|m3iZ�Σd��l�/�ʘ����=*����B��Z���7cL��������-w�:��2#ZU�n	��
َ�X�����CKV���,�o���������߿X�p���O̓L�4"ut*8~M�t���!�4O�t������R�N��N�e*�%� \��om������I�@��{�L�}�|��r��@�]0L�/�nE�hlKД��r�v�O�7Ir�[X݉A	�q����.1�=7�?�2�Э�n�m�q.|K��;�m�X)���4wlyw�އ�9N6��$�~��!��ݝ4����D�~����3���IZ�K:Ѥ_<ؐ})5�.z�W�8X�`�g�C���q��Z��99��2���}�P7��J���0��:�	������Ϫ]v6�t�`��F\�\>�-���(M�+Zf
;L�s͎�?�����zjmR�'P�vB9�����HZH��\��0taL�Ny�����Ĥ��Ѫ�Fq�W<����\�4�t%��a�A��g������>��x]���'�6�D+�e��NTJr��%�*#�g�j�k�������e_V���D�}|y2H�3��!oNJ�B��`�\��YB���n@�Kk����p�+�jd�bI������|�\8g��&�Cr!_��y<��B0y=���'���H��xs������ζq'����̎ X�u��b�ҟ�e�H&�ptr'����x},�qA� V]�L��������Ho[��q��̗�DF()�H����>���"L��S��(�+��@�� �}*�\�O�IFΩ$��S���#�x7{6j���M�RK�g��V=���Q��~l!���E� 2e�ʞ��>x�)�^������{E2Ɵv�lW�׃O���������
I:��p1-���?�!�f�e^a��+~�bJ`��A`ܱlY��.'���,���D�ѫl�L�$r�uT�1*�E:�gZM;1�s�8�5ћ�4����P�h����7�K��ֵ�tEo�l+��#��)��@��>�uh�Ր0Z�?e 4��V���������䐲]&������A�Y���T_���~u��F�����?�k��#����x�ke(�����'�Q{�0��d���t���1>]!BD�K�,���m=+ǝ���ӝy���In	"�.Q��(Ę�v�TNn��?!��8d�\D���L�a��)G��J{/�w&.Z��C�g�~UT���y�7�c�����C��p?mo��?��R6�
��%>*�W]ց�ά<�ޝB,�y�����h�r�~2�75�=j�Z(���ׅ����E���zK͜�?<v���М9�8�n�?U��%Ӹ��!!�ݫ^��� s������#X	��o�%75b�ˈ��4\��9���]����!����*��J���%���X�Tz���<P�ɠ�}��
��D���|����t���YOa�������z
y��:���Q�;�Ǜ�i�$>�v���gl5��&M�<�v�����̌���ʇ+u��2>0�Ye�篍��|g������,�ks"��L��N�+K���y@^)qz)c�4�t�Y��	�䬂8l\�=�k������� }��\r`�kl���4�ʈ�@;�U��B�mu�"�).xxa�T���M{��8#�@���uL��	�f��_0 ul����v\v*z�˾��������<;
櫄8TW����!���cM������A�D��z�B�:y�v�C�� Y�sh�2Q��^>'��̈́�cl�6xnE�^J� J"�e��{��5z��!k����^���|
��v�FQ�ҥ@Q�����!����l
�e�V�q����m�"�zE�cfn��l�&�p��*2���i%�=G�8p�6���l��鍓�Ǚ%���X�i�;��e6'�e�b�Zx� Ȼ)� 0j.�1¢ZpA��ڱ46L���F ��łr�+K���A��Fp�鞔�I� ��j ���3N���?Q�5v]~��6�W�1�&.纼���N�.����O�=��|Ё��)�/��p�<r����S'���PC�4�rB
b�z�\�κ�cC�+ R4��/�t�	^�ʽ6r�m�ѩ�&:�$be�cN	��5�t�C��`���͞�RjDYF(9�;��k	4Њ������E&�Im��s��%�]H�� T����L��{ZU�)N���lܣ�o�����~ױ���3�d}F��]
:r��<�9�q��A]�i�f�;'��:���'�9�Jۺ�l�[�*0�����Hi݉%�g_Z�����#
Vgo��{-�;��H���r��"Rz���~�q;�+B?N%���2!?9@���<|�X]��:����s���q��&љ䳁{^�u���4�ߺj�N��>?�m���D�D��kb��;Z�L��zSe�Z�j�~��}�����`9�w!�3�RJ9�B�~��a��e��7�ܔ,���-��:��
o���XT�A��Bl;�~��ٗ2��V}��DF��EpG������~���.L��M�p�pP�7�`H¶7Q� �D�,E���|��{I�i��"&��Ֆ��^k�~�v���T>=���Z��X����X_�ޅ�x����E̌pp�(��)(C��G�5E��j�|�7�-v<&史<KɧL�'��ܰ�A���������( {��U2~?m7��y��W>�z���y��sY�fO�<�3���~�|����F��<� ��|�l�q�2�`L�oW���Z	��FE����
�x2*���07jtԬ�1������r%\�OY�n��	a
I2�����Y���U�'�w ?�'qy&�ϊj���'���߯`D��Q�y*G���dw'A)C��ą�v ��U9�������j�vG�E=+�4�1�FF�U��FxB�H?
I�*�^4�.���P�����IL���<5ut쓮��	Gj�e�>6<�x0&���R#!O�OXX���Yؑc24<�q#Y���
�# ���Ҥ6G��˂����fI׮��m��𕯌���e[��p�7E�}�������Kwo�j�n�T����t1�;L�B,lZY��}4���$ّE���[�������l��qC���?�Lql�e���B�fo:!�b�!跉�Ⴞ�Ip[��Z^�%�.��� ^���DP��aF���� ���g�h�d���P��C���j&6����r.��|"	I�u:mP�Th2�g�ª\�,Տ\����.��53!Yf���lCϾp�@i'������$A�X8��;D��&|�Nf�T?�P�hI:�)s�`(����;Fp��)�՝�F�-I(��⑝ ��`�AO܃m\���`oµ&�4tU�j��\d�("��:g��kez��0��vY����p@F #pVٍ��T��^�ς1��;���ܻ<+.�3n��P�a=��O��Ie�h�5�X� R�ޣ㹉�;8D���C��=���x�a�ߞ�_���Ҋ�671<����	A0(w9~����o��a�����a{����H�1�n2�����F`��4YV2�AȮ�1���`����`�T�q��3�7�B����z��=D4.ǀj��]�YΡ��g��P(���?O�Vk��.�[�Ʃ�!*3�����=LTI�h���eV��*�u��k���Rc�e��~���A�]]X��_�g��[b���)�nUym5W�������CM�!s=r����W��PU��!j��^	«��a(�_C7Ch���+��pD�S5GI:q��Z�)�w���:�'v#�x�����={�;�LQ���)3-u��6�L�S��[��`��j�t裸t_�ax������n@��e����cW\A�{��P�=rK�I%)�atk}F��B/�	�SZI��rW�� �f��ax��ʪ�w��=($����3o/05��g�׈$&e6`��z*P-�C���H}{��Հ�3����49�C�����n�)]��N�Jh%`G���4�4գmJ秿Rj��7��Q�:&/�Gj�����wYd@�ң��=�=I�.��;���B)%7�S��)4NOR�4�l�v@��^k��ĺ������m�j�(n���NU�M@�pA�|�1@��L
��	x��R�
�����CA���fm����53D�v�h�D��/�r�A�ͪ ��Д�󀩩g1��9美 Y��Qw�Y-�������������.�����1bk�Q\��5y�O�{S�̪~	����R��XU$=�4J�ɶ��)W?�{z(s�қo���WЦ�xe�e��׻������'�6��MR�����Iʾ�Gҥh�=ton����\�Y�"7�w��=��wk��a*8�_~1�+�AYEJW]"����4�ؚ?���<��2-P�h0h�#������_��A�]u�h JLǫ^�ޅ�p$�0������+�8>�L�Η%�tG�k��=T�<X��@� �⣎����|̃9��y�����H�I��܀;���1YT�_�.m��'7�3Џ�B����|M;46d��&A�s�o���}����[�0W� ����9�}i�ax�/�>�ѽ2��VR��K�Qdo��Ƥ�����f��-6_y�>�vb�3p	�7v�Ѵ�S�9����ƷI�G���� �zy��r�nؤ���}:�<��e��F-��Q,)�6����8��hN"5���4���>j>��>!)�%y%g��Ρ}iҿ�pS��+b�~6�Y4m�L	��('5�X��[c�+RUY�,��������5 ��2�r(����0l��e�m�+�-��y��U�щ珝�`�9���j���Q�S��h�:�4�|K�Jk���_2�uQ���R��<qAܷJg�yϢ�}Av��H(D���G�W��W��h�����´��6|�i�:��|���
�IP��w�7����!�߾�FqMFw�#7�U< �^l���ö՜<*�l���I�������v�I�F�(oyx4GS1eBQX�)׭ ��Լ�����@F$ZM�D%%.Z��ٗC*!v�}˒��1]�9����ԙ4�F�k�!�\��fs�f��P��7��JrLA%\g��P��#PśB(�4���
��W�=1�x���D�&���B����Q�6��Ht�dz�.�m�.�]��;Y��r̃dj�c�LJ��$n�-mz� ܑ��t(����B�'�R�]֢�'��$� ��Q���o;@��8\W��Xx7�+B��������ziv�����d;�9��g��N^�a*,#P��_���.aӦ �3UMBowgL�(!��JW7�Z^�aJ	5 �L��������d����������v]�"��啿Gs��=�PC���Tl���h|�����h��q���R.���i��?#jO�B�`�%sr��VX���	  \D�n�D�q���,pr�s%�k��3Ҷ�
E�� L �/7V��j�!�rG.���J���̗B���/ܽ\��8-V�&��79�U.�)3�t�S�O$ش8A�0e��A��f?��P�!�z�0�~{�`�J�a��T�����H�~��`Hp<�q������b��$ۤ!��ċ�>�����{�L3���c�,/���`�ڢR� �2��Ҁ|�%��O�5"�4�|�a� )�f��G��3�A��ℶ�vU�>/�*�A]ꦯ��P����_��GW�rIxX��F�����.��=;ǃ�*j���|=NN������ǂh3k��:�+�T����q6�˟�L�q�y[F��'"��I��Nf�m��+V�$)�V�Vw|s'�7�dt�9h=�n-�v|R��j�&���Y!@�0��}�-N��*��.�G=�U��_��?�^�.iH����ӄ�I�<��2�F����}{���&E�kZ\�k����>J.&��]J㈄��T��c6�{����x�W�+)�� 8�.o�C&���>=I͌}5�_��U��ލ����'h)0�X��#1����7��\�>�VSư�D��k�`��0XP�e��� zL���؉ba�a�L���kh��u�<�f��� o ��&[ug�wЌWq�Ȯ3`��g%�wS�m�(�Z�����7�"b����#�� �u�!r{N�Q�TH'+[<+��N�TE>��)~rӉ��*2#��TS$����[o�0d�hD�ԇ�(C�eR�e��͑�h���,~�Կ׆�I��Q�'�*��f+H{��#�&+<�?�������vBڵ[Zٮl[�a��q8�&f�q�FRr���XL��r�U��Qb�������h��xG,u�rj�c�*�.��&�b�2H�5����(�m��d��kt�3多��xQ��v�c�֌Ú�+����Jb��].H�J�}�{Cw9���b�$?�:�A�z��ap	��K?�L3�nQhw�=9>� W��1��St`7������!j.T�|�Yu��~������9���?a�V2 ,������#�
���h��B!���/��Q��\[�c����|(�F4�����t�b������؂�l֬(�̉�C�1W���l���!��t����\�6�$-HI6r,#5mU�����`hq�����K��Q��l�\_#��.ᵨl@+�#���� �64.I���z	8f>N��`����+9�v%OV�T��@���=�m�Kfs�����M׭M�N�4D��<2&�֖=�����1	�m=t��ކ[��Ҙ�.&�3?g\�s�%|Wj;�W13����NQ���,#�ϩ�X+�.z��尸�H	�d"��Teir�+(xBM�
�cҪW0,fvm��1S��f�НQQQ�6���``���zG,s��8�)�þF�؏���l�p�%"�g"����� � ���$�x�1�'߈ �����'�a���<6�ۜ
.� g$h�����/*P�OQ��m{/Q�Kį�M�i��1Kuk��Η�(?�{Y�>3�@��R2epg����̎���.�#���D��+�0���_�&,z� ��,H���Eu|2�8���cW��,��$^R�mA��8�؃z����
l>������n-�I&G�B;�)�T��>��^�R�z�K������	�G��8\ �Ļ8�G��¯�6%9�f���3g��t�5�-�Uy��ӗ��{�L
Yw�g���w��L-,�!7���#�&@��؊�� �-�PRD$y[*���z�M����22.���-7���t���W:P������u�M9�OG�7l(4-�y^����5��g^"�Z��<���z#oAOƾߦ {��k ��O�b[�/��Hg��{�����'�ˌ�k���%	�2��SճS��}�Q�� �����q��������r�la:�Y
��W��c5^�����Zxt����ZmMLǡ�硹��&}��Zn�ZGH櫜&*U�(bV^�4?.�������={r�c�@��<��o´�O.�t�e��h��q�x��ҟ��w�Q=�ѷ	��^U��L���F30��<!k�<v�zr�
�rL�1��hD����@��q��zm�q�a&G_>��!������~��	���t��m/$Ha1�`f��<���N�
y/������FFR�ݰm��s�_*�}�;�����3*���a˔2A��+N�8^�E�����	/�ք�IϠ v@^�P�9w�; Q�m�bB��G��0���H"V��᠐�!_f.���w�Q�m�t�]ζ���+P�ؤ�'��
�wm�����YQ�-�
�[�a$�����K3-R~-Q"*(邿?��@�*�9H:�<�r����$r�s��Q�TZ���R�>{���'��j?H�Fͻ^x8Bŀ��\�z{R5��ѿ8b"/n�-�n	�1V=�Yjn��C|>�~{����4��O���O���O���t��.���w'>{0uP����_/���3��u����_���]������!�(���ʀFK(�����V�jV��?ˊ�K�<Ap�xRi#�!�se2Ӆ ў.�c!�<нD,�#��F%p�� �?���-�7��eW����(EӘj|I��.q�F��Y���E���e]sc7+f0KI�#�j���'nɸi�͋�)�-�+���fg ��>z9�����?v_��&>.��(��+�މ�ësIh�V.��M@Wgo�6r�P�+S�Za-���8�c�`�?_�N��6�_���A,{?OZ+�a��]�5H"��'~��P�;�g ���'��3�U SF������6�9�M�����>MT��&u��?+��[$��t��fnoc0�����Hg��5�����䬲�v�)� �]�%�4�$	P��
?�iF�^�XHm<H�̔�Ov��X .����,y:���`6�F���B��fx������^>�u��E�1d�Hv>F+T���5>���b�%�.؍Yr_Z��#�vf�/{���8��w�_�&��@T�Pjq¢�J���N��k?ZF$�م��FR?k|�ѫ]�-g�}��d�D��w<��E�� q�s��e�p�Z�OB�������<�fI��	M����
��W�HEǢ�2�j��EP�a�ʅN C7�*%��4�N�Sk��ӝǊ�WﴻO�(��ԙ,.��-q��LOF�v�ѥ�� �,?�i;*�f,BY@�TN�n���BE�:�2��N�'~T?P}�πx7F�����a���v�+�}���M�K���I-,0� |~�i��v[*J�t��ܰ��|^�����Nw���,�u<�����2>ͥ�N]�@�٧)�g�b�2J�Idv$ZMu�w�vx�I[rvm���t�Ɇ2H]�v�3]��)A؆<2*�=�E�;2�x�1\s�VUxl�/�6�S���I���J��	_�c��4g!�n�&�v|H_~��\��?t�A%J��v&%i��cx�<��۬���e磍>:އD�CB���$��U�>����M�����x-��dE�g��(tEq�fԾ�}AÉS�-��������D��'�'z�E����f� Q����ξ�)��|�l񓈿��L��8 J��/"�b�����L����;�=́�f7�z�/;���y8� �۩����K��W$��)"k?u�]幠Z��3|5��O_
=/-��	�0���H(�1Mpܸ͠T ��.������$�;@b��c��Yd����`8�n�aٖ�� �ǵp4QWqI�s~o�R��N::(���L]�k��eC��� �ɥĲ�"0C�����|鶘��~�o����"(�a��tmt�J3�-������x�S2��`DiGϝ�)2t��k����xu?ǧ�W��Q{/�ܾ��?�nB�qf��F���._�Zoݡ�e7V����~��9��z���e������+"XI��?�=����j�S����&W�E���UNIcMQ�z���e�n�g���Nal1�G��_h����%�8�X����ϥ��q㡵g��s�S��\���#"�p���PO)�z��/���q&)Gz�2��xG�����Xr��$'����p/	�0E��� :S�l�Qb&��� %�/��_�K�e|��rNj���D/S���ICk(7�\�Iʃ�|�]�g�p��y?�@���G�#��˰E���-k����1��$�^���$VJ��pɢ��������D\M5c�-g��I�w�B_&���q�u`ON	 o���*[���Ӵ'Ñ_�s*��v�+���&<�]
>	�����A�R��XL'-�
Axl���B��à�G\�'���	�!ɖ#⺇	t�Q�kk�z*X�!�SP�|�=�x�sD���`�u��!���)|3|��O5u�M*a��v�6Aϫ�B���砤�.�������;.�@����3n�9>�ku�,pK�>����M4�����c����v*ۉ����Z���|�A�1�5K{T��{#硤Y�4J8	t��/rk�N���S62�`^���'�R�\ޗ���d�����>���Pv0�"�ݖ8-��w!�����PH�� u��T(L�3���B���K���z'-7�.Ix$���e5=s*�`[��
<��Zzٖ�g�����^�|'J�`G�M�w!��.����)�2��P!����/twk��Kk�袛�Mbv(O2z�����������*l��7Z~��8t�E���լ1�"Q�d(��rA1����c9M� :�df���RUö�Z6�pM�Ծ�������X�ȭ�1�\��/�HIG�F%v
1��� �% ��)@8��n�Y>j"g%�����5, ���� ���R,��k�ڡ��P�,�-�֓�Ոʖ�;(@���p�:N�@��9���W����d�Xf���fCp"k�;��봒��X��fۻ���Sg��"G�q�q}���-��Q=�y��y�3d��	r6~)���Ps�*�K\%O��6a����d;)������.!.ȝA?r�Q�lة醱��)�j����a_>������R��:����<����L|b$�5��o��q$7�r�0����7td��}Ţ�w�}����uuyJh�R�>�x ^�u��j.�����G�&QfV���>洧����7Q@�2��eE��3���!MTl�w[�Q�Y����{�G�����������8��݂.i�*|�`tU�DBWI�+\���ҳ�T���*�=��������q^T5��LO���W���pVxdw��@��#S��4`�=�)b��S%�I*&��8���C�� �7Ed�Sl�|aѿF����;߸���~��]r�e*��ܞx�3��'�͉ڬ6fLd,���s9ybL�ڍ0X�1��V�ƛhW�>�� �-
Цn� �Yb����&� �o�H�+��H7���Ͱ�����L�Y`@�. �@'�H�)�/?�h�D�#*Py��-80�Y�5�bJ郄\�;�-�3FFݴx[�1���P���\�4K��vfC�O��E~������a�c��faG�o\�IBo��̃a��f��J8]0X澗ߋ� �K�p�X���i� ��&�[	�%g�S�f��}
���e����)g�UW�m�M��a�vQ�gQZbR-�5�V��@+�)�TI�2^���Xs|j�r��c�@$4$���C�^eT��Qv!ޫ�̔E�$���(fl(�����fx��+E��>����98n]�2�-�+�:�J�Z��Mu��c�6;��f��-Â*�ש�>�K��������<kT�=*b�o��Ӑ��q��Z����V^5�3��/�6�%P�׸ĕ��x5K�Ŀ��j�EX�O���b���&�������w������M����j��_C�S*���� ����cy�(�N/����d����~��SV��L�U��o�e�~��pӡ��T�:\��L��X�J�|6.���W2ٸF���޲��qt|&J�{We��%b�3i���(�ɶUuSݸ\�I��W�eɯeԧY��]K3��H�+q.M�"�$ �iV��_�ѻU��9�E+<o i�w�G�S�!;�(ߔ�,��^}�-�MΚ�'ߋ�k?�1+�G�(V'��h+>`-�~�$1s�P:?�ٙ�b7�32���!�o�?��,�~+�hLj��w]!q٥L�\ٴ�K���Lu��k������ix���{]���Bw����)b�k3�}�Q���F��n��-?Н�<S��j�|���
3��=j`��V�2/?���ܸއ��u$�C�?SU�hR��KxնH�Q(Q�c�$+ �<��rЌ�y�Y��G"*�dW��eG`D��n5h�&���G�s���CZNf�r`CuF�4����\����A�״���frt�Y&�f�Ei�EHaW�km���X��xI]~�Y[���Q������+D ���&��>�i!D�Ai����яR ���g����=,�]���1�	BZǖF �0;YJɟ���?J<�ɗ��o����b+�����85���Fg��_BC'ى���"yfk{� ��n�Z��M�_4��n��	��@g�p 3b����`�c�3P��=A�h���7��@?�n����M%�Z?�������`�F��OD��ю�:P�an�&=���-m:�a3'���oWｓx$��������,��uZ�U&�z����;�I��w�1[lW�]k����1=��~�k���z̏��tW�\)�'~�/���&�z۶6��f,���O�%�9���ke�v�Ճ��)�R���B��:;\�9����x��T	>|0��c�g���2��P��f��(`Y:��F.�en-��[n��|��P���z�]c�C��Ds`�o	�� �z�=u��Dw���Y�ѱ�"���L���r{� ��>
O�΂3^{��#��L,�fª�S�:���x~Z�u�Ur;r�P��y�<ۏ���U���7V��Ie����Q��]$أGc��A�4ؠ�^�E���NS�5�~���9?=j�ڕĎ��������l����u7��*J�}��Y(\�YP�{f)0�z �>�K,�P4��v?� ��Y*bxE.���k2�#������^t�T�_%�ӛ���'�[��#�~D��=8jZ��=�k>{ST�/"祢�����f5��Bȫ�
��y��7pη�=h\�Cx��j��.5늋+�H��m�"��A�q�9X(�5�e#��6�:�����7״B/N�^T"�PwmX۽��k��X���������]}��&+�%:��O&�`�uJ�e���C��O��K���:���-��ܿEY:O���SӷOA�"��+�
�T��K�,�*�0���D9� \c*r�X)Y$5K]-`��K�m�~��� ��o�;)�?�;:@{z��S�1����ʍ-�	Bs���3H�-���JD�NH�=�^/0���a�\k5�Y?B2��J�#���+�#�8M��j;6��U�m��1�S��UC8�}�� l���sTb�J���E�nS�|f9ev��z��<*��m���^o�ً���	48@��x��%2�-=���Xg�e�?/m�8z��H]�d��&3��f�����k��5��c��H�_�lŶC�e�\%W����c�1�t�P�$�@ʔ�
��謒�?�6߲w������W��2Me|��b������rd0���:-5g�V;�u�ݛW0`���� ��ը�{\���6'�4��=5BN�l���AX[��բ�$PXB8�"��Z��]�!���A+"؍�!"*p!��a��2t%��?I'�Yz�SH����Z��3Cwׄ	�Op#Eā��iq]¤�����S4�ɍ��ݗ7ǟ����_�q�8ls�
p��W���;Ŀ��C��X
	7R�2��'A ���5a��%ML�myG�J���s]7��BA��������׫�U�Jem����Y��{�F��a��L�,w�����Z"w�Q�����!�.qXRU�twQ�O�����8��,Ɩq-��� 0�t�SeX��T�t�9u��-�R�s� ��g"��i\�7}��jX �?I/�*(n���������������0l�'�A¾�CT0�#�1ax������SU_��8
�xC�4�~��{�'p��a�������-LF7k?�ORa��� |I��q�`#��8U������8(L����=x�u]9�,&q>b]Qq�N#O���,����5�	��H�b�]��o�ԭ���W:H$<�O�wإ��.����Cqd�J$�����Q�uS�N~�N ��|ťw�_�p@&vf�#]E���he)�X9��Z���u&K�	���w�U-l���2��Z�����M϶ƾ��0�i~"@��#��������9��c�{Lâ��U�K�1�k\`���#?���VKM�V���t>`�`g��G��B�QAs�:��^H���R������f�A���\�hZ`�T&υI��e觛IAg������+<���ؑz!�f��|�=c�Jlms�`�g�ۂs+���)�;��`�up��΂��}Fk<�,+L�����;[P�t=� zL B}���m����ZF�'d�y�7
��-\���Y+��I?�\�F����-ƙ$��:�%8.i�D��z�B[t�+-�3
g�!Q�	U�եc5]��.���Ǝ�Y!ʣ9$�qrv�l�Q�8��kY� �+���Ѿ�Cz�� ےE0^���U9���F4�b]��}'���G@��<뉌B���}0t��8�bXn�Eq<��+��F�Vb��6K���
��"��Ҥ�_O1u^�<��G����g�9�?�W�S݋rȜf���@���S�s�C��|�\�{$Ke%��ſ�����h��	����R��w0Tq��{$�?q�jB���o������V��'ʕ=A�f�T y$�S�ƕ�-���H��2��֯���
G����(��7�z�0%G��SBL���*q��:��k٘��� �n"@!�j�#U� h���f�L��8�Ǯ|q��z�'d*�1NL���6�� Q����ˣ�h���GCj��g]3��� y�= ]Gb�?2����nD��3�ۣjpN4'.S$?L��B�-�}�k൵�5-Z�s�[�(��޺p�PPG����c��|��)���5ߣ򔧪��j�[v.�y|�iOR��C ��Ut�'��]���I��cv����iŃ�VI���)��"���F��D���}�$���"1�s����^b��=�|��i�uxn���/,��t�P�Ӥ�u~V�8�)��2>u���	K���ߢ4��i�gϗC����pI���Ut�c��) �Ť�3�P-3Dٞɞ��'�3_��e���v�¤��L��Wh�{'Юu5l�\�9���%�.s2M��_�s��7�� ;\C-ZǛ52ǽ�z%9̼B����Ɲ3%F��ՙWۂE�-o����xff>Y��T�4pM�c�V�߹	c��uU�V�?tk.��÷��U=a�Z���R/�3ǃz1�<�;�e�#m����n�^s?M����
GN_o��N��;�oR
>!gߖՁ  H�g�;u#�i�?!s�'0L��W\Sx�K�|�%�p	�6�5V��m@�X����$�qX��h��A����L�q*�s���hTŰ,@y0{$8ܮ��䪮A��b9��tR��욷t��2O.��	 ;¡l���@_��U
�jv���S,}P����$�R8�����#�[_��pUa��I=��rk�*�^?i�t7X������<x�+��l(�FC�1�ܺ�����XBEU�#Dv��U�������Fb�-��|<�����s'�<��|A�*I ^l$��@0��X�7�T�z�#�#�r�i��U'8����$#AUs�z�У2<J+�U�QM��I���iz�r�Ps��Kq��rXȨ@Z{��%�^-ő�:��j|� 4=��5(-jI�87J��c��5>&_�hd}u��weSY���L�j���2�4��A�:���ޙ-����գ�"�h��l_{�6%/l8l��s�M�6������0��W5TRJ��V<�p��T����ki�����?�� Yݖ�r^��8f��Qf�	v5N�b7��dl?���E"�|�M��@>2�դ���N�0��wԲ�� ~�#�Ng�׊�p�<S�;~ퟕ1r��"��h�7Uq%�u؎���$���><�~;��u�bH����ΫmX	�o]~�I����1ƣz��Cզ������L���9ꊤ{�BC��:͂���r�M�v8Jz��a�L9�8�+xAx).���a�VD%�-)ك&�I�`J�����Y)/7L�Ò�64�
6W7�D݃W/)�j2N���HH��������C޹�c�o�nJ}̑�x�)\� �>�C��7X\T0	61>��>ߖbGA��ӷm�5�
OCב�h�pC��(1��j��3g��_X�{���D���禈>�d���=�����}t��³�F��Z��W2#�������#��NJ���A�Q�۝���P�`�Ag�h&)h��i/9 /Tr)`�|�p��H�6J�� �N#'l0���\�ء�xߋk��{�[�9.3N���oX.�jY+�_:��<�^u\5~�����?�?˨
uƓ�{H��O��]^�ŅP&�Ӓ�Є9�\�Ȣ���X��ĳ������ބ���#��"o�=`�*$�Z>�e���7��:^��w��O�'Ddڿ�҅�h�@L��f)�K��.{CA��CG"z����,�EI�	�g���3-�+ۂ&#RN�H��B;��L6�5�y��7J�\�x|�B#����3Q�'ss`�  ��P�K��%C�tA��i(�C����qf�=�V ��ؚA�!&�����F�f��&��Qq���,��%����/���'U����V���;4A,F����+Q��>��1`�g|&����	A��"g���%�����k�t�2�b�x�wZ��qr|�����B%�Y73�Svtx��%mk�n]�k���c�8������W�i����j����mI\E���Xl(	~ad��h���#%��MGV���	�<����m�$��ц�S,4=M�7�P9�@�����Ev5\� �R��xb�qAZ��� �-;A�"������p,^����ԍ���F(�w(�SY�+�t���,m�Mt�q�K��-�?�Awj���OgH�!�PBb~l�/ �ۀ:��o_uu2���ܒ����%���7L�T��D�a�����n�C��<�%a�ձ���QF�׿�y�WZE�pf�����%mب�����S��W_���՜�B���l���L�nL.�oa�,�T�w��M\Th_��qw��$�X��ֽ<�[4V���w��=�zun��&�͛�h	)|��X$��ޢd��Π�}�zG��~�(g�v݃+��L�ζ�K#o��/��4���U��7�oi�~Q���d&re��hO�ƫ���`r�`]�� �a$e�)�� �Q���s��Q�7;Y�_���	�D��%q�e�<G�#62��,a�U�W���3E��a�_ޅ�5<"O5"��|�J��;1K�����|G.�&����E���3-_��x?{҂O���E�R��VA���U��"I��s�ݭu)Յ������͘�� �H�R�q���<���wx�b�����,"�Ř��e�>x�����z)0�AS�}�a�
xW*�HE�V6���j����}�p3�z5ϲ�;_d�����c�\�������t-X���qR�/���*�`i�$�ɢ��d�3�zʮ��+GC�6Àl3�<�G��l��1H)l����ı��l7E�%�#^�RCq�L�EcL�M~9C���Ւ._��>����dc���~�;g�� |��>���b�1�d�+y/zu�!Z@]�E����dh^h8�z�)�F�{��:f�g9;��g pl!l�k�Y]�֚r�J�v�䬏��x�93��ZR��@h������MH�� /�\�,��S�:H�k��[{ث_�κ����c�+eR�HL] �\�eܒ'u��[��:@��:�_fͷ	�A�MR��{�T_��wIDD,%V��sC�����h�~ݭ�Q�1�`Z��AVx��+��hc?#�9�ѱ3#����Ǿ����yPz�Je�Wǳ2�K`��d���r���B�dX@��'k��kɵ���ǎ-v4� �d�X����� 9��9?<��G[:x��<7�=�ZǪ\v����| U�4 y\+pgg9T�Q���Y��B?���PC�r�Ǖfު\'���y��S�,���7�C�����?�ة��?�	��x�%7��B�.5<k����a6��L�fF��b�]0�bq1���\Af����&x�t�/g H�,�x��-@��+�ƚT���zv���G�����nI���m�&�V	I򗫲�GC&��]���JBr�6Մ��U����e�}+E��K�GL6q��|��"7�o60"y��bVA/���,IT"-��Q��X��$I����?"uU�Dj�,��D]�-�_3���R�t�f0w��Em�s?t[�,����qۂ`�+����߁�W�ȷUcO��t��ئ���#�6�}
���H!VQ� �K��n��9'��B./"����(]�i�\�A�� �v�|���4^n���T 8X�,i��#�grmN��\ؗف˫�p飭�6�c30�,s������X� j ň�yB\Gͫ���Bw>Gd#e�X?��.�>U	{5okD���	�����4Β�5�;[��Uңk��X>��ϹV��@	B$1��.�>����Kǅj���7=Sf�A�V|�Ӄl=A��Eq�`�l���L��p��G�Wp��qn^a�5�|>1˚���J��e�
rU�aѿ����9xV.ȴ�!�H$�n��-y���#��{dǰL���:�Xx����B�'C�0�!k��'�����gw��鵳󸵍`h�bm����7C�~��Sd�X��͐V���~�)Po�W]�[]_)h�YJ�>�3�O�U��WG��Л$A.)�<���`^y��L���}(�I�\�i�[���i&�Y����xRo�W�X��*�wa�+���VV;h��32-��$� �3Hf,�-p����]�4n�2��d���d�d0NŇi\-ژ����-���U������>"��y1��T\�C������"���g/S�6V��@�X*,L�'1�y��'LW��:�s8�4�J�z�/�ʶ�G���G����O��	�հO�� � ��Q����L`27��5� 9�F�K_�24Z����/������Ԑ���	�ͥB_���� ��:(7k�})z�!�K�̀��]Q�:��,�����P ܧŤ^��ؠ� N�	�g�Z� v�EA��o�nƭ,��@c��|� {%|*�&0��,8�ػ2xS��R��M���߬���u�K��r�İ��~@n�'�~-,/x��|$�ˊ�x���'���E��R>K������ٕ�Sy�f�`����R��2�d.�ce�ژ	��P�K�<tSw������f7�
u4_�2��)Q�%T`��[}�Z���+I
����'����v��>�҆����/�Pg=B$n�ڡ~\�4�� ���%Z"�w����VL��PU�δI�
� Q��'䃿��ǈXup޲�0�6�/e b{j�<�^���ĺU)��R5�z�b��r���~LnBX��/���v^�D¾���i��*������ЎM�Φ���dU��j���4~�mN=y��e=��m�+Au�Jz�4]�A�Y��c�5}y`1�7�:��v����?�	�Ҏ��{�.�^x$.hh啀��B��	j��^���Ke���fֈѽ׾�J�B�]޸�	���i4����رe��%[._�����)����{�jh��ɮ%uCtv�������	�C�7`�@��D.��[Ŀ��r�ɲS
8��2D�P���׼�V�O���Bh�����"�/��dZdtCF��H,[Z�ʂC�hW.#mf��u�d+4�O�%�PlK����bB����Eӭ�z�#VK�Ҡ��D�˽aMf��)�X2�9�|锑���I25�iyX!q�e��TVߚs31X����j�|Ș�y LM&Rp���^A�~�]��J�8cՕ�(����FD��CLzH�dX~h�pD�ۋ�2%�U�P��x^���O��8/�U����#��lpv�?4ܒ� �[UO��A+ne��yBjYQ�,��,p�I�Y]O�����ԫZhT:RnI�����$V�E��BU�J����
�F	����}VN��p����<���a�'�MM�|��|�����^(���aq��`�bK�pGڸf��l"��̰c6n��-���wZI�""�F��Ħ�N�ۈO+O�u���oe�[k�z��5�S�aPB�-W�'j+]���lb1�_�`Y�ҁXX���������oU<E(	I�7�O.�C����<a���g���U0��l�e!� ������5�<�P�?�mi*���
���G��	a9`4�Cf{.�r�x��~��B[#��n?t$^��ʴ b��1����|�Ȥ=����3X�lA���iqS@ɀ  |ɋ�S0ʣuR��6|,�����b/�4X�8;�g��J��o���n]���AP����8h�-���)IOD�軜6��ךK�A�Ҫ/�mz���۴?����D�l��(P��߻t������j���`Ʌf	K�r��ĳ3s��o,2�R�x�]��'i��<�S�hh�%��������`Ԍ ��H�Ӟ�����O�oBl�7ȱ���l�!6#I���	��b[6.>���J�I��w�cjʤ��Ո�C�=�1Z�j�K���5]���r���|�N�xt��L�1\���Q����Z�+�5[��.맗�r��gN��Nv�S����H�f[!^lC��L΋�!�H�<	�cq����z�D��yzemL�|�unXR���R�K�JR��;�d��=�r�0e�h]����Y�4:��C���T�S��/=��B�M�ރS��п`,��j�s �N���.rZ4�]��(⛪�NvX�c��{��qiKr�V_`�z-w(&t4���)$�T�]e2I�����1^G�D�N�Y[6��*����QE���f�r�?��V�z�r5���z��� J�> ս�C���ڰݳ�;��M���t��(���19_0��d����K#W:��RUg�����M��s����f���2��cS洧���y��.H��ܦT��P`�D�G+��"���������u���YuH_��� �wh�ٲ��g��qʧ
"d�����!�m�G�������ā���	y3�%�D
�/{����OR�����ifp~�[�Tk�5���,ŕ��B�9���|�IeE�aF���]^�j�࿜K�w`o�ݺ��pi��?����Tf+.Fr��eJ�:eHS+�ǁ/DAx��ew5(��{ͳ�U�ڱL�x�q�A�wFU�9�x<�\X�)�LFW4�g�iƝ�uF�$H���d������c����"Y�>�>VX�[��a5�b�7�$ v'D������)�$���|�2��̓�\4f1�^}yy}�I�Cn����t���qD�ۅoQq���4A�Md�p��������d�|u�f�Z�H��q���8����x���y���݌�R��d)`�n	�������4�">�����r��E�;�&E�=��)��~��6�I��\�ъ~a粓ɕg�u#Ghw6i�A�`2�`���ְ�uoä%����g��9��W�����A��1A�z=:���K��;;�T�G2��1*ݔ�m��x������j���6�~�'��#"�]|8V��h���J�)� %w~8&��?mc��QX���|�öf"@�K�`w���N$Y���l����k�����N*"��5)�栀���?��QVJc@�z�B%]v��Z�[����c���9�sBk���xP����b����Y}��V6�wh/�s_��yCK~wGx��c(�C���A`a9���:��Hd�E��(�'�c�"�B��"�[_����DV�&R
��E�̹� ����T�*+��ܧ��eK�u�ȝTnP���R56�ns�s<U�!�{ׯ�@\��
(��"It��#~�����u_�����;ʪ+��4���a3�6kxw� ��U�����"����A�ࢡN4�����e��S��ƹ�U��1�U>]ɄT��l�/�s=��h.���iE��A:���&��Ju�ҝ�p�B�J���?�~p�J���&L���{�Ю'�ň����3x��O�+�h��)u��&�战Xy`n�8���5��In���2�?�r���E�	�$�������{Wܣ��0�Nw�i5��x`�9���`
��q
�v�%��>Q�{�`�p���8��"���g ��<ΆT[���,�F2��_`:d-Nc�;����{I��o�z�}&��&H!k`��TE$��������^�X����}�����Ȗ�+f4�/`��{�y/����
P ¶��,Ϗ���%�)��A(�)9�s��	���HiyͿ�1��1�|Y�Y]����l��O妳�:�_�\sۜ~��!�4xQw�1�����z+9������@�5yXp<�ʽ.������(��4
�OO7.X��Asx:�9<�8�;mV�_I�3�$���'�u�!�֭��Io7q�e�Z���ڴ�K�J���R �FԄ�qP}�tz�ٔA�[M��6Mw�;���T�)�+�[Gx����Ӂ�u�5��.X��N��e������>�ʵ'^�%��	�Uj�]c��9$��):���D�[u����y�@�H��嫴uF�����-�C�Lc���TΔG�y�����:����Y����R�	#dw�`[zu�@�W�+��pH}���3I�e:%�y(%5c��ә�������;2�NW淪�p�M�R��8<ga�^��B!U!�P��c]��]��$��~T��ŁrWO�kEE^;�	�u�x�Ͻ�ʧ����F���P�ea����9��.h���ۦ:7���q�ί��3�873lc�U��AW�2�@A�aJe�.�H�|�O��=
�c��F��֔M��l�<�	��ʷN��V��cV��Z��"�"�ߑ���)"��K|�(�yi��0&��PJ���R>j�nK�{�nj!�ں0�1�p��@򁕗�?�A&Ŀ��T)��i��u�(�p�)��dGƢ��܃���!\������P�v}�����+��T�\e�t�X}�҈.�ٷ?)���I} g*bR;�O!���U$��ɷ�����_��i1�\I���ȣ�~p��N��8zV��t�n�����j ;�uU�$V��_�4%vz�I@
 L vI����Q8����M� �o�7��t�COb�D���a�?���߭.�Я=��4�ʤ���z��#�������cl|�[;�Db?#i�"�Rĵ���`UH���k=��������� ��Q��K��6]ψ��#���3_�;)$��X��Z!�#�\&C�i�Bҽe���>Ѻ�<���?%Dn񍹓+K�u/>�� �&@��&{ޱ�^
#�H/N�E8�(qf�
(�x�q�11��;��t�Q����ũ�ͬP%!i��i ��Y��5,��udNpY�d�\����+=Ɵ��K#��K�)�!�&���/���}��Z���QV�m��pz5݆��0E�g���,�~�0�hVٳL-��?�zlY���5-q�6қ��N���3��a�����z�餓/Sx����b�A�Gd�"�c�VhUU	���Y(}���R0��d}p�K�V��Q_/R���>a���['y�'S�����Aɛ�(�Tgw^∑��;3d<g�Isl��=(��R�J�����=� N6ņ�a3�y�Cp�Y�q����� c" ���$���8�9ޜ�\B^d+�ٌe�\��LP��_1� W<��S�8��_UQZ���Ŝ�_ǢNhJ��ԉ#�{����k2T9k��Q��ir^6��W_U "�<�=� �����8�Cl1�U����_��ɭ � 5-�l���t"��)�H�:3� jd�K�f�	�2��^���8K��4t�Xɰ
�M��(v�� �t6eQٜJ�,����5�~���P�U��ɭ����h�^����d��_İ�u�� �5�OC?j��_d1�?s�������j�W�����ffE�]O�2��ݽH���Ǣ���b4���
_����9��1G����]�w�:6��bq�m���_1���+v�C�4��t�������{8
+��F9X2a�R�ٔ�.�u�[�wҀ_wXnjC"}x��s���+�j�:����J��N��:L橓��pݦi��,"�QP8����tVb`[fev=;���f'�**��Q!.aR�w�F_!�o$�l}R�&�J!������D�b`z���xo�j��,�t�6_4̬��i�A���.k�5����qL��� t�ɡ���E_��Ż\�gɻeYJ�(-������ަ0aj��i�ɯ��n�;�6Fd���Z�'�5��E�a�CÜ%�=��y��K�$�a�_S,�=��<ǗGf�ep2��>^����*b�v?б0�)3��U�	a�}-����
�g�uT�<��w�?ߗ�L��������w�k���8h����������V�QTfsݕO�%yNM�o}��=�S�񈼆AGČW]��k�����Tc6�n�u�;��r��;�{c@^��He�ٷ�,�S.(B��y0��A㐸�z��Vf��$
|��kܣ��\���şd��{��NmJ�$�4���	[ch����?�2~������Dݿ+CC���B8A��Jۖ��͗�[���t�Vmx�Ԑ7W&���|�d�k�^�[�H�V�,�y��-)x�ߪB�t%�W���A«�?�ꡁ��G�0���1H����/�C��G�fBxDf�П������u��-"���p�-&�Y)t��u�y���%!J?���� �)6~�'�f��_�}o�;�=7/\���:O��	&����-�"?)Q�D�t�O��F�1�U���Jh��@�L҃�6��-�'�g���c�+��sܶU�IielJ>�S��la���A:8���l�]���C��dK�n��@y�rg�F+^�A����9:�F���| x��]���xP��-_2�Ы|md�O�;r�/��j�2���`����ޘ?E��Oz��|�H�C�O�g~��}^��/,���������7A�/�H\n}[�q��W�`Jwg�lƄ ����X��e���q{;�Y=�.*[�8����(��9L$N�D��]�i8/.��3D�/Jʁ��T8�P�M��m�M����.����?�����bql�~��{ K-}>g���\:M�� Gl=�mK�{u>4F\�羧�6\xk���[#�K���;�u���£��I�
��$174"������kGU������SyK�?��Pa��"�(�v�\o@�_&�Ɨɴ�����S��J��x��$NR�~�o�E�`��G������
&<̸����p5� �c����[�t%�nS�<�T+%���#�7�(o"!F?�mDְ��4y��F�%1�z��P4�}�ڒ2��3�(cI0�����T����aΪ�f��òJ�����/}�Y�!�0�C�.}����5u��
ċM�nB����h�K�R	��%�E������>))$Owg�;���Q���]�l%�����y��P'�0l��u�:i.(b����8�S5�R�4��߂�|�+���º�?�)%�U��ݫ�q�$���'na�m��k�v�Ũ�nT�.}�kT^�d� ��d��i�I�ћ)j��柩l�,�6s�,vc��BC��:�iߔݜ�|tn��]���-ۇ�Gݱ��O���:��ZI+�͓�5��g�X.�~<9�/P��͓��#�MmY�g,�R��u�L��!���<q}���������=�T�D��x�q�OM^r&[w,�=%N�s�!�r�l�Y=H������jHY�@���6�pC�3�7�d��>�YAwQ#+���>����P\�Q�����pF���k�	�A�hT�)�<ƶ��)	��Wz����y��qi
bK���g�i�w��s��tl��ct��l�]a�������x���3z�%��!t_�_�)a��)x���ȓ�UR��@�p���&��=�d!'s95��f�a聼����8?��i�~i��M�3�\5|C�B�s�{R�u��B=	�esB9Ф$�1S!�\|v�/Siw9)x�<N����A��VDv���-e>(Ŋ�ؖ_��~�	��(�U���ߔ6x�A�ͫ�>}_�|�_����%=ml�&�q�r�d�
���M�D��
�jy�L��5�u'�(o��I&f���'���8�h�i&2�Ø�i�B��*�X
T!�_�{?䜅��:���օ�픰2������s�"�kZ�&�|��2�\�=�_�.������^��zV�
*S}4���ZB�$* G�ړb]������=���̦Lnn��'
XP0��K"'\�Ȧ7U��؎Xr#���<wk��n��
���Lc���o�Jm�f�3G���V�^Y?�]��jc5�ټ�c�E.dj��2����!W�W�!	���72�gj��R� �h�yP\���hؘ�谜5��N4�����v_f<u�Ѻ��L`���|�,>���q�M��^�/�l��s�Β�`V���nveh�_�{�]�P��⾮����w���3�X�J���K�?������-,�~�i��S�ǆy�����ε�į�R�y�I�=;}O&�ZG��H�%��[J��Ԩ��������v�Y^�Y��%wI���iEkP�yX�w^~Z�E�݌���P;_w㘀7���v��>uM��d��
�#��o���T�@��g����FE��ìp�R�s�'K������Q6'��Q8ER���sA��G���?w��۠�|��@�x[�7�b�=��%��s,&� +�v@u�wB7���N ԡ#~��O�����Ij���4s=#2�A&�092��H�<��r�ڶ6 3�?���4�P6���ئ�?f��5ĦBx��/���A*
��̻����<�і�(���/K,�x�V񚔭)2���c������� ��>�_cbs�q+)�1� � ������W��X]�f@Z���kn��QA[+P㠾�̕y����������S�P�^�3������>0�����!
=e���Gh���a��`��g��-w0j-��ނ�Th/`�+L�*� ��֝���H�F�S��ˇ&\ǻEF�*�x\HY�񀊒�)���}ń��w����s��"���"C��Pw�Nf?�$��"G��k���]孬�@�a�&ۯP�v��<�	�Th%%��\h���Ss�R9��>fu��Ǳk�TO�C��ޓ��ln�6�]7��]�ȫ��chb>�N�����I�-�	/�y^$�jA6p�fc�����M
x3a�����6L��͞����$iq}�iHG1�qQ��ؼ�L?PE�I
�9�������f'&�2����A�ľ���q&�O�Ï)��%�$L�~�d�E��
$��D�0mS��9��6����u"�ʎ�u�%����܋499z��x^)�oˑ��ӄ�D_�(��bJ&��L�ׅ�T�t��SO� �+T��̏� �Y�C?��M2�s̪8RXb
J)q����qΟ�A������ˈ�n����g�
r�#��1i��I�~��5E�'��5�>@�T?���FOq���}S p��8���x��_ےΞȪj N<�������[7�x�Ő�`h<z�|"E Z�\�9RB��yE������J�@|E�8���!�y�8PO�3�8��a#� 첤���J��akb���{�Ew��ρv~�+��M@
��p	�G���\
$�`&�0!:G�	�r���V8�6�T�7�ο��L�ЩRF;$�R\8������^���ɧ���DFZ'<�q�5E���EDEO���3�c����`��1#����8�0����>'iE�|���/tc�n���8f����VB2'���D�&嵽��G'�Op�}	���w֝�-=!ǑTOcq��_Oa'Dz�\�}�V��D��^�UaS=�t� �{�>���^�^����8���2���oU��z[L�T�lc�p�C��!��'�`r/���|-y��G��Z� @��`�-��p��޺�K�)"5�2i8Eb`(.sh�赊�b�%�"ؘ<�`E|�w�>���,��ҠӞ�G	��6�&_SX̵,B{{���0�WfR��e�z,N}ta��~8�S]|��}�䕭a_�br�h�W+=�8��)���5,�������i9��� �1�c�4�����V�n#p�&ـY��.�we|�1~W�E���_\[
;FvN4�D�������)#�A���:����Հ���}���5�q�;�������{����L!U.h��(�]��`Ǯ��D�F�N��h 髭δ@�s��O�6ͯi���;���U���\�}��l@�V����Y�57'�'��B�`��Z�5���N@�����9��R���+�V	�u�(0��7~�ө0��Ug������UDs�-�xV�/�R�~��.��3C�K`��X�H"�W飻��U*]a�Nn��y�!=�΍�5{F��CI�f�&��.��E<�Ի�)A,Z~
q	�0�W�Ȑ��ݨ�r��!���U��^��#^}4���(5 %9{ɉ�,�D4v �C	p��f�@�}=~��i�un|���o�2M>�d�6��ǡg{ч	"3�h�?�P4�in����fIv;����?BaJLH~N�����E?�V�Z�'ڟ}�� gCyA��x�9�R�	J�@�&fH�ʅ*m�E�kk�������ƲoQ�N�x����R�n�ʿ�:�׌K-2�X��o�|R��$tʓJ�(@	��=�ɻ��4�������[H͚1�\�;+������k�spq��=`�_�y<x�GsF���D�+������9��g�AW[��~�`�I�(k8jq���������r��˥}7�D�9�����Vs.r�]oqךj��=��gu�H�����E�$���O��i���m���"IC6x��_ڬ92[iY��ܴ+�|cyҎ��$Ǿ����=Ԯ�%	�S�@�EeSF�Ry/9\��6/�7<zUg< ��`C�&�о�e����,s:�0oN�Bs�%��w�0b�z�6D%\�N�|��؂�!
V���WKzv�h{��10U�Xf����{vA� 8)��g�m"ds��{�����$A$�� �죐#04}e8�_�N;��%�r��՝_�g
@3n���(�a6������P����0]�GmY	��l�e��]����3���Jr��T���[J��K/ݡ��p`�g)܊���tN����wŠ�<�P��1�'������M�\KO�ߛ��� E�P�U>�;���Ӵ"�Z��ϠP��$3����1q^49+p���n�+��to9p~���� a<��%��[ˀ4~��FSL��\�t$I�ү�̷�����\X�)���R�ɯ%pu�9�}�!8ENl2�AweO�Y%�糐@��\�߾E7?D���~�&fbe�_���HK�P��<6�j��ʽw��_�� �'�(���92��D��9�JH/���Q��h#$�g�:�0��k�4�x���_�JI�S)�`L^��̰,�xlEm�d�����C�6�N�d|���c�ѷPA�QZ���s� k\)��%ݒ\ԶfQ��h�"�e�s�}���S�-w��*�,!�&�%�V5'�T��WU��:B����S%�7
�UH�����C��=ktδ��`����i�V?�Y1�ӭK��il �g@U���J��k����'eH��j FN��o�oC4L����Pq&���u��#<q�U������R<ʴ�o���0��^'{��iD�`u-�V�5�ǲ�B��ո���d��Ս�^E���H'}�cO�ܝ�קs�L���DW�L���J�7mbZf���Z4��d�Y���a����6OH0�56�����Xeo~U���W��U�櫩޽[��'p�&Y�א[�`>?�i,էç� �u �e#x�B�_B������G���ˏTl��O^B\Q��Y��ԫ6/J<�W��������i�GN�N��f|E\(�^A^2���zH�Y�����'��$���$��{�L}8�8����m��ɜ����~e1)�S]��K�j�7�e7"���=O>�����̰p��,4Fw#�ȇ�J ⌦� eɣQK(ͿM�r$��@9a�k"y&K�H�n�}&.�po2�b��$�W��#)?�ũ��$/�����|�/՟;�)1J�΅Ĕ�����]�CLX�c-��j �8fWx΋0��\4DӭkR�����^;Vv�4����I���;���̂�}M���pA��_
I'���5!�ܰ�>�Dla�EC�[$��L@��p�EA~O�޲;w?4�"a?Cj�B/�&�S8*��l��#ڸa3Sw��Ȇ>9%q���fBH���`���2�u���W��`���v���zۦOkP���L)G\s��RP�.F����,�%�����[G��^B�@��+����]$I%�mA����"D�5��?f���K7�F���!�U˔�11�	�.�;����uk>ʷ2�Ffx����el�5�(ş㏫G��R��]���jb`k^���>�>��g~\�5ҳ��lJG�˞.{vxذS����8�v��]��6H�F9H8Q��.���>���J�@� 2'��-�%�cc!e�c�L[��Ųe�_��[/��z��{�	@f1pɑ|��j��M�O^��'ӒXc3~�(m<��Y�Q1����1�ɯ���K�sfZ�|�y���t!7 �K��(��xlU`�\�DG�����)���&�5F��1Y�g���[T����U3!Y��&��=�E�(�����oI�9�^�'`��9��S����1\#x�WM��X(�9�����_�q7J�.ߒ4�� �ڐ��k��g����F�C����Z��p_��7:=Q|��>��9�=���������Ժ�i���I}�7�1p�///�w���ϖ�y��\(/���CiA����~	sA&�i����Ê�\�f�
XZ����1�ĸpk�c��%{�N(�ʩ�ٞ��r�z3#����! �mZG�j��"&���	a���M|�q;���^�3I|o�kV=�y��wv��d��
�85�h���Q<
�����Ћ*`J�N�6����U1� �Rc���|Z���>�������jj��	j�&ڈ :�E+�8�|�{�\�B��ϗO|��'+S=����`b`�����EPH%)"w1������^�D���?C&p\{f��^����`�tAsu�N��?�u�mf^O�00�=!%��zPa��N)|.�{�"���~������F�4q�c~ӛ�Y)�1��Վ�k��l�)~�<xZ��zYj��} 04�P���CfY0OY
RC��`T �f�7c4:���ԕ{��,��ݡ�:pf�sa���5 @Y?]�C�E���s����욻'�z$n�S���/Юd����R��,[���ʵaDp%��J�R����[����D�-Cl^[���7�?Km����0A��K�MDsƫw���ev���8����-�B�����K~��+ȇF�8�Km�N'�>R��uN{j�I�����ہ+��ƭ���a��]b� �@���%@U�X�ǅ6~�l���g���X3Ct�7��I��|�&��y}{B#�SH6*���jqԠ�b�P%`_���-d�����ZS/�E&��ڌ!��W	�r���>�4�����2��Dm�8�mSoDݤh��(W\���i�c�4���©z����Q�@-[Q�{��/�^|�a��ĝh����"J����.k�@��e�=s&B���"'�7)���M4���9�r(���D�o'+ \:�/jS������zK�6*���>��'�>�����P�pi?���q�|C���(��@��"�R����S����n��#�DE�t�&�_��,���'�n�������z�|
r�Cw�}*A�La�n�Zw�Kɕ�=��TOl� e?����m�AJ� �����$#8��/_+�]�!f��k�����z���s�0^ �t�Ж��O�HbO�Q�YtU�IN/��^3��G�@
��(b�6������|�S���T�Zf�dY��h�H-��y�7�N֥���5�%&�s�|7��<����b,
�$��<5VK&�d:���w���\: �0uju7��UጸA{�?����]�U�/4���%]����9��"*�{���O���.�����W/Ş6|Q�&���`
1{q��΁������Z��h/nE���Q���M��5���M�������������/�YIT���m�46d��J���)ʡ-�[��3ϊb�9�9Q�
	����f`��?'�~�2A=Ոح���jVgq�v�?Y���z�{7J�90��\(����m�rS�֤c��ZC��vJ�)b��S�Z����eRm���&��������v׿I11Tz��p���y�����=�ݣ+}���0X�1�kf�白j���:�Hzb�8'	��fZ���=:�Ϲ�l�:B��+����M	e���w�S�y���朘2��P�q��؍��OYӼf5oJq�iy�6���$�Ow��S���	Թ>���Oـ�H(ҟo\J�-P-�N���{ +?���������#AE������>�1��{
R�;��D2! ,PA�ɠɩ�%$�)Bc�����i�U����Q�rw��n#���=�u�bvW��uG�O)��4S�Ca9ѷw)t��A9�\%�o.����4�#/�!���%v�Bp:�	�'?�l����j�|n�.�<(\Ժ_$>��e/B�6B��Jl5��1�Џ#$��g�Ω;�lE� l�T�X`�����)��BNR�n/���2��!�����;�K4�������,o>(j���*�oeð6Pg1��$ŏ�?������7����{9�9K�˞��Y�)z\^l��Q��P�!j�2^��Al�
Ю헶$і�}��������c{FG'� ���@՜�e�C�����GE��"*[��`T,*��%|_c����^ք�����7M��O�-]k���4�����W����!Z�F��D�^�T�~Oŵ�4��Re��ʌ7hc!�c�w�K�z�$*���#�Y������_��jvy|�˻a&E$&�X0�<ߟ�qxsG�4nhS�z�\ȩ��E�l>����K$�]�)�5��t��BuX�]�e	q���`��ϋ�:����U�����Oi�����Sy��O,��7q��8r����өn��	�=y,���fB��ؠ��kA�5	�`��t6 ��2�R�4���&�3Y��5W�qTo:=Pj���k�y�E]ޠV\�����~K���֏����=�؛���E�+@ {�f�Ռ)y�Ў�߸�����}r�Q�.����w�V��׸���}�3����(�7L��� `{�(�|��5h�@k,2}/A{䉀�T�P���G!��Y�tr3��zê�[g{��L��n�$+\��X�Y�0���hk	��+\Y�y�O����u�s�'Ԫc`P�<�m4�����:ف�"�+��/�E���Ǒ_�Q�}��}�wP�7mm
��O��Cu�q������`)4lj"����YI^��n0l]�Zt0��F�i N>�.)��/�/���-���-�t��pVo/=�4O/�l���Ο�a�h�4R#��e�v���G�5O�F��.DG�ln9��S����}]ϴ�{��aG��)���B��o���#�[`��,��D1���Nf��AY�lp|k�2"\�ό�S��+�����m0��x��F���t��:�<�U�'V@5��a��l�$�G|�n ���q�=?�.��3_y����˓�%f5
�/��8}���y#%�@O���I{4Xj�m���m�8xRl��	��W S���מ��q���]�w�r��.�2��;ݳսA�7�d|��J��s/�_�=<~�3���%jw�8W�3M�Y3F>�B���w��oFME6{���kvH�6*��Mv����u�����S���4�Q�|���y�&����H��I�ũ\g��X	Uoxn�r���tK�`Dv��w����24Ѭ��r�'2���j��o�I'?�;u|��9����%]�oԫ��g��� 9�2���A��0�����Z�\��V�2������T�gq8���Y� �A���K�����:a� -���YDf�����5��8���,�7���}$M�{~�V��Vs2b�m��5����u�B���#��<��g�.���$�Ϲ�d
�K�a<�{@�f���R�XM��g������r�~�vN_c(%�h[��v>��U��.z[Tc��ӏ�t�E�Y�����̇��v���>\0E��in��g	v�֪V ��F�W���a����˴¥C���9AC�E1w�c�������cćIW�����85�G6F�]Q �<��ށ&&�̖4P�IϬ�����=;���X���1aNL��K������EL=�rK���$b<�V���j��Z�aG�N�d��?��N��|Y��k�_�U�L\�]����u��J��C1H��3�!̉�Ĭ����[
��Yn4�v��j"�h�m��������Z9T;�}.��}�������0�bU�&}��3�,M&;�{!)�UT=8��N���5CB����)*�V.��~���b�ŧЦ��_�C�M���N�<8��ԕ>�wxjv�w��T��~�x��?ӤB�^t���䃀����X:�:�5�mo����3Q���j�RI�koڕ�aߛ_9�6�Ri=d��O��k>&�0Ӓ��NI-�Z��=��!a3��J���'Wm��G��L�����阭���@~�_Wծ��p�:<�a2�$�u�&��d7�&W6�O�j:�e�R��U�$<,�ЂL̥a�$�<�_�s҄B�JV�=E�-�p��f��1ž�{PKt�l�p�B�u�1�I�M�Z�Ɲ۱���q�(��e:��^�Z� �KƮ>+����z��	8I6O�]WI8�|�20���N����5�1[�&j�J����0��
�չr�O�	��w���r���ޝ���O�˫#vz�p��@P��(���a�E�v���p5ʔ�v�'��_��z����-Q_E��e�ىg1��GA�}������� ��%̓\��F⇋3�ޠ)���6�h�y/9!���,_�j��{�TQz7��_����F�I�(%�HJ�+�D��&��y.�fp\�n
���7³�\���w��K�O&�6�s��w�
+Uzq�j��5&Q�rHN8HalL�� ��|9��zv�H9��(�KJZ��(���"��bQ�V��F�~�R~���X�T�!m N����	�`R��B}R	���!�#z����};�ۈ���&]�U������ڸ�R���U�-�5ԇX�.e~3�ٞ�+��F4R��/��/4�#�9���� 3�0*�T}¬c�e_@zh�ԋ�Z���C߲��x�V�q����j-�C]w{�{�7W�i��|��杼�#�ʄ���)>�)��C\�>	���"�4�{�t�[J;��Edi��j%U��u�	�q���iw�<�	�J�}0KU��M�u{ �cU/6����t��l=��I%�P��ߞ�{J�#]�;�Kw���,�R���:^�t
>}Ă��"����׶J�ˁ��H&�~�T!�4hmz���+�B�o}������5����b�!#[��E�w���-UM��?\c�K�gyE�.�s��FF�K�dUV�
i�(,���E�β)~�|S��&|RSD9�]k�ZШ���ڒ�2��׶ه@߽}�� �r�I�Q���13�e�3S��v�ȸu��gZb�)Z-g�L�1�v��ES����8�&�_���:Z^QF�/��4�&��i�S
KxÁ	�yn�� T
\j)��qI�D;�5qJ�
�{
��݂�iqډ<zq�0'r�)]��9�R2����n|��BܠKJ4��2��Ĺ��{��A?�E��;��"�T�D|�ۇ>RA/�8�.�v� ?8�`ͭ���z��G��mЁ��X-�IW���J�/$������R�f�7M$6&pډ��$��1�{ŘD�hC`Nn:��Τ��%���fu���>�h��bv|ފ�����L�'���@�p�}�p����5�zk��D�T���Dt
��{���lxŐe� ����^I7&?�Z<�^&x1CW5� l[6�.��>�`Ǜ�Ʊƒ��Y���ŢkZj5�-��L�-k�y�����2 ��
�����m	��j�)�b1���{j�:�>騧_QZ����gc���r�ޕ��2�'�y������(R�-*���-ǲ)�-QU�x�(�C^Ov�Fql�j6֑˯e6hY3��R��)���/~ �t�D5����	r��F��XK\��D������.�V�������ot7Z�I��d�g�d�Ĺ|Z:�Q�/,u>�5��^��#���f,�M?{�S��km'|`L��#��ܞ<�}�ӹO0ɥ���q�VH_�:Y��L�
��%s0MӉ�w�\��Z�>��>�E�Q�%cD�����F��
tT�S��?P{ˮ�� ؈T����N�^�i'xk��Ƙ�M��<U2R)�L��*f���Y�&4���� ������s��M���U��f�F��|)f<&��X�uN�oH��ݼ_˝����e�q���5�0��d���v�OL����4@�c��I�L{JPnD�G碠[�;��&��z-[^�&�i��h��|��}��9�����N2P"f�nb඿��"<Oy�ͻ�/D������S3�S �1�z4�4�Iy[���C.���&�T��<�8�HcLm��x@���Hᓠ��)�HpW�W��A5�����P'�&s��o��j��ob��1�G�}�4Q�h���R�� �)��?l�mJ�5�p��	0�����A��yU��,��P9����[WC��CpU��5�W|�
�cV���"0��Jc+-I#q�R��8لk��6����P��*�%�w�V�e[�`JN��Ӹw),LtiR+�%Ԩ���K�@S#�|�-E��4�����-S�4Ti��,�Ñ��Qv>�m?,�JlJb������4ԦΧ~b�0Գ�������>���X���R˒�=O��*��:Q��G�/�W��s��2�@��g�׃��P}Bz�����{�_�LM�B��)� �z�X���c`�������?�Ň���'c]���AD���6���B���<���"�]��[v*�P�f8)z���VࡌIwۅX�U n=�Fv�l�G�%M�G����b���n��egq|�-��Z�n��O�T�>�*�O��aO^"C�µEr��My�K�f�|3Ţ����kuy���%Ɓt�\@OFI�>4F?೅���.�RT������I}��W����;��^HZW����ţ�o��ٝ6��naT�g����;8��dT�V�F�����)�k�sb��p_��2���'{O�����W7śrv9�7��V^5����=QF�$�)�0k���ũ�r��·䋶�� �\|� �T,��P0���s6�VU�����A��rV�m�2�N�˞:P%���Ʌ��{��H��#-���V��;>��t�69���Ŏ�aج㲑WH�22����
��q�O�eů�).�[(�l��֍�THN5��P*��QɮD-4Ȱq��(ˊ#y�`�${6��˴��P,�a�$�nDx�&�jLf5$�f$,���ZK�+�+-��l�<�M�:�����h���C�HY���"�dB?�A���{:s��1[�V{��*�k`���RQ[c�����(�w�!�e����m��˜�{{!ژq��Bmw���^{���$ ������[U~fB<���R�m��қxk^����� ���	�r(j����a��W�'�-6�3�&R��E{�.�����h�P����<����}��wk%���E����'����9G8����C���W%���Ј�Pe %{�M�}�����R�ϊݳ���N��h�����У=�=#�ٻ3��Kbz�࡚S����>�?}�9T�{j�M�3��N�QɆ��'/ܾA3��� "ؗ}T�ů*�v
x��`.a����P���mc�UUϑ�;�=8Q]c\J��Sf�u��k��Q��TE�1�r�>�����*�G[)e���#��к��x�/�x:���M�K�`Q�<�w?���YɈ�w�r�MU�c����qsB�}�L'C�}�����fzyz:}(H�V�� ���.>�?��܃*��LC����N������2G����S��b->�>�}jJ�#�0(�{��@�WC�$�:}+���/`��IGh�j )��`pD��D!�Y���&�d�;b�Q�;!�4*�L����#��mHt,��<T���f]������|1����q�|�y��}����dR��R��
��+��O����������t���2��a���x?^�)��|��&�=h�39&4�0f���(�b���ӎ8����s���S����}����63%�\H�kז�z��0�U��[��G�2�_"x����Xit��RQ�y��M>׌诶s��ҎZ�k�oso˄�'�l�В�U�/&$0�P�th�|�Df�M�h�ُ �B���L����տ���tT	��-�$��~���d��O��f�7�x�y3:���mOY�Y�"G1p+�W�G�E����TZ��MhES�l�����:�Ű��y1չi|�p��z`�?�䆢�S᫠d� �^R�D�6g�'����Ak��ʈ}۲H�_Pw�}??<|���
��t^��@a�v���H�!"%�a�һw�m�������΃��;���ƋA� #I�ՎF�!#��+�][���V�P�4�áY>���$,�2���`���R��
z@�S����\ �P�����"a��RWrh���ˉ����z�=&2��oe��w��2@�l����  �B
n�:�G��W7;g���l��^(����٢Z�q]]�Phw#�n/�]�l{JQ�乧��4c,�1V��G�
��'`���}dv0��o�d��-�RvG�ZI�.s�,j��FE��-�����C��I�&+�-��j&�>]���~Y�:�s(�wZ4�Ѹ�U/bct�8(�P����n�do�wz1��m��?��g�D��PxY7�v��휈���v�--����\��3�T���<��!��Ͳ{�҃�2�_�#'8�ߐ��촬OmD�=ú́��DT
u��>G����O����ۛ�N��Ş���'���Q�݃*��C �P�Щ�Dv������ڔ8pso���U�y&�+��݁%|�)��a�X���־}7=�,}��]Ԍ[tx�(hև����!Q;�!�C�{�m��^�^�������P�P�m�Q�;2��1V
`�x3�~D迳�q35�.��xL7���xQ�J�(7��*�&}���^����z��%׬� �ӥ���h�������b#(T鄼�>���Xx�=��jn.+�P}��Ĕ��a]O��KԀ���'�v\��ߛ�j�sa�UR/?�J=�,��d�̤�_-al6v����r�3��B1���ִ�c�DcH�J�����Ĩ��03�ղ�ɵL��݄i�R+��UV�_��n�y"0��H`�Jદ� �T� E�HB��W����U��n�d`p{N���7 jJA �F�=��.%^S]��R��-e7{�F�����!j��ҝ.�ݝ`����	i�[���w��2�%j]e[��X���8�1W