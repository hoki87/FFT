��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n����x>��r�_��S��7s�6J�t���/9���0Q�W����=b}T�-�uZ��)B=%�&�8|hnv��F�3�����V�}�ѧ4�B@F�jP �\��P�ο�����]��,p��2n�q?&���mGx�{#��@�9�_���nʠ� ��p��pJ�kA�9ӻJsk4���,�
9�y��w�e,��cS;����4P'7:O���w?�Y�o�������LǼ�l��Z%J�]�/�u7�(l	���l�\�Cod;��'<>��]��W'&���2���d_ʹ�r��c,] 8�t��s\�.�1m@E�w�t��a�걷�D�V4@�2���ʿX�����ڧ{:}�,�n�{&(}���:�s�!�4r]��HX�DI��7�ͫn� �X���#��E?����7PX�E���0�8���k��������X��p�����g� 4�>�K�e"�6Z��X2Ț]Y�s7S����d�0qod�{��E	���Q��|��-��=�*ޫ�bM���ҥ!�d�.�K�7��3�h�����bu�c+9ɓ1�!���֬D��CR�ayT�J�Z��4+� N�35��zW������a9XV�_�������d�X~���7���_|ԛj}�0��y�?�7��m��3W')�������N<���Ō=�Yf>+@��P�*<k��=rfj7p��
e/R:M>���Vŷ��q�)�%k�j���|	4K�O��K^����FYk�+M�v3�~�fU��
�'%�L���k4�m�tZ4��hv\��]3_���0!d���f·i@���1�d�+���{Y�?��"�86)�3�R~��`�l��Y�s�4��;N��0"u,p�������42����g�i��h\����4���X�^F�"�����mX(�����4]�����t;T�Ad_z���%��|5�?m�#�7�TU�����{�ۤw(ʊ�F>=��мX�d�%��b�he��{�_�b��v�.�����6�ծе\�nv��R�ԐR�#Y�HZob��X��m�O(Σ�J�	�OM{%�;
���@��'���9WҬh�_J@%^)/t��R�mȐw��-�>HW�Ɍh�"��Y2�8��v�jꓣGu����iB2�gM��=�F]�V�Y�K2��#0%�����E�ؔ�>v���#Z�σ�4�I�9={I?�g�*�o� ��n.���"����t
���>?�?&�=d0���᠐�����D��f�D�z6�;B�x�1��!x^��y��z�sk0�E&P}���޵��^?_Eݴf�ܟ{[1���&�S
�����,ǀӞ���Rǎ������X�i)T�k0rJ�A�~�� ��\�H�=j�E�:����4�����[LYk��*��5�s�Sz�*TZK�Uiј������K@���恑�#�d�h(]�\��� &;�X���ٺ���`\��6�^������M`��c�Y���(4�]KI������렗�*D�������|���.�d ���=@yc�+�%���Vk���.�~쨑�g���~��k�{hDU\7��ok�|P�8�b����"^�����u�~���f��}}DR��C��aC�\�`���ߠ����]�d�@�Z�������Y��I\t����{�,0�EǏ���V�g7�z~�g��-G��\�>��O���"��J
^�M&*���������F��>�H�Y%���d?�u>���EoUA��� ~��J�1�y��&�"?�yF��I;�\m�o���9K!ܿhs����_�#+�=�&�e�V��)���9*���^Xԃp`���rb��Zg ��1�S�`@p��Ӻ�C�X�Tw���?�+3ϵV^���7dPe��"��a'q�#�
��Є�{��{�hSOp4�rt�=�X��V��8�c=Ge)����~|����(9�Iۢ�"�;_��iP�S�̂B!��1������~�+�֟Ѭ�"�F�ئf4����,���v}q�og-��L�<x���5�{~�N�����8a9r}��դ�^S���K����2$m���|�û��8�з���h��H��K���D�G�E��Ncr�ZQ�u���ƭ%�G@d񈛛�&Bc�>�u���hb�;Xsq0����ĝK���O���8Ip��`�N��E)�)�����E���GI�`0���Q%�4��r��������2�~F0u�+0��z@Ѣ�)�5]�V�@�|��iԖ�Ppl�A����|hyC��xv�7Y�u�W\�v%���bmRŮK�#+�֞apXj!��m�ZX�������Rv׏ظ]S��:�cz�*�h�0�t5
u�'�9��	���7e�z�lP�>��S[����7N)>)!Yt� �biʮza!��B�>�̙�R: j���W]I�丛��n��Ng\��4�H�5?Υ�(e�N:���}���yzC���8�=�n&1L�c���Y�W�fz<U�u{�:���2��a��!O�݅\9Bi��������!��qv�S�ӱ*��������P�����{� �"�<��ޥ�k�:M3�Ɩ}R��)�)I�K1Aw@�t������e��|�:��۷��!ꃭ�0R>��F���*�̛O��QuIe�Q|��}si���V���$Rn,Iz|Y.9f�zM��B��{�J�y�bZ���&Xz�������
������?ʖ7|ТnCr4{��U��Qc�����x�Ԯ#���Ⱦ�7*z\����x`.�iϵ�7I;�g0��[E`�zΆľ�]� �<#��V�܇�"5cl�h2_�a�J�d�A�AZc�T���+����r��ӛ��(�e��o���1Q�� �.���V��V+��R�el��\���tX����s��=�h{�٥#4j,1����4o��h!�x�C��䩢�d$���"��ە6�lO���L�[i2t�Xn������2�kM ��޴��EDd�q���cb�L�̼���y&~���ԊI�p�fK��ܧ����7�<�����G\�H�w7�E_�n����u���4eo��3�X��QSUC��>��_���W&�'tހk6���f��c5��̇ة����/'!٫N&��z8��uX��a!D��ҭ׎�4���k�(�E �/1C��>���w��%̅��_�6�Xutpu�>?Q���d�P��s�Q2`�M�Z���S��[����i�_��i,��E�{���5NC�uV�5`��R��2�nа��cO�#��'8MS���r��֚�e-�8���J�kh�s�f�Nw-����*Ħ�X,̔��{���#Mm�q�,B,fD��h佞�����/~��w%(o7��l1������0h�ZOU�</�(Yrkb�e��XA�@$������t��^�����Y��aC��| P$�Ϋ-a`���Y�Ь�Tx�<���� ��Zj9���V��P�G��-� ��Q���!�[U$Tl�eg��Q�#�A ��R �=�+m�Q�^��D-�"�,��eIZ����h�a4�[���f��e��Y�8fوy��� �$�4&X�|MI�p-������"������vAZ�*=HND�;�Y���4��b�rS� ����
\�l��k��S��C���� %������y)r�[�XA�X%�&
��0;Q��γ�s!�7���u���Q;Qd|F�l�����	� _kωѸ<�:za�*�7��PZDύ������4�V	���Z$���Z4�'������+���<Q�m*^L�w���m":U:���@U_�K���C�w37�%�������D}�����Yp�FF7S$��zȦ���w��B[<Zf�p������Z-�u���yP���=���Y����`��S�f�1uHc7�H_T�����x۾�9����1��h/�.B$�ULbt��6�ۀ�tş&V�&����W@��j�s�r����إ�N��=�k��^�f=I���j��C�qS��W��7d�UZ��/΂���W9�.9��y�^�7��E-8�Wa!�l:��)[,����zƁ� �����i��(ƣ���9�d�=���f�h\Z�AfLVa˄��4N8xem�܄?���ҟ��מi�;��²�ɇ���[L{J[��@9 ���7�Ԣ�h����>��L�'���ёeJ
ͫ�'d�M7(�1��V�:���1�bɿ�4j�v	�/j�����9�F��%�vi2�d^m�mg6�J�-�i˸ZԻ���L�&�h��3��g��E�C+�jr(�v�ó��c�����bXwR��+�,V��n�?��q�|�crk켰M��d��w�_~j�0��ʙ����k�cB쭮���]]�=)��-��<>��s��M%�2�M�G��íg��\<	&�<��/K��U�E��:�XIj��ƖV�L��vFyQ�$ �i��q�+�CK��vvu�u���������!�<Akǩ��p���ή����yk����6򴿵��xAȦ/�����FB���G����kt��_���VV��oIx����ud�e�ʇ�>�4���s��#�_���tl�?K��{j/*�JXGW�ؑ�c�z�n>s獹�˯��3��>xv�ǜ@�,��5B��S�5K�q`�-8]fD�MԢ���k���&~&w�^���z>rD�C����efD!J 7���0�g���{���&�����?�y��3���}�ƺ]�;�Q��2ĩ<��N6�q�=8�+���w`I4�����΃	��{�<��!�b;6������D|SZ6����?M\*�c�B�#-4U�G��^D�!��آz�ᣎ}"I��]�:;���%� ���]��K��Pﱛ��z�Љ�0%C�G�TN���=�u���Y����^��5-\�H�x:�*!�K.�����!���6�^XN���p���q��z�Py`.f8�#��f�ů���}�P�����
�e/���SWG��M�F	ǘ��� ��|�/k�!�ZME`��w?@�XƟǁt)`���mD�FU�z����ẟ��8�u��i��8M�>7��8f�Q���%�ָQD�Ռ�zPPKT���W����7�7�h8����]OK�19��p��Ɣ8%p�ަ4i߲	5����"�|�%���Z���慿3GY'���v�RR�$�)�L��"u��9��,���a���r�ђ}�V��M�wK������W���|�{ �`��
��U�(R�M1��#�}\���W	�}%s�O(����k�TAb��Gg$�2� �8K�鴏�-�!�����o�`�#�?�81�$>U�����T0k��1!FOy����O#�i30�`u�0b�����)�o.����0N��-��k�09�T�8eG�7�1C����,��Hs[Q�;�woG��y߄�� �=ˍǙ��#(�#���`Q�2k���0��*�����F���g<���](�7��L���W]:�1��8���.n�>��dL1k�^�����~�)c�"�&A剏����c���[L(o�{�IZ�j�aݏX��f���m�$	�N�јH7�U�
�l�t����o�s��'��8G����2a0ݿto�V������*�8~�S�hגƟ�����*[��7Q���~������.ˁkv��fcU���+�8�ꋝL�=�j�{�v��&v�Z�"2[���=�����mp8z��r�g����z��8�v�����k�~U_(�jZ���k�wV��y�( ��П_�����#)or��e�n%�>y�sa�	G I�H��\��]P�Q.jߏ�њ�[�Q}��z�袒:]#�g�����oU���2,�!�i���_'8��}����wMW�}�-dl؇E�=�}[")�.t��c��l*����A=wY1��즪8� FY?��C��%1jj^��@�r�6����l�($ؘ*�\T�-�K���e�,Xe��#��N�&v��w(Ҭ�ħ��o�\�}!'iկ���@*b{>�	�5oQ�Y[b�6��~	s�)��mt6��V~O(e�w���*ǚ�}I|$���*d�}�=\9�IKX�*�= �f����4�\[�����-49F
��v����uC�(	
�l�l.i���PH���!;�k�����O�?aCY?�>��y'B������k�>�|���G�KI���O��'��i�M��IͼOd Eg�H�+c�����7:=ҵ�q�[L4��m(�U��P�R���X�ֵ����`B�D(�+�D�\=iL�fO��N�$�ԛB��_A�}����֐�E�<�#�\p�}8X��8Hg�p�W���·�2��˛����yӟW��dB7�x�oe���g���#f���03��6�c�D
��w�w���m�r�@(Ү5��Vbx$qY�tY����K�?�=te5e4�i��_W�h �}ș��>%�zsa �J0�D��[����2}�����?:E��A��Y=Qcs�5���q��u+�8��J1j��I������1sȦ3(�0c��m�=�K���ȳ�q����r�u?�Sh��|�>�W�+1�@kT]�m��Ftz�d�����Ƣ���U�OI'�P�|=g[�U�F�h[uu��EO�hV��P�ɘ�U�#���ș2�m���)���5a�J���	몤�ۀ_4D1��4*NeaB��3>X�j��X
�t�0������8���Js�s��/���H���-���dK�i�Z�Eb:ޢ�4����t\�D�r2�N����$�%�*''{E����Ձ�/P������E�y�����%*�R�Y�~?*��R�#:��뢘����6Aԕ�W�v�e�Qe�h�đ�/i�E�`SVCoٹA���@���@��������YV^{�sPY�������KK����,7�R�b"����#�J�� ��|�n\W��=���[�-�r̀}�7���3���F�����I�i�p�v�K�	/PعS��*��U�
s��M �clX��1'��ὕ��^�����+�M��D���W���]Z��֒��,4�rO��vϽz�B�w��5'���%V�0�3����C����b�g�Jtg)�!��5Ӈ,fQB(�Rl�4Z��a U����F=�%��ZJx��b��M""zS2��M .n"c�S�B{��G��5�	�LF��'����O=��ױꇫ�a �.rvq�Q�Jl����~�jOe7؇~�h?Y��A�$����EfbF�&��h��i���Te����>]c6��<��&<�.�9�?^
��#�Ξ��Fz� o(�w�6�"�u�J�u_�:��<�%�[�?2�}޹�,"����$�:!c���>��H0h�Aѡ��X���7
�m�~j`��ZF��]Y�iG���X�I�8���,a��56"��X�����_Ʌ(d:������P����;>�2HAU3��t;R��#^d�n�r�X*�����L&����)�\X�[��w|�������t;����Ƴ�Ƙ����U�%�tp���q��'v<����5������0���R��4ǷY��>�.sHV�/5&)lB!��0"���T2�ծ^�4�z����r_�/u�ȴ���|�pHI�-�������C��|�K��!�K [���!�+n\@�+�)�4�*߯�|������pB��f�}FCJ�����%��X���L�!�������{Z@�C�����p��ް�;I��/U$O�N?�0TK��Lpz�eRڍ!��Z�rXpUy�2,��!Ƌ��ǯ5�2U����k�|u����~_F�z
w�Ŀm*�!w�3Kƀ�=`�l���H.A��|�T���z]VSc�#��(�pu��(��<��0��q^�s5��b�z�`#��%W� ��t��ݕbC"w���z�UEe^%:�-%Q�W�k
8�/�آ!?�>`� 3�>>����Z�P�'�!^��u��ߚ�{�#�&K�mBm�$�/8�=�<�R���T���U�6�[m,�"^#�V\��U�jG},V\7V@�����Y���o�@���]��&�ȲB�~['
�����r>��LV�����j��:��V�n�o7����س�x肞�A ��i� 4�Ṣ5?γٌ#�\r�Kr����{� +.�ԕ\ļ�L2VH�����K,ʌ����C�k���UJ��^�k��2�-{�b	5��AeTׂ����b^C��zX�n���0�u"��[�\��1�����>I[������[���J�f�	���8K�Ȧ���=�NV��bq`��Eb���5~JQ��֞�Z��+��v�����G�1��^3(I��9�&rH����s7��G�6��l�|8 �OR3���>B
���6_3L0D��Y�J��u�.�؜}J���G"~�S�$�2~����(������:$�>��K��u%n�n%�	��b���8^�gg�v;}}��(�7�.v�z�L|h��ҵ&QLIrVs���J���#ϔ�z	���$`q��!�����7Չ���A�X�_�&G����������q]���J6d�p)0�YS�yr�R p�~���!�d\�rZ���@���g|U�Z92b���Uk%�x��(�jܟJ�U&j��4����&Qg����M�ʸ�IK��l7�w�q�3�5��;߇2U�����]$�7;b�o�g4�~�Oa
���eWƶ����2�)�%p���w˻犒�J���n�P�&�w�?CF�/.pD=UbBx7�B��m��X��\��b��٥���ٯ�<փ���n͎�	�����>�@鱫���7D�j�up"%����w���1Oh���'��雯³э�^փfL��0�g���U��1X|5��끓�f0p�D�]��CB�pٷ��y�K3��8.%V	||�上�pj���>�q�BNzś��q�U}=9P�6E����l�'�M\�Iš��8���u�Q���k-�����[�T���;zV�'��Q�n�	_�#d��6g����vkp�����ݭda�7�A{�!F���/�l[ge�̶J?>xbI�ڻ�)�d����ƥZ�d�-M��}-��4싟H}���xŴ ��U[g����7p���!��sy:?�L�|�ʢ<��M��{�T�L,0�*��_��j���"'�m���f�P[�����W�<��T�׌O~)�t���dޖ� �đ���-pɈ�)sz/��/�E|��15��hf��Ρ��^D�9ԴZ2��f����J�f3���n���J��"��<�x�=�C�e�a���Vz�W�zHX�nB ?���:~�s-q�m%��hW[hK���/�����>��Ga��N�}�l�V�fm���X����LK�c.ܷݯ�T�"8�)�I��z�'qO��(��Sm(wzd��6U~x���-f�v|�)�°�X������8_N�a��,*�W8���d69l�@1P�S���f���{�AB)D��=�G�S��Ҳ"B��|]a��S��B��,���V��`�ZC���}Ԙ
�~�x�
r�Bz �ӡ�=Ss�:dc&?���=帳����d��]K�lF����g�YH��b�u�	�P�����#w�Ƕ�1�%�/���Ð#�.j��/�g�T��k�N@m�����H��:I?���	0�IvI���V��F��H�^G~�:��X�P�k�N��PL�uW�6:����[�]bMp��.o��;�|v��}���?JS�Ya��;F�9�D����jܠ����NQ���9G�.���$!��!:�[>#�c�ܤ9�m>��C���@������ё��J�~�u�5�(�'u�����˾1��C��L���s)� ��V����c:i��hg���`r-���X�����3��F�9��'*�ɑa�Ϯ��J�!���ڷæ�<���%w����e��yQ��O�-�q�G������~�j��!�FuM�h���~�~���?)d�g"��R=|C�2f��D��1��S�Q��U&]���L���=^�3�����;��-y���4�:F�E�`��7�x���A����;Y���յ��qw�q7Q��
?�w�BU2�p�K4�Ռ �.�k*��<������o���J�#y���@Ҙ缇��w$&Q$X�]��V�y�,�1H߃�.�MLx��#K�Z��_Bk}��ݝ�J0>�j��Dc��V��� ��u*=#)�jb��4�������-boHF����k_�eA�t��*6��<gh�w"�����Q�GE�ǫ��K�t![�$z2rH	Vé�
 �@`r��ע�寮m���h�g�P6Y������G7�ʹ��(��Kӕ����ޠ�.3�qt�k�����1+�e�w/Msp����J�s����rj}:k�4�Q�:Ȇh���Nn���e�2{u13K5On��eo�`r�����Eq�kXtϴ���a@������Aׇ��ḅR�/��+���"c3��)�Ey�Ga�n�6�(����[�1'1!���ԛ಺b�n�h�����h1	ӡ�l-$#�=��(�m/���:M�$� ���TK��E2�R���݊�����S�N�ۮ�r¥���O�:Ҳs�~a�҂m`$��2�+m���j{�d;� ^�:�ܥKa��>Nن�3;j��|(Ac���˶�~�w�_�Qi� ���|�B��p��ӭ�P���KcU��i7&�Jߝ쉚��v8&�g����gKW���a��Y�Y�8A4T8�Df����*�u5���4��>Ί����B��a_�����݉T����%p�3M��rzDLF���p���ܤ7��峣y����22�y�oC������B縀���b���#8sWr����4P��ϹE>�jBo�J w-�Ż�m1;[-uD��o�ݤ��[�U����S_-�g�%�!ӹ�lޘ������+'b{P��@̤�2l]��*_),�	�X�����y�!	��]��Ǯ�	fg�R�3<�n�q�[� �i5�c=���v�QIYoj�n���
1������?�lB4�b�,�#��YP$�����{���I��mR3�:'���tt3��h$�~E��Ӻ~waE�ߨ��&Ә��Y��9Gbpr�u�`���w2���@@9��9���}-ʛ���T�e�x��)!��wռ���lY3�v���7R	4/��a���p�	�f~5�'b\�} �A%BK
�JY���A �*�ڃ	1&ﱆ�z�0�mW	�5q�34$;���C(�w� �A�Bd�yO�Y�>ξ���J>$Ǵ��VJ�R�oQ��u"���\�H�t�|�����0���= $�����`�-����r*CSټDJ`]2�Ҙ3\�a�h�zM)9�[�7@�2�Kf�����y5��EyLȺ���$��#��o򝹎�ؽW�C�8�!=V�);�O��.\5��Ha-+�i .K$�O�n�nx��:8�%��;6襆>��g�����р6z�
�����{H�� 8Q󤀙��%�h�?�����	L����(,x
�%��.�/�����h:���<I.-ّ$O��D	I�~E��u�i�5T�����
2(�[�KB�"�ku�7���f�S��o�M�nh��ʽ�1{?X]Lz��8��:̈́\<dw�{��-[t��nB#F�JOa�����T��\�0�&�4;dWT$C]����8^'F�ur
��"и�"Z<X�T%x�l������vb�U����E�C�-A�L�S��ep�
�4��^}_G���:��y�nAEh2���������"�KZA��T�O�ā��@�A�3l ٘\<����L}��L��u�:��Wc�ХSǑ��N�U�^�c/��2���m�fd�^�
������ıX��;���@Ý5*D�f�$�}�څ��_��c���m7���(�GEQ�?>�R�&bu2�d�tu�9(M�:��,P<P7" e�ﰧ?�ԟ;	��82����Z���� h]��>j+�#0��K(���cm�����JF/��5�_�ϯ���ܺ�[�	���~ �t�u+�" AآǑ~�\����W��k7�64%U�J�evc�):ϑv�j�s�Μ�E �+
�v��Aㄱ$�?��j�Z�A�c��6���_��7?�~����[AP��?Z�iY�8�r���t�E-V�k�K��"UU,7���G�������t�Չ��������1�8��V�I��O�`�qk�Lw�ၝ��~�Ƨ*
K���������D~��⍭��������g���Ltv�M;���78M�]�в����l��7�G��.�'������S+CՆ�`W�e�{��A�S/�/���vJ�k�����f瀉�?t[���L������gNZ&���Añ�w2s��|���+�BW��_#�/��6���YeL>�-.�c�d�)\b[{�D�3Y�:�4���EI��Щq���z>lL;%�,�;�v(y<�[G���iYޫ��x��.��b`�am���%;�@	�Nt�%�o�&��Baq�����
8B]Rx{d���s�	Lص9�����v�D+���+��{�:rsCsI��߲��V�� �����~d��_�qk���Tإ�?}�4�~�+��3�|�r�Axw�y���{�P�?2
wԪ7�{+��&�O����rQ[*A	ƍ�:k�ޑ-f�ݟC��v��KɦW�u��d�'47W$>�ߣW���'���R$����{R�2�R�tA�|�wk�S��v��8>*K9�3������jS*ټ�~)Ga��Lۿ�����q��|�
g�wT���obc��t�i=�YL7�I�J=�[�`JY�p�auk�\Z������VK�G����sGy�MO��������0��y�=l!�H�*������#u���/k4��"L��r��@g�ȸο��"].f}̪�_/�1D����tԉ��tn�}:��W}�{���e5�h�D�-'�o�K�g�94.�۱�2�u����KSWJ�o跽���5�aE�Ɉ�9�2|�N!�L�@%�Rˋu��x굤,KtA��l�Uz��Ww�r��xFto�)&�D>p�f��D=��!B����������o��clMY#GnH)9KH���ڇd5rW����W{�Ш�|�M�W�S*.^�Ng	�?#��bJ�����8�;Ok�O�`8�e���hwKCRǄۨ�n}+��6���ƶ7v��� ח`��#�R�M:���~z�DQ��� ��w>=����}ww"�|{�6\�=z尦��#�R�T��.1���a��R!.��D�����ՠq���~�XC���'R�d�o�^����� ��9��Θkd?WC��*^�
�i�\!������PFk�� ��9b2}�������Y�Fb�a�,W�a�!�
�j?��b;L �K3�����Iu�)�E#3�ȃ�q�[��<(��v8w��E��8�l��Ƨ?��ʴ�W�"CN�m���*�*����93�b�H^�e+r�eפb/�q��r�2�#*�}��:V�..���a��WE\�q��{�e$�+σ��:��7�`}$��Z�fE↕����o�(�R��K;�U"���l�}X�_�p�]E�h��$�*S������As�T��s�%� ���pGy5%6t����Z���f���X�����8u�u��&�h�p� �R�2m�^�rvSD�r��t�}hEl������>XH�y�e0yg�@�4l����3��~X���FW������B����^��[} >��Ҷ7���� ��Ȓ�%L$4��bY���e��9�9�=~iVC^o+ae�ޓ�2֝t�._H	��v2��b�ş9#ɚ4w���R��7z�,�`��¶j�ԩ�1<I�s�� ^�n��S���jtʞ;6���c`���8
Ə/`0�t ]��黀o<u���ق�Hw�?�'���~��� ��Pi*��`68�/��*��K�.�1��|��y �0,U�)7�|���W�������6���{�K$O���m�'��U8�>l�IO��L�IBe��^i8|���j��d˲������d��?(N��i4&:�uv��n�������������Z�D��_�zH#���U�����Qui�u��� ��Z�bzSkH|%Ie��A��`{�#~����k��2��w���._��� 4y�7b����Xpԝ�1$ǔx��!9��B��WV_����aĀz�T��}wc0����25P�����Ww��e�%t��
�`G��3?K��bP|�'�;�����37�NW���`���C�J�e�A���L���TS�_/ˮ/0����G �w-a�;wG=8E���kz�31���3��5�a��oɦJ>N�wv�������m@N�	&ϫb�V�qH ����aW|bn��?U^��=����q�--bO�ZJ䇠jfP�]�A2����8�?2W����z,xoi�~j�3W�4F�g��yk�#��ZCXސLfR��)T���˖�:��Bey~�E2����,�h���2?���NB(G��*�rGOYȍ�~�7<�����
�n�Nw�f��s��#y�pGd�?{k��Dl'i)��d�{���֍@�40~ڊ���R+���x�!�����.�M°�[���<�C���Yړ2�� �8�O�>x���:q+��Tvc�Ҝ�Uc��)�E(2k֖̆���M�ĖD����z5��)����+�2Oثj��߯o����U����s�o=w8衂�z�w�֋�=�.�gD��T���*�%�ۡ>���>z�F��ޒ�(�` ���FV����{!x�.x�����Cx�ԇ*����ީ2�@���Qe7����j���xn�Tg+!��p#��-(
孥#H-a�����Ԏ�"����ε�H�$@�ҥ���츴�6��C�s��!@��h��kn�y�q�}��nu�(��y����e`�4���3F�]/��ߣ��Z�ݞ �6j�5�7�K�2П��wп�zrF�JmF�E�ETߙ�9+M�Cg�f�0��� ���H�ݐ�:��oæ>2�w�`��y�'�Gݸ��y�����S�nB�L��M��;�����ܝ�'�Kܵ�竮�]���$V6>��M�dy�:�	d�a)����w�����|�cy4��x�#��2���������Ĵ(���Մ�6jv�ϯ��u�v4��um�{7߿�[�"���MV�5�p�S$q��wO�sK��1)��R`CƆ�y�M̘l�ol��Q�95#ud�� `��t���Mj*���2(A}Ax�j�>@�t�q�^!�@&0C�8dW��v������._�ܯ|Gx26~ۯQ���t (Y�����8�����t�8}T��0�Ԋ֯#����(H�@�@��IaB�noY C�4�$�����`K��	k���W�;�3Z�Ҳ<���.j�������*���x@�)��X��CNr=0�>	�ȥ8�\I-�������$�5�.En��k�XxW{8��E|5�j�'�Vf 0�8�γaa�i+�$����Slق�&*p�W\���X��ʳ�V�,����bs�l�2�Q�JÈJD��'Ȯ�&9�c.�e�V���1�v�Ad:`�_�E>�b(�X���Ɠ�HK#��1/����Cz��^�~:��ޮ%�1�:۝��ʃ���6M԰�?��.:9�ͤ_�	'��S��N1��������7fW��aQ�����+s @~�C��4C{�L�
C6�e�d�r C�����};�BxR�"�P��n���0E���={N����U���XXT��(�yK	����+�ʗf�,`ʓ��+�L��U$ytg��#&w�"r�'�>�=xL+����rc��@%.��l���H��3m����KC�r)�6���G�0< _s���j���=��9�-�:��@�M��L��������b�0�5�1(��'��% Ɲ���zҙ-Y&�ҧ|�"87kϣ�̹�����G�Q*J�č������j3�K&�Qe��ǦѰ|���V=��'X�y�j+�S��V��m����?8/}ZѪ�7\�_��y;C!a��4���I���= ����@HM	{�|�\��r���p�UF)D��c�H%Km��Ӱ;$������6�=�fY�~�P"H�Dx65�i�\;�
�4�g\�Q�� H�ϬֱU��5
Z��ވ��r�������r�*��K�!��/["���9v��+l�&	75� �G;4�GB&���_������Dh��:6<v_ e���Т�G�'ϐCW���֓�����U~��柢�lB�N� N!HXs���A���eF��7{e���[�ks�XKЛ���&<\��h���
=�J�/sˊT�z�-�X�ZvEf׫C���N3D���CX|` )��J�|׌'�Ǜ�nY�]}4K׿q�2_�Cs;���z��N��XR�� g:!�n�A�648=��dF�� C��q�l~}"C�E�"t�'5.��o����ߦ�V#�/��h���}<o��ۋa�|,{E.  �[HPZӾ���d��A�7sO��~h�u3�C]��qPO+� J�<�~�3��!�k;�F&�7{�2-��n�?,�EG"e;C�¿����|��[�=P�QT�����2h:������_��~�I�b�?V��;�F���5xVsf�ԩ��'�NO	l���t��gJ��Ҩ�R$K<�*�1;ɐ��;�s,�F@�M�y�ݔb4�:ڜw_�G�=W@(�����\*�����	�����w�-×L�(�j�b�8ܯed�ub�ܪ�4�?Y���/�^�n;M8X+���p��~%tn�?�pN_N�7�O&]<��i����A��]�2��,���IWl�I��Pz�v4�����`'��{���f\�9�F�u�&��(z��ѓ!p�6������p0����˗�-��i
��,ظ;���[پ��Y�HSt��:G_��+��`d.g������Z����J�(�?һ���7t2��;䅌��hA��y��"��V%pt��~���>4!����W�=�#OJp�/�;��2Q�"槐\J���#�[�z"�#Glhlg	F���'W~ێrX�o)\��U1���Et�+,`K��ݥ1�aϽ]:@����z��b�>�L��w��A|�R����s��FAu!�G���ej�q �4W�"��R[������5(��X�h�=�b���$8&��γgV-am���#f�	%w�Z`4���x��%7W��q���1t�./ �v��>��>V�qC���.��e~�i�mMi ��*X�+���J�I�c��P�W�<#���p"�t�lFItx��������\��~�0RE�vA��3:�s�
�?�(ҋNB�X&�nc�eK�I�"��|�:�zrk�R��)��9����#�bz�K��}�O�w����2Q^�[����f��nW4�E3���uZ�Hw�	�l��"{�i7߈ߒ�x���~�K�8�;e��v/fw�\�4�/HQ����N���r3��B�EWӳ�1`.5�l>YE��9�0t]�:��iD�ၥ�%I�17x�����4��G<��2���@//�!b��Ix��
�b���y~�~�+��c<R��j�n�q	��GShn�~i��3D 	C˶�jޒg������[e�q5Ҕ��Jm��-�����wԪ5F�4�%�����k�x˺Ш�vk�}��v{���$$Ol�b�o��[�"}��{:��x�6IS'��g������������s[j��L*/
���ƺί �T�547کB��dd�Bǧ����W���Z�]�n����\���0�zLz1�������H�j-��2~�;к+�g23��j������_Q��2�r^y}@UŎ��RL�/7�dIÝ��uHd}���v,�.CyAs�y�x1)09������p��0w.�t��
��ã`h��.x�o'l�r��� ��PZ�VU����OD�������h(b �q��f��7�upV�n>9��A/��d|f��ލ8�����J7�q��~?�bS��(������<*��z�@wMH�ö��P��Q��af��Wٹ:�
��vQ-�5�	 [�'���w� Rc��dB���� �d9'�'���
}��'�m��OF �f����F�5��#����4�֜�S2ź뉯Y�@�w~���ˍ��d��8�6'$d��dA��`�UW��*8�N�ǐ�H�=Y�)��h�ˁ���a��,�vTU�&汧�(C��ߥ�0줋O�Q��۞U�O�X�˖���Ų~ؠ/՝Z��K��u�'Q8��J��	�&�A��w��\| ��(:J����~�ˉ-B��=̀��x�v��mEqs�~�lhb��Atr��f���]�e/�sH�cT��K���ze����m�����s�WQ�O�r9jH(�U�]�^�o8t�{:+��vh���&k��f�<!uH��HЊQ�%&�V�c�3ϒM������w �K���;���x�W�S�mg�И�}q����c8�/4�����N(��X�D⭻J�����PGb�?�Sk؂m�%������;?]���U �$��]�35±^B�Шж����B�gf ����3#��j]`C���	bZ�H5�Bd�Vv�]��[���:�;��9�i`x�A�?jB	��ʡ �
!Zc:a!��p������!��r?D��3�"DB- 6�dk}q��f3d�W� �����x��	v�x�a_���P��D���|%���ԌH�Ȓ���� �k�q"�u���ħ3]w��I�-/��"�8_�z��ϴ,�B/4X�:�t[Y�DK&�Uy��ـ�^�-ߠaC$l�y�&bv��)��=G�p1Xk��~L%�d�K��P��/�n��iڮr�y�	G^�a�ǳ�P�B�!n�1nvQ-���뚲��XʮtN�gf����ɜ/�^3$I��#���r���=��������r�~M	��eڭ2?(����D%yL�E��[���X��c�6����Wma%�=��
���%��*��а���r�
��Z
�� ���{�|�[X��kb@<�'&lF�p���G����d��{r�'���ƵǛ�0w<P뢻:
t8ک���5c�>���S\�g1����ӵ
8S��VK�*̌�R�#`��+ �M�9��f׎���̤	��	<g��do�<��a)����N��P+����B���Y�``���1�Ь����m�D��O�~
����w-�ɶ�* ��䅞bɝ4y��ܳ��tw}�1.a��N��Y�y=�t_~�A:��=E�p�a%(Qm��Gw�n�p�- �kt�΋T ���YG����;��S~�t�x��n����s���4�ua�[���e��6�[TĴ������fv��M���>��L�-����@�j�a?��(!&)eU�a���G 'N�T�i�Ë�����D��|�љ�\�tHd��'�b{�WĖ�LٶF`p�}ᥛ�v��j?-��j�G��Ѿ
gX%�l%`u�}�$)�?��#Z��^"���/P�/7���T�{[�޺vy��0	�E�3��P[�%���>�H�"�>k��mU�2�;�Ǜ��٘)W-^�Vj����t6魍T)��ypK�xIEk���*l�3X�1���3׺�)T^���G$��L�����˱%�~���j��4�u���K'2����4�;�뀋�뺪��+b����C7߁����@6�8PK��ƣ"�-.K5
� 8�;0'�P�``9��k�L�/�&���^/Tv�����3g�Q:&����>�xli���NR�,������h]��ٟt��b�j�|�q+�}Qi����.:o�n���$�1�O���'��6Yes�
��g޹����Bj
�U7ɹeߪ�!�k�)ݥL!oSF�1�������
�js<!���h+�>�@����1�g��3�_^�Q�.٪���!09]u����^���!�1�C���-NYD��b�R�ƫ��i'naߚ	�������l7�W�W��|H8N�*n�V09�,�ad��j0�,#F�x�oVk�\�7)Jx(a�K:{���`�㳫� ��U_�w�澌�Q�p?���cj�AO�@[2��x*k�ޅh�������wѷ�.W$�Xx�'ŝPE]�cy��E`��1y���l)\.�CƇ~bS��2\mE��|��� ?~|�3��`��6g6:�?K_u�?�C�W?Ӕ�ƌ���>��|߹�:��5�w(��K�M����Q���4e��RL���p�?����HhY]0�������M�\�)\��Fg(tBN�Z�F�.4&q��(H%�W�����q/��!��H���ЌN"]&�rH�
�A��rn��<�F�����#�$�T<�5G��?ɒ����p��/��&±��{ŀ
ݤ��x�(V����yɈ���s�?����b	k̎^b�h%�(�oDr�[ʁ��gAey����c�0�~�ۙK��& 3��8��|#�b�{�"��䵵�ב�`ѯ��ۗ���~6��u����N�Czgٸ}�R3ǧd��� ��5��ـ�@սN&Z�}n�Ԅ�n)wm,(��5P��7��k��jG{�Д��`N�����:(4��6htX�I(���@�2�0���\Ʌ8�NT'D|���{��<̹���L�T�[qϝx_���y�*1[[��P1fA��B�&�/��nep�銘Z��2��A����"��Q4�#�:V����KO����NTl<��i���ޒ/rti6�i�,�p��#s�B/#p �u�Z�G����2�VH]T0��Yg�%"�k# �腡"��<��Y,fd�7bz�����'P�/����N�]*�iꔩ.�T�����!��ve`N��Y��
��PU��\u�`�J� <��N~��G�y[������J��Y�V
���@Z����Ђ�<m%�M=�����?V�x�\���ݦ+6/.r'×����"�!����{��0�k��$?ʵzPU[���X `�oZ�JU&5Z���X+�5�xeb4A�$%z34��=[��LS�T2��|�3�U``������t�&��u�½�c��I����k�\�u�4�����<aP�O�W�"tq��+�%��ƛ�� 1�pi�#~�8ֳ����e�Ϛ�Ug���b%�Ds;���;ܿ�8x����oo��<��<5%0�2�%�Q ^�!^6ȶ��j�DBL(T��P���k�:rF]K��ͼ�1��)�W�n2��N�e���ڳ��L�s`���'����FѲ��'zz��iBN A���1o�B���}kſ/L�Q��O��s;��"0����g ơFN �p:=��zY���-Ą2���/��)������&v4�w����n�O�F���f���+�q��9�kG{�S�� ��u���`�+�_[l:�;LuL�͡���Al>6;a[z��;b��A�I+,�{·�c%��U/��R�@�#��K���<��[����gaа/z�bIX�Cgt�+o�p{e *n��F��Ċ�Tě��W�F�]�P�U��Z���Y������S�s���ܻ�Xz,��-RB�Q�^�Mh�_�J�BH�{�&C��S��@�Q_��TB��2��p��[P��YI���Sf��g�K�w�|
������߲�u|	�J�<P��
�?\vMI(C2��}�N��� ��EJ�E���M�w;p/�a{7���1²��`{�(V]4𜛟�/�-��-���+���(�f\͐��f���( [�m���f���}�iK�&�`5��U��znP/�a��>�dV@&d�˅nxib)
�,��ɍ.f�ko�ֻ�W;�<�K�7��KD9�#�qS���GTZ� J����u�4nُNy(7n�F�q��b���K#��8`�eoP�V����T���>�����;�~��:er�a�Q�X�Hx�x���I^ jE�Է���]{q�,�ؘD����!e5Ӧfi�9zn�� �Αy�|��F��N�� �N4{�\�ݯ���N�$�@������M�pYDRGo��D���X�K�7N��N�kT ����␩�O�i��c��=o-F��W�L׳0�e_i�Z	�Yş�.\��/��2�$�O;�i�Iכn_aI�e411�<Mcb�*M�qM��p�i3����3rF8��D�qҟ_Vn�OpV��8�D���F@����6�)�M}F�:���㐗m�����y7�ׁ�N�DrFK�M�KLfo�`��:/lLYq9pԏ�d�tL�<rYe��U�;(�R��DoH��Uwd&���ئ3u��v��d.���(P��H\��(��h@���hw��J�����yNt�xN��˒���2�T��v.&$n�Df:RpI���N9m�c�m@�9��6�/��#��B˦�����E$Ӕ�)?����j_)�aݥ�X����C�Y*	:˄w���D s
�E"Py	WA���T���ue�ϑL>k���.���w>>#��2	�L���E}��`��No�oY-�����xF_+��/�4pZ{'�:Z׵Ek٭6��p/f�O;]����	ʝ�H��){v�0�P��-�����|n�{N�xO<%G��֓�?<�3�Eq'܍fY�ZR0ܥ�_�-E~�M)�9��v*�\y(R/R 9�e��\A�!�n������π%/4�R{	b�;�6���.xJ��Z��[QҢR�^UmL��k��A��	���v`����s�;Z`�����e��ѿơ���¬���L��Ȣ��j�ڢ���X�i��hni��M�Ǧ�e?%���s�f>�dx\{}x���$�P[�Lv��Z�gh��7˼�ƶ��(N�.�'���V!�q���BzE�=��ڱ�^ݱ�����4w;��%GNؕ�!6����2��3��u��e��`��(�x#e�W�'sf+��䨝��L��'�-4ρ7���$ ���2y���v����!�L�m�1���RR����jn��eĳ�����H��~ۆ��l<V��ݺ։Ѧ���k6��5�;��Ϣ�6��N�5*;.Ƿ�]-زU��O����>"M.`��$���^�?�X]α6ǉq�g���ߌ�Jp9Z�Η���̫$�������1r<M>Nӱ�o9#L,�R�A��n'�LF�mz1o�w0J*3T��J�N0�pF͔����^��Y�Q�^&{jp;[�X93��\�D�����ķU ���ԍc�\�PƠB�4��A�!h�0& ����`������02\��e�~:���m�)<	�Ǯ֡/�z�
��DZz�S�
A�|����n�f�_�b\�^�PЀz�RTb�*�`���<����#��I��R��ҤL19� '�XyI�kh��Қ�U�"��B{	�"����|�pV9���e1"�k��ޔ=<�'�p�|w���֩�@,�[�-4�c{�tv?��}�p�`>J%�1�?�h� �ĳ���-�S���G���*�4^���3ҽ'T~-ʊ9H���0ݕm�Y�i�����u �M;݈Ι�Κ�}%��$i�$)�|�����:�i,i^�1��|L��˦?#���`�q�":��'����-dA4pm"z���O�[)q�k������w��M"�<~��BV1�b-5��ٿ�k�Sn7+��I�Y�pUT���~.�Z㞍^tk�a�o<k��,X�����j�(�r�����2���v����u��ʣ��.��[\���W:[��L4��f����
I�ۜOv����MK���[�oL��ʞWރ�a:�,ʚ�h��0х����|�z�%PI,v�� SVu��E)6+��!�R���|��[�;/�%��x��j�[�Ѥ
�'^!#����#K
�D������&Rd���a���}�G���c��SH�@S�&�l�ԋ����7��=<9�訶H�A1m�qՍw�#�TA_`��QDn�(t�m?�;>��E�.݃R��̑�B3�km�2F�HN<^H}wA�-�r`��W6���aǧݵ7b��@1��A�;	��d̜P�J���������:��m�4��Ǎm�Q� 0�Kw���ͫZ�WZ�|&di�0�%D�ʟ���:���3|�w�Օ�A #���I���tW�r�NY�j^7=n�$>M=�\���-ӵ���=yZ�^�r�S��ĩ����D&�oh����Jj�(��v�֣,a�.ZО+�m�����	����}�K�	��;l��_��uI�luf`���@��y-��t���K0(��`�>���c��V�S�o��5�dJv3��/��d��_&��	�A��CC:o7�Y�2����&m�c�xր�HĿ����2"`�\�Q����	��8��&���"v��Q#q�(����<�	z�:���^#i R�R��^nt���ɪ2��ȣ$��V�0�*��X?c�{4�"�u�0c��b�L7�F���K��â�QV�y�ܴ�D̃p��M3����0Kv����3K�����y믝�zm��6XG�Ğ��a�΍���W]Y�y���٭�\*>��"l���U�.5�_�2�F��3��k-X1�V^d�gr����|�[ۄg=�@���Ω<"�KMF�.!b#׋̗��s�A��*��c�k���	.��||�mx��&`�PU+e&�Ԩ�v�Vʸ.��m��{�wב�z]8�)I���m?M�5�N��t�F��;�Y>䨎Jl~�S9�����R���f��Sn�(S䚂w�+�I�*�NR�;C�f����iʨ٨/���n��&R(/�|��E�ƅY�t�J�t�K��/�����q_|'������ι-���+UQCfol'J�E#��ȓ�ó���:c��vOm"H(�P'|S��w���z_ �Q9X���-m����ț���_c�몖R��Y�'�+%_���g��d"W:{'ty�x,�߈,*�+8��l����*G၇\1ː�ϱ��y����#xM�}bzg�7[:%^��d�B������~���ϻ�E�XNxlD�{Y/3|�ȗ}�`�@�HV��B�dǁ����@��r����b��$3����ڶ;]A�&������;ϡ��V|Jx��\��{�em�q�����jI�i����9��2����N��)/��R�/؃�ܓ����*�l�+K�s�=Z��Ti#� �~���B�;�ޡ+^������"z���N˛2H��f.��wU�_8e��8˿��h�V�T��m�|0���,�`�.�)[�T�l�S�q�d�A=t�-e_�%�X�����l���/V_��@~��B�/����+���B��{��Tx�z�\�
�4�ݻ�t�b~G�>���
�ˇ`����,�ĕ�-7�95zz���v9e?��彯�\����~n髓{&����x���S��~�{)LM�º܅�g�ΨΦ����Ar,h�0d��;��}S�j�<e��凰��2��n���Khk?`�O@14�&����+��,*v�N����kmH��f�O@Ѕ�b�2��� ��]�#��}VK�c����嬐w*��.o?ThUl�!�s���qo��2�,�@�<l9MZ$�߳kU�ؒG�g�=,"��1��D7��C�a�<���e�_�t2Q��MTjk�O�^V5�=x^٥i\اS��V�E;�O�V3W�Zi�[���'4o#梳�8��i��`V�M\A��N�#������e� ��3d���*a�L���)L��[Wר�_Q���9�d��'=Q��$�%7���Uޖ^|.*n�fN&!���X��jSH.�������@�A= I�8 qY�e;�<i�7�H�J� �,a<����3؛�����.��n�t���8{�VܖP�����t���K�4���)u;ud��)[�I&��aM���Mi5�C��CK�����|�ȅ�0I 
S4���7��\���;���y���(���m��֭Q\j�L����D�O�B��X���zm�A����ؾ4NkD���qcZ�YO��Y0��� ��ʗ�2Nj�^�� .��{V���j����ؑ+�C�M�[U�����e7Yp$��O]�Hm�����!��R`Pz"�qI��|��UZ ��Stv�vP�T\�u(x�5��suXK'��ɰ���4`$�����k��{�	PF^T�<���+�#NƱ�P��Q�VLb���?�`ã'ikG7�!�䑐����Ş�[�y�%u�-�dd�����ߊ�*����ǫ�j7�b5j<X0���g�]�T@��uC���)�U�Qh Q�V�O�	�~[%��/���^�Љ��C��ϗ&cW9�sVV߀D���K à�?f��ISJ�E��?�?ؼI�J���?��ΈoA���ʙNسE24NC_�Y�,�k�L	����J 	DUl+����� �tԺXI]9F���G��c�n����I��K��;}�ΰ��]�gno���g�P�>!���@kdy�P3�����w�>&�>��
y�@zmşWŖ����cZ� f�����ĥ���{��y���&�J���ֳ*Qʱ�6��>zm	��{&��)����p�H(GG��YGcg���~�����A,d��;�pF�cyq�'ȶ���au�w?9���[?ׇB� ��
�;濅B]���v'�g����J�w`$�����O�oS(Y�L�Y�iÀ����� i�O��Qy�X(��߼,�k)��������h�:�⺃,&���p�(v�'�:���j=��������n����6�u�H�ܤT��C{yR�e�,��p����[!���kZ���ds���pHȶxS�
�¾��@^"美\-7���<XL��E{|Jyd$�Y7�s9TE�d��BF���ܢq�q=���=s�
�@�v~#y�����R�k���m�^t�o�5v&=|0��Y����X�%}:͌� -�3�D�V]��|Y���$U�%w�4��@���K"�fyL�6X�مT�Ɲյ<P��O���Iv3��o��R�0������z�r��B=r��:�x��(�`h��T6��(@4�黚V�R#"~%�=��ܲG��Q@b���=b���es��OR�����#xd1��x� %���b��j�T^���B�_w�@���WaQʴ��kc���+��ƅ8�{ɂp������p&�1*Ιp�\�X���řJ�i�ϩE���|ݑV�<���IW3�;¨��0]��eu�㣜	ҧ#��'���J��H�{�&��ߘ��	�*�fB�xv	����Ɂ��\޵��E8�9������6���y	��9�8s��������Óh�yw걷b�@C�����r ��85�e��24�cL�Oܚ��cz����"cߒY�|o��?��V���^��	+C� 梾��y�
"|�E2:@V!4��Am��� Z���l��4.�2
C���y<�E���Y�a����aT���8�F��e��D&�	�se����Q�8�`��y�����S8�ӡ�>�ҍ�����Ĭ��곙�1t'�ܞ.�Nϖ�n���Db�˕�P�E\lj>��
�b�VBH�u�:��B �)ג��� �C��"�ɥV����J?�+�/}�^B�ء�r��e�7'`�)�"�����$\��~�K���U~(bpnc;��DW�`Ӏ�`�)�th	'Y\�ut���$`3��
����߷R)�0�2(e��.j�T#�q8ŘM�mb�6
�gxf���)�8�h��3��`�|���v� ���!���/����q�SEY�o�H�D��7�����1��f��U�s�f����Z�/o�e����Lq�a�pY�ϟ9�u&V��9|��#�ٓJ�^��U�)�{	��L=R�g��
�:+�Lp�y�n�\��v�Py���ӊg�4{�t7���S�w��k���PT�җ�����gbD�E~(�Ta$�DDDv���0+	��N�G��s���A�2~�+3+��?J��|��Ŏ�[;X=jv����ՊU��樧n��^!b�70�x�V8��.m�]�H����i�x�O�u�|_�W_��z��gԮMd�{��S �F8W<��"B��#����R�nsUl�����ʖ�� ��S���R	��T���_Mprf;�r��l���lRj�<n����GE��p̌��� G��H����e�Չ44�c���{�F.��r+�֩]��@d����.��H3"�Աd1�B�VL�Bw��.N�@c�z�U�0��~�r�za9��*�yt]� ,ӀHd	����@�裄�_q�B�]}�$ؐ�4����-@�DWZ�}B���R�������=�[8�f�� ������X�Շ�P?Q(,ӄ�$�dR�+W�Gg۬|X-Ka���+��fā�tJ7#B�2w�.}:Ϯ'j<���e	����L��X�w��S�1��{c�3�݋��>>�0����f��Gj����3ֶ8�l]<�P���|�;�i��U�d(�;J����b.���/����+��e(Ws5��{h�T��A���*��iTd(����@�!`�H,(u�$��<� ��'T��޵]����r��(&�č�I�ץH6 �B��֎\%*'.Y�	>͕U�h�=r�,����z�r�'e�[����ߵv�ZWoc�X��}�F ��42{�(wY�{0���<|e���1��4ӠaX�����Qo�U�,S:t]N?�lgO��c�ZT���Bx�����k�[��?��"7��K�4W �yR_����v�sau�όטȩc�t�1���6_�4�C�o@�p��r�g�|��z�����F��:�!a�	�R�]ё��Mngys�E��А���rL�������ƀ՘�K��p���Hw��զ��k;Ć��Pnj�{�$u0�rh�Ƀ��{\����֔X�3��^B�Tէ��A>& �6�IO%ms,dG���f`���D���<� D��%a��V��M��X��)��;y�8'kH|�Q�g ����[�]ZE:Y�#�����z�a～I�y{�(��Y%N��"1�Ww',8�����h�Q�,U[�v�m��ٮ7R/�������,-����KS��N�Þ1S3�H9���Y�'� ��ݎ��:E�;�u�+�|}�Ϫ���lD�HXuE*=���TA7��?��륂�v�� ���XF#/LE��2���m�rCˇ�i�z���Z�膢�z��m(~��c�b���Ϗ22�yY��D�	����>u�l�+.���Q�B��� ��9���3-i��q+'�&�)uP���v:�W��5����#"L�ע�E`j�Z	�d���f��i���ԸA1<���<��i�W�(�x����l�E��">h���`�j���{,'(	�>w��!���-o���Ԍ֌]=h�[�E6,YiM�*]օ���N�{'Ą����&Ѯ?�HB�*�	�-�s�P"4����mhG���\?X�GΝ<^M�����fP��ʏB$u4q{$���{����Q
�PP��C�$QaRͫG���*�N�Hu�Kڭ.�K*w�����I#��߿�d� x�J�F*	/0�3~��ڳO�a���͑X� ���������Z&���1.���%x8��B	��.��g�%^��*������R�{lX������w- �VRh.ƀ�����< ���?�O��G@82�|,*�G�p��]dc�w��0uJ�O(����`[+�P���<����œ�g�ssPhRED�����xKOc������Y��00�,9��� ߣ��gLF��3����f��t/
/������u���$"�<��r��K��@f@�}���Fҹ��eⷤ���>`��8T�#��c����X=&��2����������no?�yR�+�CFbe�\���R�M��V�Y�Gr��Nd�Xiha����N]�N�B��{���1�"~0�7��[���;8ɳ&�g�lk��3�/�Y��B��ˁ�ӓ˚��j6;�)`��HX<gĸ�E���h�x���6�*O���s���B ��=�ܹ:�!X�U닰�hA�"X�/�Zg�t�q�bu���PV������Y�Ѻ���;ƖgD�Q60�i�l�6M���J|�{�g���Z���펀ݕ���
���[�=?!k�U|%{'��k��ŊW��冀\թ,�Fձ�%�ʹ
���=/�L� �B<B:�E_�u�*Uם8EQk�M��])�lh�Wr�޲!�j�Fi����Cq?&D����lI����Ҩ�~Kb�S�E_��,S?e��i��{^�S�|!)\�|�U��e�߆��^*&������D�p
��>�9a9�Ȅ ��TJ�S���3��ͥ�d
C�D7�ȋ3`m$*����;�n1������/\�l��/n��ziHLW��Eo_�,R�g��[���X{9Y6;%��2r�m����c��̳ۛ٨���iv*�-QU
yH#�)i���H}�����l�5b8D&�A�H�k5Ȉ�=Sz{���vuq=�]���.'��E�`�5����̜��cÎ4�6�]�"M��o9:赫(@��I)�B�� ����"���px��4��� �<���r���ftF����k2%���p$a׮� Qԩ 4�|�"EWm�r3�e*lz�f�wyP��پ�����klY�X�vj��I`�9a�4Z+� �/��R�u���&�S���M�&@��������f��b�Gd���q�
����{���J�� ��H��!��k4��HO1a��Ϥ�l�lD�'h�ؤ��k:�����,��.���Zd��{"Z���(��4P3���NP�O���J=fْJ�=T�|����:�^'��, �5u�W_c`W�i"c�Orpӏ�fY�B!9̺X�ߒPm��� ��P��V��Sٽ�=cO���W�uޭ��I�M�0�W���u�4'����wr�+E����nXe���U�(�rD��	� f�6�UF�����:�S2/��p!Y�j� �J�dn��q��5Wȏ�_#2��	���xy`�f���΋���>p�h��>�:!��0Tږ� ���J
Ն��z�k�r�c݃�x���B;�{,�{�	�u.�;G�[�:�[J�+��n����-���p�a��irhO�E�#�����;B���a��)���Q
D7��3�QA{Y���n�?lz�L�)��Mtq�\�rO���0�11pˬtj���ZR��E��w/b2����Nh�z<eE��"���V����}��FJ���a�7��p���F(
y����#��8њ�>L����D�	`�a�!��畮�{D�	�P$j��1"���3�U{�3|�6�ͳ3�$��\Uף5p?�obd�$/��P1�Qw?�U��O���?��>+�xc�[Dv�=��*�p�N��W�L��{��#?�{Vn�"&���T̑g�Cl�]����ΈS���m���� \\=�2%(���v�e2n���nN�J5�GF�b�zk0�S&��h��P�s3IğV�3����{��rk_%8�G���M@p���.R��ˁ��9D����y"�h?�����:6�)E֪[(�Yk��8�$B��f���K�v��oq@Č6"�j���Rt�g�!�!�Ue��2ܡG���g��� >�
.�����՛�fb&�\e��*ɻ09����k��շ��y�P7%��<�S>a�淧�ϐi�@��p6�j�[��]N��lt$�غ?ٯ|��[#m{Y�h���Od֖����� �)%p�j���W9�v��]M��ϖrJN�@n`��菜���� ��m ��r�����&�U��z".�`b�;��5�4֮�CG���~`+�f�d�o�=ё"�\�K��F��T�,}L��_�]O�z���G�M�6<D@$ПQ��R�ߕ/��e�t�w]<�)9>n&q�֕Q��B�|���^�	�nRwnǮ��,��@��<�hUc<܅�Đ��Ɣ�r�/@�n�=�Zwu��:��>ce��~�~',B�E���Q48�  n�E�o�u�ӌ���&q�������g"�4�tY� <R�oՒ��Dt5���`G���%y�]�j��:U�ͪ�j�b�Y?4{"PD��/�}��M���2zR�%yJ��Rs��W: _�u�
^��H�L��J��W^����S�g�S�UOÂ~Xb���JyZK[43����{���<;Y	�˩`^6jQ,�QX� T>�e�H��*oӪ�z��"N��:H�M�I��H��Y �h�ҩ�����Vܘ���9�Cv�py'.��=ȶ*Xl�XbD�>�`�i��H8R���$:f�IV�CF���GE�p��X��u�}U� �u'PGXFR�:���d�`���I����V~�d��M7v1
P�H���~i���4 �=��\3���~��|okΟ|�c�9��N?����i�ٚ�rb�0�Dߨ����ۮ>�_0���0���xn�Z�e}��t����9�M�L�2q)���ss�$9�5���dp���)�^5Zv��db�{K���K��XH�_ ���ajIO��I5�@�=I^g{�A�1��� 1U=/�����u{i|�RZuN(o�C�
]�#���iL�Y�>V�BP�B���J�PHC��������镇SAg���X�)��k)��7\���(��O]~wz��K
S�e�Y�[;����SJRs�Y�ḶUfT:��L����f3�	��@}u�ჳ^r����������ϸ�\\E5@ Z=j����������@��p��p�J��GfbgD1��P�V�4�Z���,����E�j�|��J�%f��P���X�wѬ�H��ě��V�O#�c�3��#h�.��Qg��l������x+��\����חJ��H�+oX�^q��?�vJ���r�k���T���ʃ�t�g[~M��kX�!�\	�y4a t݉�J���C��[8�?Z���eHN�r����u]`�G9+�gꉇ��Κ�N��iȲ�o3��0��O����Bp�^�������}���ы�V��;#�?l*���B(�Hj���O��Ycu��u����
�X��Z��`��2�wX�-!_JE�W0Xw}��ν[H(oޯ���+!�:�(QM`ͶӥI8���(�1U�Nt����B]��Tx�v��fmU�'{�����������]��Chl���)ܧ�
FW3����Y���o����`�j"�%�nӘ�T sˊ��d���ȶ��C~n`i�u��{'�>{��54��վ�.r(A�1ݪک�d�L �&��>%�a�nӨ�Mq�0B�`�t����As"ρ�
>�B̨5�'��Ng����0(B������}�%�.a#���f5/"�g���#��.(��e��k�p�>M~y�`e$����,T�22¿�K�w��Kv��d�ce��b��X���A�Oc���9.�o��,�xy��W0�7���#��,��`v8�"�<#�{��ڠz�W6T���ziڭ�h����w5���� ����F�{-���}G�R�>v<��q�ՏW��J����#~c��޶�푿�۩k��*�Q&)�χ���?jܞ���ظ�v���6z��#�XG|��S�]�(�z��Cq�����0��F0ab�I���G�����䠡�����{b����B�RB�Wͫ'Ӧ&�͛��Ϛbp��VЙV#�_������vz	��(��)��]
�
(X�a��R�K����dT�9�:�Z��t�����΍��lt|)��Q�봳�}$
Qahd�1ۊ=J�|���"�=�Ezy�	��B�+��<LX�L�ԁ��%c�xvRq�T��ZL�7��W���M>��,�	��NiO��<}�:�W���_-��Pi��8pe���X���ջ�ױ/����%-�/>�+���ƶ�-{�RE�� v���.�"��3["�5�wA�΅3�ִC!�	����ͤ,�pjU�7j�k��8�Ƭ�}�J�~�f[ʙE>DVoi��U��x
4��KH[�R@�!;��ԙ�ydX>P�X���29�;'2��rЄ�6{V��ڝ�ȃk|P;AҺX�P�{����Ei����P�Z�P?�^�Ub_E��6���F]j��F�XE�$��Vo�ֽ���Vd򸄤�3%~GXS)���=Q!�=w�rńo�����A�u�tb��"Z	9����+*Gӭ1늺�E�1�"���L;|ٴC��"N�����|	K�i������Нdk�j첻d��ˎa�P����R섛'���"�Ű��ؓ�e��O,�Y
����7�"�ݘ����ec�
{D��U��}T ��K�$ @+0��fJ�{A�@�]8PZWÍke@��r��-Q	��U\�`m��h�����}�[k��ޞ��ަpK��o� �7�D�����}��:_�+``4��l���L6'��go��;���﹄��W&U���,�85bk��"�*H8%��w%r~1���0�/t��}����3ż4�Ao? P]v�j*�P������.�_ ��F��ˏ[��62���`��O^kY@����,Ţ��!��&�)F<D�%0>PQ-��g�h5��F �܉�.]U?V��'h-�W��H���e�>Io[uys�{qǐ�'�ݍ�RQd�aw��;���������9��c���ӑ�g��5ͲE�Ik]��գ��X<<�1��Q ��}���/�,lm#
ɧ��2w�C�:l�p�!o��Ƀ'
9R|{D�8W�ψT{'��L�7��&w�
��lx���p��˽tv�@Z7v��K~����TM aq-�Y�[�����ꡍ(�H�0�%��S��w/�V�o%�g���yX��<�^KsP������/r���JZOi߲���Y�,�Z�����y#L���W�?(�&���"�\�-������d7�X�&^~��N6�`�ۜ����0���	�зu�l�0^f�Н�~�*̈�<7��J%VY�$5���#�5yC�z%Oʏ~��]���i�� cЎX��ŹI���[�i��(80>B�!ň\��& ��h14�Misbţ=Nѵ��-�k��ձ��N����7A��Ym�ά�
�c��'�B{�d.�2���r�+�5�ͅ�O�tj �!}��v\�����:gPR��P($���P� m'��L�PK���襁]��U�9<��I
<2��1�zmQm�]a�8�K���q0�51h�s�v1�C��~��>zL�WFx��|c���`8F�����lla����������@u� �e�~��x(tlh6K���)���s�<Y
�dҘ�a�:�t�y�����y�]9
��p�S���&%��Nl9\ ���v=��}<�3c�΍ቪx#� )�|�d)�`	;�l�J۾򶔐�d4`d��1fH��z�Ks��L���0�?suPB�Pqb�aD �+~�_'��}�`F����z�'B��G��+��3b��x��?���Qo��` ǛV��lD���Ry����T�?��� "�L�����{��'�W��.}3o �t�}�o�H�M�oఱ��K�Bt\ji�i���ޒAad��T��?�G���x}c5��WB����fk�C�H�5�/���x�'�=�i�t���*eRε.,i��M�[���T5�UU��$�/4�9��� �3���ߛ�n�)�vA=�x����J����O�<�����;I8(��-��Α���oʮ�硖(�u8�4��Z���i�Fi�o�q-�����f�̻�B���h����F+��$��]/*�k$d�b_ŉ���B�[5��gT���)xz�"zj��^N��t�C�M5I�y����昉�a�q����z�s`/��	���@�ޓ.c\��p���%�`h�u;��wféw����n��2l�7�=�] ��74�]C}[2�.l��������c����wz__>i���v�50j�jHϖ�й��-f��!l}���1��B�c��-�5]����;��:5{}<��8!�O/�p��
P�L�2���^h�-_�?����E�}|"�����c@^��S�{!�=4�n3`��MD��Vo�Á�h���O�>�%���y�e@�D���L:�5e�:@��7иEWT}1������W ӆ)8���iL�ԙp�VnAB,�-��xM���a[HC#,m2	��*Vz]�5�Akj���*��� _t�j-uo�R��/�N�YT5��X��Jb�]"萅�_M9�ƭY��%cs�}���s�,zD}-v ±v�a��qRZ� ��'��(_]��zO���nP�O�h�pЌ�������B�Q�%�s
���ϻk�NgWd|$��R��}��O��>fRB�fМ@��4U,Bv�3 OJU���6n�#�'x:�B�;A�|���Oyt���y? ~a�=�I<������%甃޿%�i���܇W�����z@*c�+�c�(hAs���W�g:��iE!/�¯Mѹ����E`ei~>-l=�zL�zI��������C���`)Z���e�c�����62�= ���)L�(�/��*��P�Xe׎i�;b����S6o�Y�J]v���䓐����t����Q���ٚ���P��m뗤1�$�E�S8���$SN%oc�w��e�[�sOQ�yx�&7'W����E��ߣn�=f���*�����"b���-��9`�J�p�e��wf�ʫ��N�����t� Pj�e�t)ק.!��IL�<�'Ψ�^Q��e� ����U`�`^��l����~SWdض���]�t��ɰ����o����lEν�N������iHK�^4���H�Y����ڪ��(O"�vU�̿\����٤NG��^h(�%�9y�A?ๅ���Aݺ�<+����Pl����T�쨠Ty�Ѝ���%K_>G�UoVP'�.��X�r�q~i�I��:(�<�f�ia�eq��Ӊ:Oۍx۫0��@���6�'hVmq�:�����K�31���*�S��`�x�Q��&|] �(bB3�G���7pft]����z�])[�����΋g#z���<��~<4�}(}���M/@������S#���|4K����f�LW���o@�"�d�g�HG<��!clM���lx�l��%����VNi�&.��,yk2������7��f �����?h������B.Xeb�o�8@%E�_��Ԇ�ϗH����t��;���>h��D�p�V������
���n�e�����~�C]~�#�T�@��R��#��mL�DT���x��aa 3 �Ŏ�"/��_@I@��f��w2�ϖhT�UDK���P���kH����������ҊD$��|��h�V�ڄD�:? ��d�D��{3���>�w8uV���xs�T�7��ta���uԐ�W�E�~�^�_��!�i)�VD����'81l�k46<�R�N�Ct.MN��%]���4Ҩ̍��cV݄��A�1ϔ�DtyNj��_,�uII���!9��i\k]�;�e�N^��~�K��K��@^���)~��Fq�g����\���n�7yy�u�՗0�䖼�Q�H�ئ�Nȅ��"���h%v�읹>�體�Fj,�G�1��]���)F}��Ď<��*��07&����V�E�q H�������bP�N�i(ŕ��=�Rj��F�5注+U��' �b�����mD4��v�/��cK+ל��g�|�X���Hl΍�
K&�+��(Y��k�B�0�����CÚ<� �u�%.��
�_:�z�D��,�Y�g�H�ڢ#� �MRU;�Ї3>����S4u�AH�5�ӈ@�K�}ؕ�g/��P��^o�Ӆ`DwX����`�^,��3�Mj,`P�Ǟ��'*I{+�j�=��]�<���V��Ou~��K�� R�{�g�֧�1X�T]ŷ,$P�� J����><S���X�5��t-A3Q��D�+Y`f���>[ #���W5��5�KFoZF�_^~{�.񹵜A~�s���f?[�焇��o��5��ٞ���H3n���mf�ٴ�f�B�i�:o4���D�!��Q�39�!���~D���(�
c��Bb&�z�oS�<@�7���u�o�:�=��Si9��ĩ���R��r�@�J2N��]��Iǃ@<��Cl��<�熓��b���gW;�9������5o�T�k��m�¤,:ڕN�0���yFQaإ-�0�Q͛���ؼ�������ˬ/�F����G�(�9��Ѡ?UH��6�,��.��V�{���-��$y����,!��ܛOn+��@����sy�;Q	>�ي ٕ�״�RJ��}ç~�r�Y�{�VT�`v�ǖ�k2���|	v�3?�3���kkh,O����Hp��o����tФ��gjW��)0c�\��]�a�-�b��e/���;��ϊ�Zs�37��f������wL�&`�m��g)��I@�6ք�VZ�]�+�LE�_
X|X�Sg��H�!�w���+b���#Ȃ(���[�I�0���f_����w[i�+�ˊ��B�p0��B���∊S���V$!��C�����<e���QQ,�8�Z�xr�!N��QrPw�&���I���6 �W���Ś�lY���&�Cp����Q��|��B�uU O��F�O�	�*NC�侒u��^#b�8%�:ӏ�����.�?'�\t�p$g�d�˕K�k����g��*���o��޿�8u҉��{E|,���_Wѝ��Hδ��4��.�s�Ňe�A(�����g#�,��c�z�h�3b��@�}� ���Y����kCU �Ru�(�W�?�if��O<�`GE�4T�Yش�R�R�[�@�yo�/O�i�	0�_z*0��Z�A���� ��=�f4.ל�c?іz���s�1������A3�c���M�M��rf�G��]TN#����D��6��	A�s빴��	6X��lYfnX �@.û�L�I��Ԃ�З,���P���6���_np$�CI4��e��&�xW9��ͺ ��|�ٴsL�JU!�HK�X�İ8�����N�yNw�8m�[�j$�\�!��܂חu��$i�M�>eR]�\5Ђ6c^�dj.�bAiH�+;Q" u>x����n�I�+�qN�E�9���Ky�#�y��ŜS��a�W�+�-h���)`8Q�YH�x9/KW%�s�z~�;L`	�=u�q�������M�nZ��:�U{GJ˥��^���5�v&_4��
l���`wQ-i�����8�&-��#a�|���o+ϼ9���@�|U��W�9��J������Rs�΋�$��������'Ɍ/�
nUc�>4�kL6��XQ1*j���F�hx&s�� �Zr��s�hZur?J+x<�=zl�o�WZ����"��	|�+�눔��4~�2v��[*N'k��g�	,���� �g��'x�=0�*� ˵}Pr�9�s�&�d�����i�<^��ic)��L/a��r��?gI�{�@%�|V�W���~���@�E��*�P�/:��)&���pm�荴J��<�:=#�S�2�v@�d��eao�m�H>���	�S<C`����������>�k>{XS��;��!s�r�4r�k�O%�/��%��b
)?�{
a!;�K�̮uz�q�3�rmE�+����g����[�H�m�CeZ`IO����r���N�[S(x<I[�ۡ)�D�XOЧyt2���L���w��S쎼%`����5�_�o!�U@���y8��uT�4 �����@��S1��٦g���7⨖�j+�196�| �