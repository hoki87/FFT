��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#���������l��U�~�׏O����j9�PY���`T���x���s����uí������P��"��b%>�1eτy�<�gܰ�N�Y�	� {��I�ɍL�ݫ�G�R�k��Q�!E	�5E��.��:�͂2��y�m�-�.E��i�����YS�
��@�H�ۼ��nD��Y�l"BU�.TԊ�=�-�����q���Ǹ��j��ԋ����tr�a�ٵ�]�b	��%�ɔe�)rYOjX5;V��R�������M\�	D��ҏ����9c=�Vͼu��Ro�P�Jf�tRvsY��c�"n�XO��	3g���Q���^�Bʹ�7gQ+Г���$�-��t�8�����A���<����l-��*�|d�!�&�J1lWD�9Y�$E'��wܚ^C��j�U����G$M�����ؾ��O� d{��Tyw�7.�PV_�-Ѻ��Qꭸ�@��5�������Qd� �ӈ�����T����R�\O��-�/��C�I��w#���R]�،�#���p)uX��p5���䩠��RKH����b����C7�̗̚��s�	��)�rj�0�e�9�� �(����N\bۋ�OF�y%�F����M�Ɛg_ÂU�����c�\J��u=�<R@��63{���8q���S��R����	�-�|L�Z��T_>����ZSK��Z혻�~Tة$ �_�p��C�pT�oՑ���[<�5[�I�N��15���8�l	����@�B�T���J_���Jv��Us��If
��S	oc.�!E?\�Z�������䯖�\��_�}��u#Q�8�����P��n|lv19z��W{]�w�E�'#�MG}���Bn������O~��'2�����8�`ƪ| ���M���F���@�n�4��H*��P���MAF�W��3z�?�����*��!|�m?��7�7���aF��L�Ý�h_�[q&w܀��d��Jlck�i��
�&�Eѩ�_S��1e��+j�OJ��b7�l̨����o����M�2��h�ھ�h�	�>������n��v�iX�6�"���|�n]\zJ��rm3:dQb�uT�lB��Fx�ow�r}l2ݔ��K�l�CU�@��������O��׋����/H��1�BJ�w��4Vf�ƾާ�΂|+6�L A����1(�5x2�{��,��z(xv8t"y�[J�9n"��ﲾ�W
Th��5�@U��Z��H=Ҋ� ��˭*��{�x�������/1�MS��3��h��)(�yvf��	!c�Z�f��;��/�[�P$Zs��h��N6x�|�6PR^���V.��6�	�1l��:~�=`�� �3��k�=m��H�a��5�:��</Y<D�~Y�"���zFuQC�*�,}�/�㵢K�@��2�?8���U%�m���ܞ��{ ҫun���I^�|&J����lծu�d����<� v]��p$Iv"��b`/)5���G���Zi�7�.��%'I�6��fk&SK�o�ޘ��Xܺ%[~w3����ґ��� �oMs��|RU{�[O&�0�i/[ӠI�L�>����z�T?_�~Q��Uz����R���r�#��A�4<x��.�1��U�лP���|aS�����pwp(�kv�D��|N��`u�Z.�p�~���q�Cp������j]��T#oM|���>r���/K�o@� ��>�x���:����9q)�����g\�:�R e�+��� gv�F��>+MRJ2��E�ӭ�|�g�lbw�L��ʐ����JA#)�Hni��P%�V��*8)�[^�������E�&͖)N^�{�|_/<�¸�L1P�(�g%�8V���P2�F�9���\�%.ELڜ�A\�
�ӌ4��&��I�O�`��#�q�E\�hc��8Ս��
�9E��EZ�R��N���0`����?O3���3����A,�ϒޮ��s�p4�	LR3+�S_��?F���T��G�
��g4miwN��g�ܓ)��}
�Ə�M}]b�c���J�!z��q:����J�e�t��g�~q�����}�:��<��Uv�HH�t��J�8�V��?/�q$h��G��͑��}g�E�E��bf�}T=m����R5h�qVd����`�0�@Hݘ��s�yn��]#�k�4p�Ƃ�0�eH�����%:-zl{
t鈤���z7���A��cH��y�߁g%F!�d.�hEQ�9�x�(�c���!*�%R�Ѵ3S�+E6O�N� �������j{�DQ��(�$hc�%��\�"��s�R@Cv�1������JR&ΡX������0�&従8)4(XN�]��)���v7�>wG��� ͯ�!�ͷˍM�M��́ʀF�G��u�����q(O�N"C�`�k0��T{?[$��M@��\ �N켪0��l���if�W"E-�/v䌣���S���dAl��f�c�-]Հ���"4��Z��)K!�%�}4x�̹F��Z`Qء}xa��d���LVH0��cTJ]�
t6h�׻!����g�\�GO%!�d�YA���uT�`C�	��.D^"��+qi~�;t�'�o���<��i�������a��/��vEH�����a���fm5qH�� u�����
�C�&Y��k�w} �*���d�#.��¹��R�jVp�4�S��]��)Bq<.��ld�%͒�����Iu���,�m6�8Ğ��Z�c�+$��R�,F��ܱ��B���n�O�-��̩D���~��X:g�7\�.�}81�fbwx�#�#����L;S�EH
o�4��'�.,)>����'��a�����:��%۸�}���(Q��VDL4ubQE��]Z:B��q���^�M�_Ͳu�#w�L��dn�T%T�Kõ�J�I-�|b���_�����W�"��~��}�z�f�{U�]=����N���l𾩔�,O�g`G���)�4�b޴���(�.v���	B�����)�A.}	�{�u����Um��>+`H�H�,&'�9
�by�n���(U��A3�+}6!C'��U�Ee�K��F���ԫ�.|�Q0S�J��N9V���3	dؗ��⠰3G��F��,C*���U0�۝���~�P�=+P��u� ���PHI��<{<A�$���X��T�`��;Q�b,o�͝s���8~?tU�Q-��P�Y��nfv\�1�b.t4����%-&�Kks"&^XF���`�I�]��H:��Y:�T�[�P=մ\�Ӄ<�3��V��!	����P�<�d�M� -��z.������Xfڮ��`&�b��c!���#��(��؅�-�s*tǴ�~@�9��$!� kHQ����$�}�N����Wy�?��ÿ�pbט'm��8NW�� ����W~ h˝�/\F�q�|���l�ew����	����)���3��z����+Q��¾3|�� ^ p�G��t˾UZ��HMu檟c6mN�x�� �w���;i����ݞ� s�g�kb�Q0���]e3�x��|�NJ��U�:ژȆ�l'W  �YYB����L�X�ӻ�܁�R~�ݿ�_&k5I|O)6�'xX.�n�=�8���;_.�<��j��^�]a�L4��y����>�YS�v�!��;ߢZT�b��^tb��V�������ҚZ��o���������2�2bU����Ҕ=�c�M�X�EW�
ES������%E+�z�(�z*lA����)��&d����xe'�+�%�}��Zȳ��	�u��l�(,N�)��|[3�Rf�=9�ҾY�ʬ@��a�4�Z�8��Y�l�h�� ?J�p$k�/Z���g�[�6U3�rh��Ӟl�0^z��N����l�F��T�����*�u��/�Y������cx� ����d婧@Q�3 ����{=f7���<qK_P�`������I%�a�b�7GOPR��G�(@�C��B��j�1P�{g�'sDpcR��'2;�fWD��놲J%Ǝ߾N�H�E��6Fه�l
���|4N=��Q�� ��'?9�ū�%���<�!�Q���K�`n�����n��k��`@�F���Gq#�p����~�����*����'>j��e�k�x'��$U�E�MObV�4٠��r�:�LN8���A�5ů���[>�b8�b���`t�I�;6��`	��p�k�x�!�,Y�,��$5�	RN�~b�&S���P|���\N��.�. V�}[�T\��a��t���Aro��tw�e;�!:�����m�cE�f�bEԆ�zG`u�ƈ���a�w�m捩av�����vg'j��9`�g��}�I#s۬ڗG��c(�x��r
LG�i/GEi�]~�I�S<}9R�d�\$2��@��x�v9ov+t2k�>z��IR�
��@>�PIAA��������L믋�/+��М�10��W#�\_�0��DM{bܾ��	c8�ئ*��V�n�Ӽ������>��2�74��c	�����7-���jw}A6���%��Z�n4��f$t��y���vݩ �H�J��L�������x=���_%�MQ�ǭKd�+�Ic��Z.ń+fc *�,�x����A�\Z�TKUl27�Vɻ���{3%ݱ�t�~��*��r�{�n����|�P�6�ɘ�l7��X�0G�Խ�''��I��"j+�D�+\1�9^�lJ?��14�cp�\KW�~T��L�D��9�)"�"#~3a��ʶ`�1u��� z)0�����hjv&�J49�K��Uӣn{��j}�J*^�r��b�8�∁�st4�W/����mE��P7��RL���C�#�΋��Ta �����@zE(��?9Q1)�-{EFd�/Pd�+Jx#T���Ե�L��r�4�݉��l�2��kOOݣ��l}�Hpr�?���-lx��V������6d�����И�|�25�`CGm%���1/�X@|*¼鴼B��(
-�m~������%����bvB��tp�VK���i�L��lo�+�XvN��s�É���t3 Z����z�>ǱT	��
�I�5C�w9�?�2�WA8�<i�7��d�>�́�y�8lW;x�F�G�K�FQ�P��h���8x9����G�y���Bˈ.�����d��Eg3S��+��#�zȍ���(1^<�ﾁ��پ>�����F����#pL�e�V`�!x���#?3�P��fc����eZ�# ��9�ifI����H��P*P���S�~D�(gŤ��-��$r��V��}A�{Z���zi���B_"Y:t�A��;����P`]\�T\�������92�;%'u��Mb?"15�{���PҤ#o�x���9_8h9���������m.,����F��l���5����Ne�R�M{�H�KE�TA�%��gʨ��|��]��֟8X0��W�1���<�3�4�
(8��J�c�fc	�o.�?2���"�QZA� H/�_�2��X��&럤�.�_	�j�h-ID���/�
&����J�IFX{-;�?��=
�ϹL�?1_#�K��ٛœ��!����1�7��op�3.e&�A�J�Y3�(�����)�6�X?���Q�)�f�$Syh �&�+-�EF��:a�JZ/�C��D!��|y� � �*Sp8J���u�#��@�o�&��C��`����f�`��N��Gc>sX�*��K���7*����;ƅ�L<7H�P����r�v��H�q �m�����hSÅ��(D�}��}��O��˖�L�0)
�\�enܙ����[sj���&.���m��pB6��i:]S�-�M�.��!bb�X�j�=�J�;u��/ы5�>0�\�R�E�%����L���z����|yqz���n!b\�:�L�(%{�Ƶ��k����up�0$&�YSF��Y��T[�R��_
�Tɻ�c�G����n�vU��@Z,�#�
�
91F ÔQ;bp�ۿ�̓�j�C�����]Τ��9 ˄�P��n��dI�$�]|{�����(��.���P�"�,Sw	���F�Nc �9b#zX�nb�Ha��z�R�`Ϯ}'g��y�&���,Ptj0�v��� ���!�{�'����{���I��0���l��Z����Fo��OŰd��Ǥ����;�dJ�7�c�uS�d�;4��{v�2�.���o���.�W4w���T�m�ŉ3�+;]c?��Z�r�������U>��-�Z���}��x��8hBW�x�_����HY��,Zp����Y�H�K�œ6���掌�Q��N>!F�5ͭ*N�5h
9 �5ep~ ��.ǿ��%�|���s����
o��
�8'w]����z���u�3�\ņFA�I�������Ց�i�����G�\tV�ԫH�nWH��I���C1�)���i��3R���s��񆷓��a�m
ϧc�G��o����<,�K1��?�G�jc�3E�}HB�$\t�:��E���ᢨ�yp��	���R����F�������M"*2�D��|��x�N 6`��e?�  �gڼ\�s{�븸9�r��*�tE���Z�f��j86m�f�(s�`B�ˉE����Z�����ȇ\uq�Fc�^*�l�AW����.�YJ��;�����L��;�Y��׊��>��)�w�A�3�����ƼJ%�,�y��s:�Ķ5��Wƭ	V��T�lQ�F}�$'k�+1)0x�q�@� �Ay"."s�l�F�ߑ+����Q"���j�qC��{�j�#�MX�?�	��]˝r'�*"�W�����@�-��N��{16���� ��%�((�����-�5�ʏR6�92ӽb��B�F���̩v�m�xR���6~df)J3c���52_;���݌-h_����+�fE ��6����K]{��.���gᰍ�>��0N��Gҕ�K�2� ����6�h�$fԷ�Iϧ� ��*����s\~P�2�Z��Hjģ�q�w����A�4��E{�̤��Q�d�9�'/��)k�����W���h�L�w,A)�3���FЊdSn�"�/��\:�p%Xz��� ?�'��w�e%���=k��Md����d�l�m�kT��G��{
��/1U�Y�F��5h���v�����86D��rܩ4rN���.�u�X��JN8ci�ģ{�u���v1���Z�z����,Aۿ-�{}R�14��OJ���D{����6E"1Щ#vN�k��MA���5k(9e�ir�=Oc�:>mem���ɈPTڔ��C:����
����4�{�rF���l擎B��}������y�յ��P�a"����iǁ�/������8p��D�h"�)�J5n�T:�f�
�D�uN�#0gL��X����Zj@)������T�q��JyNf���n�s|�D��-
%Y�	]�|?��F�C��T�*���������1�`f�w�"O8��	H*L�o��o�<E��y�Qs��)�=�
�r
�9�^I�^�:{ �����+v��w�%�3�\?�p ~b�Z���ּLr+�x���'��hB����YH�)s�s~�d�r���)����8M;�e��-9��r6� ����;�`cё�?3���3�7�ÀBff��зe�ɀ��s�K�QZ8=/��p�$�ZV]@t�j�zz����F�N��'��X��V�#�*3m����{>K�R��l�nb��M��P��qr&��ުSd��~��G��0�#�� ���߂�M45YT֛&��{�/���N��G��z��Ce���ؚ�@o|�dot�t����ڨ2��=�eڷ�.�X�Z�q�k!����ڊ|[�����B�1۬��Q1�Q��Z(ٜ�wL~昘F���j+;deAl�N���I�������c�W�b��\�ʦ�4�~�nUXƘ���%z��M�?p�7G{��� �	&��zv�N"��ڭ��IBm��ؿt�9���9��x��]EXj�i�Wb�"�5Q�B�2�{��y�7�hr�����Q�Ңf�����l����2&�IB�'t���\=\�v���`y����X5U{��C��iϖ��GGc��L'N��2r��8X:�J�Px��o+���c����Ң,V]-���o�ٕ.xid�^�MW�]�����<*]�C���~U���sէf�7����+��p���#���R��+.�l��*`�u1���]8�w�TQ��v�'b�E⥗J*�y���JEa��1L�;�P���h���{��`��G^�=_
q��^ۘDS�����&��Gf6�kV9�����vѣտL���m�3�Z	�rX��̛z�}�'����t=�/�lDS_�L~4��.%}U�_B43�(�#��*�^W���{��ż��#�Ӈ#@(?�X��ݿ�I|YJG� M�Vf�Q�Ł=ɔb��G��G�7�K���Z�oo���5hP����ś��~-o����\��N, �W�I����?�C5~E��t�����n1){x��L����4�
��e:J����l�ڎ��n�#�j�3�&�� 
��7�@�.��'�_��7�x#����>m+�ҋXݎ/&���Q.#|�ͥߏ�Ҡ�H�9�:��F�_>��S�C��:r�P���Ǡ�Փ@�--ΐ��/�%��a|oIs�9��W���y�r�����ֽ�3� ��$;�$���*iO����t���,�K�)[����q23_�[����X/��� ��5����E��B�GuВy��\��Cn��Qr�����!Z�z	iC���h�s��>13�G�}�V�9ݸ�n�e�l�w�Ȕ�ذ{�$)��f��*