��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ����������h�j���%##m����Xa �� ��T��Q)Kh�,s��s�� X����π�@.��E[JLv����ݕL�2��ALq!��.�ڱ��Cx����ߧ�k�)�>9�x&�a���Z;�m����8��2�� �+ *A����E�FtU�PH6Q6��"h����.c�M7�o�
>��;���FRS���J�n�\��>qj�%���L�R�>���	Ǹ���H+��n�`β3F$R���|.��p��˱�r�U�� ������J�b�����*\��Qw�=�G�N��ς��J�7�>��p��ru4��^W��RǙ�a(����1�Oc�8$#���K���d�{��N�B�<���;��`�
��Y��Ⴔӈ�6҂�l;'�C��	V>��s)b��2.���O�A4.&��d&,��\0r�?Ѭ�>�"�<�z����T�*o�[�
nf^�J�w�0ª��ߜ�5����Y����U]_\�=��������� �s�=�8���Ǿ�C<����ߘ$�	a���)���	��t�X�e�M1����S}1ܩ�����C]:�OЬ��wm�~0:���F,!f��n��跡��$��?I5
����ݢ�
�X��]mǚp�ԽEW��~�Ʀ\�0�r�&Bk������z���JáS���%Vo���2����ZJ=����8��N�50|#fr�`�k�:�]�,ǯT.��5�A?综���l0W&�Js��_���
^�{6�[��098am���bI9׻Ԉ���z��ޛ�[�48�ƗZw*��5\�n@��w�mz'��:��`7(��/y���"��5c�t˙i���R�?�.�CǸ�:!�&g�E%��vK�S��\{}{���؛��9�t�OȾ-	��nN�l1���ue��)k��藀rl4#N�d��=D�>I4wS�����c�'D�C?���Zo�An߮�~y��=���W��ti��]d��P�}�����^Ucc����,���['Q:�};����r�~�O`'���"�Q��F�l�F���i߅��~���W�1{�����4���#��ZF��j���qXcd���H������/u�^Oz����#Z.?�o]a)�H˹R��F���a��Ulجq�->�S�'��榀xAx�# �\��Ά!��p�����:�2Ѝ!��E>W_$d3�a����	�������<d�d��x��RB�P�%�nk/�}�Kܭ��{�q�"��K7n�SQJz�dD�3�<�#��"�P��g	�����P��ӟi�������)�>���_�/���@�����p?�,oݳx!�6� rcy_����t�>�ZS�WOO���nu:`K�*W徻��S�m
Z����^u��GC3.9��	��<߱��f�WGe0�i��f����L��K�:�BE�]��;	��\�V�O{����6���=!�Y'�k���i�_�{��	ֿ�ӖI���B �HyD�@T<?��(ژTG����9 ��¨����"��r���V@r�g�uP1���{>x�K:�Wo�ʜ��\�2�$o)�S�ο@?7��ٹ�f;N:*���?��on��f�J���t�/�u��:V�.�M�)�҃�yq�l�jX>�=�mÅ�;}�ʉt���c#���7�AUȰ�o�%w*�P9�s#�q�IN�Fvi��������w�N*���;KI�rKB� ��$e��3~h���9R�\v�E-ID��?A��i�Q� c%#g����l/O��SqrǤ��%[�z�Z��*M'}�O�E���@�6@��� �b��>a�4#Z.� ���4�J~)�.�V���pRQ���5���e�옑s:��s�}ϧG�z��&ѦAV(���]}c�1����n`�ԓ��*�������+�e������j���C=Wٓ=N5W^#�m܅l�����(��W� �	��zX�Bap����^z�3�Mb�q)̨�ߎ��N��o
Y��i��sx�~�_��U�[�=�Xw]y�؃\�#�W�A#wb](^����� �I�ͣ�������M�`����. �%��e ��o|Nzeӎ5itl��SP.�h3��#w'�5ո����L�0Ɯ�'�Ue���Ξ�����`�I�C�R3�Z7��+G�h_)ڞ'���=�ͅYN��ҥ�߬��?���hm��,�u��{�����!=ș��B���2��"g��$����k{���)�k��΀����|����*�g?����+�[ۇʭ��*g�����~{�C�Jz&q��3�`�g��E�&5��h_ִ�j����LvX�O[9a拢0��}b��d���{; \bl��ȼ�s�r]�Ϟ�e}��e�^X�)�r�Y�_�F_�cF�T��Sp����	{�r�N:�]=�����}EB���<q;�~phЪΫ�c4��q�@G=q����M����;� 7#�����'����� �$�c�R�N't�C��B�"!�5�X�΂�l`��u)��(@vGh6Q{���a.���q-�ƅƁl�W�E�G`��%?�}�����/�4޸�ɰ��;Ҟ���w+�=P�[#6/<om��#�4^��,�@<��!Q{�X��+8�<Yz���vy�m�ƋYIsn�袛ϧ�@�n��p���;�QM�$g�#�JX��"�J�� 9�;r Č��\}bxC���O[F/J��"d	�m��L�
}tL��#�j|`��Q3+���YE����?"Y7������ѵ�
2c�Ȼ�7}�ʜ� ��fRK����Ey���^/��uHe�F����t#�[چj��r�%A��p��([$2�����<]�� N&32W��8oR�$�s{[��ƉwjڦuW���ɩ3�`�v@{}����0BM���1�KhU�e��z��Z���	����q������腶y
~jÍF<2VΖ���B� ���&%��&i �К�͜�>�ДG�Fv��`��f�o0�;���s?b6
��I�;�v��[q���˪�bG��~�Q`�����N5�&z�#t�H����Յ+��[�/�[�ayͿ�a&���K��7�P�0 �u/��|��N/���9AZ��J�� Vv4�)yM���i��7�8Z��]W�	��+�*r�Ǐ�SH	���K�ʽk���Weԃ�/o?��ۀJKy&׬2M�%��y1;O��Qc�$���T.��{�tp�qc�Z�̿L7&�g������J�U~L0+ϊ-��%�;��Q�1o��	��3��������)ypBl�Zn���v��v�җi�Bh������f�uk�^��n�p������y5�����&~Y��W����t�P�)!k��MǶ&wG� �V�~�2g���c:��7Ly�\�D�*5����EK�p(e��VEe�(3����0�O��^�~hӍY�Z(�PN%E�Ē��������f��1��TDBś��]�#��Q��\���|�hJ¡���iv�ۧ֯7�jvz�,��C�H�6�Df�%h���a�#�?Ѝ`��X4��IG0�1��ї�j�9r�5�xJ�q���\P�{d�'��\֙:�{��j{?�8�K_��٧�:3\G�@��uDZ�0-�m�����&G��̭����x�cB2D5����}�{���b��DVI A�{Rj�[�*K�m�J��&ҿ/t�9���ȋu
c�Y ��3F�B}��4ETQQ%�[��\������Ft�����s�+e��.5y+NH.)�J�a�)�zS��I��on)I+�&L����Fƒ���9�2��v��j�����q�%&}�ԣ�
��\�&�n�(	aZڟ@:�Ƥa��`�z}eno���~~�xY�+�3x\�@��d�f�}�Wِɇ+�<�#l�T>o��Ȑ�� �bҹ�R�!��ϳ�����!�p�k<�6�+Qk�~�%HIHN�3V
d\�s���!n��7R1k�B��Fאr��_���^� �tӾ �� O��.0�w�ֽ��m���~B'��v��BT�j��4:N��-0]#fr��>�E7�*/�Ƙ���d���t�`��!�l�Q��u���['^���cݻ�3%�dD&0o���C��y�
��a^s�݂$���Ö;F����d*�[-�F�=l5���d�(S߬@�T�}̃LҘ���%�k���пG������}�9�n�^b�Ea�=��7�a��vn����
�s�� �-���	�G/�rD�b�E|���i�(4�F
ģ���*LU�#e{O��i�놋�yY��"�z�i^(*g���~UR�,�������%`?��zAJ:���N�V�;"K(J48�ҕg��03�N=��mC�wf,��v5"�~t�y�DLn�!U�����SA \TJ�p�;�5������z�:+�~o�B����!\FYy��ܐ��D�����%Z�8�nɢ:(5e]�6E=��V�r�����������}|�<QI�Km��zz�>��?��l����z��+��ed`�>���S�W�|�d�� A�ݹ�`M�����ч���
��nN^�u8�|�w#�~�Kx��E��J�p����' %laА| qSI����GĂ���S�\��A�0�@��#E8>C�G�)H��ܮ]\�i4�y��|\������l�a����{���L���Ub�u����\+6��y`��02�\�fp�̐���O�
>���,�p�S���ަs��1	5df�&z��w/(=�i����=f��GrS�����X��4��h�+���>������:��9_@�E7��¿�Xe۴��}��c�ҙl�	�q@������J��o����t��^��y�J_e���� �T}�����,{Z�O���fU��(0h$��s��W;���tdH�޺ך��h$В��-�gS�AbLq����2G�UDW��7�*���P�N����b"/:Jܵ���:�Tf���)ϵb�D�Y݁;��O/�婃�:(��S4T�@�c"�[s E����E���|\�I�t����+AټO���ܮ����ЅXSQT��A�'���4t:����Bp��IDR���;����U��=�M�&W�_/���5{�ޞ���Cz��<�k	���|6�Z$&O	r��o���G��8����R������]��D�J�i�&m^���
�/By�l���N�B���V�Z`!Mn��iY ��F�ܩ�:��h<t�$�����"V��Z>*�N�2��tz����6��>��5��]kI�th\#�}YA������V&N�fc�h�)�#��^���ձ����"��b�� �L͌�
{���S\)�zٿ&v͏��1v2�T�G������i*��XD)���W���=�gd!���z(��XS-�������5�AA�����.�}��5�z��U�P��֒�+a�u9ȡP4���P��=�2om��q�:AZ	���.��2�`L����x	 ZJ��K��������cC��D�aS4,�����P�G�+�)�8���|.��_x��7Mg�(9�b� ̅)v@�\�����f�d��q1��s/��2Q����U��ܧ�G��bs��oA���L��̩j�u�H�������G�a�9���W�x�!n��A��i^?ɀ���FB�Y��rk|M�<��t��&��ik/��iB�F7�j�@����
&Ѫ�L)n��^ vJ��m�З�X��B�	�l��"���bL4��M���i��D�*B��KS6���Kʽe�t�]\����m�N�4q�h(<Tw"es ��-<���&�������NmL4f߼��EP%X�j�ᘟ�������F���mt	���omB0��Rnu�;���a�Y�R���$�����	3*߆�`ɝ8Y+��wv����U����<�*rJ��m펌�%������� ���X���	e��D���R�y���+��z��p{Fa/��p�C(�g:>cD�Q�!��_bS�����{�T2Y��]އ��m?�(g���8�L�ޏ@��2ݽE�Y���`��w�m��,F��`�N2�T��eh1'� Wd�5���t�T#oR�0:��ޥ�}�f�@�-�#�8��}0�w��f���V�b��$���-�_��t��Y�� ޱ��������8M/�+�/C�_˵"&t�}���<CD7��k,��)P4֓X��K֣ hTT��f�GJ*���Í5(���|��m��`���ǚ��\߈���йN��Zd��{�k�����Uv.�L�X��1�1qj�
8)Q~Ŝ��`i�6��j��!�@�Pr�>�)?X�ԜG�lbr�%M��T&�|?�t��V���9S�?)���{W�݁U�bnqj�����BI�sK1�4�b⒈/��7���q�[�|WB_��9�=o��_�C/ސ��"j��H��V>o+��\/i`��r!Sv��	`aPm,�
&�����\�i���#$!����8�����TC߬�3����|����$��fR�ҏ@��xI���%̽�Nj+W�+�uq�kZ��	�p݅���!]�A�IR
'����{�p��l+O$ќ���������U�����+w�p�ivR��N����7�����$o��5e r�ͼ$.�-��6�����*(`Z �k KQ�'�x��`c�<�N�L���;�2�p��e��8Yg
.դ���<��MA��ł=�t4��3���=�%�Su�<q�C��@�%D�D�V���~r:A|�����!��t1�,� ǖ)N	 ^�*�h�ӿ��^��\�Z�_�_n.�#Z��C&���X��](&x���L� 3
�9_���M�>�n�#IdO�~*C�{�lk�����	���(@i61q��P�1r4^��_~����oF\�b���n�Vu�P�;v��s���
�/́`�����jy��v��a'm{���SΎq?��P�����0%����,�I#������S�� �q&h(�R��A�*+�k�MYL}^�5}�����D�In�M$�
�\��~��v�7Ex3ݻ��-F�!�f�!�� ��]e�(�(����{GN���D����Ʒ�-��aPJO�
���I(�9��O
����45�Du��@�_Fa���N��k$�`�J`:"��Zܞ����"�"�4e.��$E�#��a1���E�������<�d�$��pr&t#C� ٌ�����Fr|����IQ������P�Vr�fQ�y���_=�?P?u�X�D*�� g5aM߫�����@���c��ҕ�2< ��Zi2��5sx�JE�m��_9��/�QWR)����h��L�����y�4JŅPp-�xI<%E��"�E$�@)͡���� �x�h�w#��G�L~e��~؍Z���J�>�0��
��)8��"��W��gȐ�fؘi\Uh�:c.�I��2��G��Q�Ґ-�i.[���}��6ӎAu��o � ��=
�>�_p��`*���o�t6�ǰ�Hf�҆��X��0�*�!�<$�ZX{0���;�f8�6��q�S��� �N5i����g��'vH8n��-�1� ��F�L�Z�;�|���
���1v +w�L	y��C�Wo����f%��2��jD3�1oS`��C��Uɜ���JS��gf�_�.��� ,�'���Eb�{�	:ť��q��9YXg�����~����2w���
l���A����������sbW0
�P$8��:3.�1ol�dͶ��'&a�^��I@J��/��j�C?�>G;Z��1�X�� w�l`,0�$���!�ǬB��͑,bJ�9��=^]��nZ��H��Ǡ��\�f� �����O[��ݝ��^o�X�d��z��9W�c�Ao^����2>�g�<�j�P2;�ٖ/����-Rl�>���R��-%� �^�/Kx�"Ǩ��݉]�2'��O���(a���%v��4�So<SƲ��"-�j(�9M�X��+�Vڞ��]M��"f)���P�ji�,��N�44�Y�e