��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�#&��#�<�����d���o	�i�Y��ǢNFKR�r�d�Pє@I��a�ڒQ�6�: �m��H/S�ߥ��x5F�
��,�
v� ���U�͗A�^��!����f�f�Lx����6�|�G��ӗ���.y�o�Ke�_6�Nl��_�]B�����8h��,�GK��:)����-5�%�D��#�8�b5���=��@��Q�iH:7d�߅P�W�U6���<�%��6�8�2�D�uһl^���壤E�_$r�������ƋaKo� �)��6y��  *4��:���G����t�w�n�96J��A�.�&��:hRD�$��aS�GAkk���C�G��6	�R�5$z1]�)E�]���hCP�ll&��\�l.O���� ��w�~�6��D]����ֳ������Z��6�Jr���^�{#|��8E!�F���/H	�äU�$#�����<�r�:��J�ȣ�4�:E��B|^�RUbHM�_k�l�5���ߓ ����A�P����������Z���>�eUn���HmZ����e�p��f��kuu_��f�V_��"�r�2��K��f������񭇮�i'�+�Չ�	��;�5�|*X#�j�1Q��O�{��b���3�Г��e]�����b�I��o�s�ק�w�FYZ��<�.�������s9�>?���vl���K�$]��t� 炷�ߵyP�o䇓� ��ɇ���ȏ��p���-F<���I�>���
Tj�1��`�\
�l"fv'�6�F>��ց�O,^�z��k�����e[���w�X>�=�Q�#n5�4�a�1� >�����یM��m����!�n�x�5�.�SB']��tm��8L�)'zNυQ���3�m�3f��R���'�V���1��=������Z%��ZǙ,����4�I���/��ىǂo�dA�.]v�����!�C���D&�TF88��:���ɨ��.9��*�^�d��	�#�%�t�!2B~Z�ʾy+���L�����;����RǠ�\Ժ⫻޽M�g�K�̩9��X^���l���8JRHM�1R�)�<,X��Bk�١Ӳy�.F.t���������\끢֙p켟�F��3��X��vyI�>[��ڭ�`~�0���Q�+�2�%<��{�i겭p�����2�I�^������F��!��M�	�5H:	^�h�3�>�[��_"�~S�ׄP���)������I[$��ZYm\�Ί����(de�:�k���k��^�!>��/�̰�7Fu {�m�O������(z۾ _�놰�%�gW��?��6)G�َ����k��.��S��m@CES�U:fC��	I�n/5�&�m=�U|}V�̅»�&
�}��T��#���2iw��_A��ݞnNh��z��۶�:V򿓌���g�	�饈�L��IG�EK��I��vX�F�����}�����/���`|?�\����Bk��ѿ�Y�I�~wm��c4��9+��WZ����L0p���0;�#K�+��-������&T~1��!��?;�դ���B����ϗ �sƛDegE�o�hA�.��Bcw��x"b��<y��'B�����;�tZ�3�`�L�|�4m�E���N�����aMۤ��ʒ����XR*�n��~f��ޫ=x7���t��}�t���f%�FS1�e��&wjHyD Ǡ���G������G�.JJ��|l�Ȫ+���xݩp돰�{���u���ʠ?�<T����� ������X�Ѽ	�Q�r����� ��<�b�jLKs/e�ڼ���L�d�Q�h�� �k��:��GԳ]Ȕu:K�o�-p��=o�0\h��Ogd��"��J�ꞁ��ȍ�y�L+�Q�	���i�����ϸfD�k|r{�	��Ex1qd���gwNj��C��]���8��T�IZ��	���C6�oȃ<̀ϟ�[�.Y�t4�%[P2f��c�7�3c׷���4�2��¡�Q}W�H��<�+��=�׈��hW
�T�r�����5���m�6�\�D,�H&�y�}^�VϷԬ��f�O���h:���q�^X^���pP���#�ń�uw�`��1��4P�[���B.b�u���
�k<-gq���X�ci�wV�������-�%O��!9d����Yo��T/7���W�0V��*0�ۂi�9U� ��!YZAI�ї�J�ֻ�rȲ]#�	�Z�s`]���{r��J7���h�=��4�J������}�٣���H�K���
3%�V���������r�t��j"��k�5:���;-����d��U����f�%�GZ�<8B#ң����ᡮv���y�my�TLu�{UR趣I�	���m�y��U�)���_6p2��8���:�n�S�@����Qǣ���f�:���=�?����bS�P0I$��5�p4͆���Gv��%���.��,�W�K������1b���q��!bj�{i������>��1��_}﯄#���@�Љ\� ]{�����Z��/�#���:�<V�gXq�1~�5���G��6D��,B������L�X�%dd�������{_?�7�01�a=����<�����f�DJ���� �߀-��Ff�:D�1��+�~�������"����mF[��C�'�GJR!3�}Q�8W<p�*I��<�|��	�͝�� ���\#�~�:�'��rJvϴ$j6V���Dث��ޙ�T�U7X��^EF�X�^W}½kf��2ԩ<z$*X;�c�"+��A���-(̨��Ȃ>C��>g�d@6"�W[�!�lτT��g�C�����ݾtD��3�9֙%7>K�i`+�C���!/�����OB!�/2�CB��k�ĸz.F��s��{���F0�4��W3��o]�&PI��;���Y;٨�v���*�����U��k䰅�@��D��&�Gh�x�t��:�aY ��02�c��L���GH�O��`�0�S̨�v��H,�V��׏�g(apsV����2ތ������r�>k"3���L%�͔�(�?�܊4���c�b��h�vId�Q>��|7�ᒽ�� �m�h2�3!w	�v���H��K����c'/R���l�-�2�PM��^��6�CD3��Y��3.�F�yp���R9>���f'�ij��Z�������������%��x��;{�O�����aX��y�ڭ�~�	ͺ���H^뎇�Q�`=��t����7����iX�mq���p
����O�*��� ��ʞF4�q�I�Ʀ4b��v3=ձ$���ӒE��������t��D}xd�?��d�􂆺я�lBy�V��q6�&�
��{��ɛ�����o7	�5������O =l�=c �kڥ/�x��6/��,cÉ	���.8_&C~���$⳽��Cw���+���-_��7i�ߦ���AWZ��ɲ�$o{�g�D[�+󷔬��n��i�U,쎊�^�[�d0��!�v�@(��-��M����4�`'͸*�Z�~yڄxMK����m��{�8�����)�e���$� ��CtP�A��'d�V�O�ݒ�7�s�t2��.��X1�;����aev�Qg5�,�`�����X�����Ӣ�1N��	F�9MM�J�Y��-qO��x����q���.�F��-}G;�)��������V�eo��G8=��$�	�=�q�ig5w24��.^	W`}�m=�b��z{�/y#�(���?]���K��\��;/Q�b^�����/�s��QV�=q��aJc�J3�=D!�v�7-���y�(��A�e<H��QG�\i��c��LY��C7�:DE�z�R)a!R&�,�k�{(9��(UZ�y����K��^�/Z��k�hu�p�N�j�U�Kڊ=m��=[�s�[���+��Fp��+xF�����U|#��&tx�O�N:S�\�8[q��uaO5��0�)��7�H�+=�U���`�;�F&��5ݩ�C�S �;4����f��՝����B�7�qrk0�TM`�/�Nv���w3N6Fz+,��5>[�Z�ɵ!��y�@�W����Ğ�=*`��X�!��!�Y`��!g��+�m��}	���7 ��ʮ���.F=�/�Z:�	�\:h\ �Ы`q��g�Z֛?uA�mj�H��qf�{!�>�17ƌr���6&B-�"�6͏�Mh�D�c�/�)̼������:lD3Q�"�2��u(�/����%��L����zVR�n�=D0K�Rb<Rg (�}���2��[�����#���\R���'��ʭےQL��,T���3���x5ux�C��_���ƹ'��r4e��JjH�oD�&��`��LQ������/��/���Q?��xr�j!��!�}
�C��E_����k\L�0����BЎ�w\HB���/V�t�|�s�k��I~�Qv��[}e�;]�0���lv���:�8L�Qi�×�Z9u_����zz
�n�+���12?�:R6�2~x�����O{� D��J��SOJW�{����>(R�ʆـ "�rf^���GER�xƓ%��:4֘U�qVC�1-�g;�N�ur�a�R��Rv+�J0ΨY�_��*lyY�q��6�{�i#�B�I�2K���Ѫ��4��-q��\����x�~s]� ��\��nF��ʛX��i������ >cK<�(|�`0hD�c�,��襒�>3m�m9,�zL�~=�M�s��a�����*f���=���G{���8��d�j߹�����ݼci?����]�p�7l��jw��H��D
�{�^�u�aTO�1I��Z��	b�z6ts���-B1y�Tۚ��4f����mj~g���X�f'c!2�s��6 �$�y�@���j�Fn��5�.-Ob��������v.vx�O~�&3P����:�o�*:H�-�����ix�k�xL�̜/�k�<3�%t��r�B�p�i�|e�= I[�����N8C�!�������s2��?%^��p��;�U7���` /���<�:)�Q��z���u��l��P \N� �ވY����ʦ1&A
v��]kz�&E�	-�}ރm�+�)�+u:���C�Tu����/r�P�8�3�C<w.]���%�/E:[⇵O1<V!FzeKz�^��&q�Q&����T�z���#iB�P@��Ixݢ��=0+����l����y֨k�,߇�N�sW�<W-�[�&Fw�B��)8A��q�y�=Ŧ�| r>�ܔc-�N��Z�j`7el�@d{��6��i���=�Ǚ�MW����4ӝ�z��sF����g%���,ҧ<7-[n�=g�z7Qr�	�~�S]�&׽ ��An�����j�޹ �w^��*��y$��9�7�X� Vh&]5�9��i	2��6�Gw�+�.h9<�T���a�N�Y�$"GM���m�����;z�	)k����M�3�(T�h]�)v�Y�Ǔ;&��^P{�K�w��3a)s���<��~`�,�U���̿j�%����bÑeQ�{K���H�d���>HOF�3|��7��-�:���W�Œ9�E=���8���.E+DM����Ѧ�}@�y�N0y�;PR���o��=R ?a���=�[ϛ�X�$���M��M��do�JǦG ~ɫ �p� �W�1@k�ь%���}�k�@18h;b��0>M�s� �q�NU�u\�uݶ��z4z�~�G��f��.�i�r�S�Я���&[�P�9�)�j��`;�-�h/�L�D���&<Ur�v')��d�*ܹ%`�`���� ��UIQbF<�2Y�p��w���bYs+iI |��#���,���L����b��jA��8#g' _����z��E��1X��+=$�@��z�^k�@�łu7��L����p����<� �d��0�{ڂ����5�����
�^��y���n���I� ø��Ĺ"�誊�T �̕��8�Kk<F�T�[��e�
l�D�Z)�q��(����.��1k�q:<:�K��ˑ,=�th#s$69�G� ��r��'Y@�ǐz���hG���p���i�{���:��Pm�.�.8gAEYD7_@��9iQ��`�L�A++���	 v�%�Ю��%�.���?`��=��	}S)(�z8��v��7��l f��3<Rۗ�����]H����jI����H�^ccE6�����b�7�dxyfIeqg�U�f[����Z	q��ë8�H�=1���y�f���������l.�F�OBֳ�*1��b�H��y���k��o�m�z`�ߑ�1��Ѧ���8n����b�f�C��+�D�1Z����Y�/D�9�3��bW(�ˣ�Z���٨�C�9���{Ú��(�t!�ۢ�(d&ǚTNI�q�^{�8����:z4$����#����f�S3B�?'�hH@���M�D�l�҅q�n�k9|T�LVhVolp�n?U�Đ�C�{}�f��x�ϙdk
tK	g$�9�'����̷sC�����#j�nF�]�]FUz�i�* ��ӯT/e�y�1^y���D���;Z�g�]�B2x*.��*�����	<��XXS�ë<!�O���<�1��=]@�V�K����}V��v� st�~�m�<6~�ն�&V{R��Js��ײ�n)��iv�5�V����{��,?k���̅yW3����U`\�E�Ȣ�l �����:n�7��.�>S�P>�4vz�1�]p��� ��mI��)0�PVC��yA�(��5QW6�����Ѥ��ZD6����p�?��B�,�m� wܕ!�H�v�p؊��̑xH��/��'����OH�h�HQ��4�p����豈ڛ[ �͘`y���6���k��V-S-;�<1ҹ�:-&�F�P�>>��!}�E_MQ�蟣u%s�n��e(3��Щ�CC�G�`F�+��M����5��Z��7����=��L\cNt����4_4��!�{:�|��иJ6��z��M&M�XwZT���0޸2�٤WA�XFHF��Ra �N��EA��tk޼Wt�jF*�cȊ�|��	!����v�喾�V'{� �;T�7S%4[=�d��^�x�II'ݞ���Q�_���]f~��y��7���ASVt$��Eym-S�qY3C̚F�St��w��>�б����"���_m���F�"�x! kN�cԹ"�[а�bRE8
�i��[4a��¯��[-�!�����ƝA?�k���:�f�(��d��<k��}��]UI>I˻X��%�A�b5J�D����@�F28�MP��y%_pk���,9�d A�S<46إ\̏�>,O�]/��,�S�K`~}ϤD�����썡��AM^s�w<hT#C�ƑR8��B8�
t��,-����]�!��l��X�W�B���he���x���,U
��g9l��)D�^NZi���Κ����,E�)y�J�Gd�х ]!I�G�Z?N�[-1�o��	��*��s]H5��C/p�eDn�+�yϧP ���}�������,�3�e�����$��`6���	wc��w'�|���81��De�_|�|�p��u\[K� ��ݛ;u#h3�|e�uo<ϭ=�?�H�#�N%I�S�e�~oӡ7dHG3��mXm!gA9�{���h*U��\#l��C��ֺ]�-�-�\-$������jB���ё(p�Y��_��3U���tB%��Һ�8�@�`D��0�q�R]Vo��e�бN`���,hpN{J+c�l-�h���4���@�ѫ�n/�� ��+�7\��]�$f	//�ը��e؟��٫Z��<��%�U�:�n��i�F%����eȤ��i��$b�k��˶�(�=!h![�X}]���|Zʟ���J:���
gi����D��f÷߾68�Ҝ�;�I�y:�%�c�)<������#�ط�V.'��
��yD�J��}�1��kN�䥛O����Hw��B�����U�p
���ɩ�a�nD |$��B ���1��;�s��+��/w���c�O55��O^%r��yZi�0T(�M�x�G�~@��#�^k��P�2ђk��q��ĒK(��+�u<�h
�*���8�1�<A���A�eX�oiu�%ӂ"�\"�����v�2`��N�c'�+]����!k��*�:�(�v��K��.i:<F�U=1D���N�W >�b���&;��6Ƥ%S=���<|��,�AE�y�+��v�lS��|lfAnѝ�XGU�+E*�ߝ��pl�6'z�_g�[���w�#h�
)��2vN���
F��&$8I�C1)c�C��%�z���M��j\�by����I�p�_�As�ޫ[|_o&L�Wms�b@�o���O���z�|�X��ճ���B����;���9��?i<�ր���/��&�����h}(�t�n@�З6�%�  �
~1�ϴ������Ɩ�
v�7�]J�.��ͭ	�wddL��T/��h!�U�;���R�'�֑r�ԑ����������=���~֔,�@����7�� k�Okݝ(Л1QiJ�����Ӯl�pXҬ��f�o��D��v��q�D�t�uk;ٷb`{���A��.L�Q~}����k�qE��؝�P֓�����e��Z���Y�NR���>��уʫX�*tR�=������9[-5��x��&�3�H(\�b��,�]�B���d��7�!���_���Үa	��_�r�	�a�S�=��t�ί�q=9��Ŏ#�,�![���qb���Xz�t�Q�?&3�$JY!���)�2?�b��ݤZU9j��+���U4�m��k�˞[��'�(D
��zB��f���s
~eS��̟ɥ����5��T�]d6V)l*$濤��Ļt���8��o�)�?[�Tg�3b��&��N���҃����̌�' r��B���j�;�[���G~�Z�A\�qm������ �gg��p���qq���ʹ�k��w�{|�n��>L�tF� -��BH�G��N���K��p��ӄ�:�����"债@Q` ��B��j��r�D�����+��L�4ș���|�T��fn�T3��N�K���s� v�4#ny�eh};�����3��n�6j`�#8�<��hyrX+�x@��(��(��<�@�@Ak�GJ�Xi�Cxf�ZR�Ko�S"��k�9�(�����rnD�sZ�O(���l;�^�N�%'�j<+al�Iq�1�Ȥ�1�>�R�2�+:Q߾��4)^6i��@��;���6.0���(�"{eW��:�����J��F�m�I�:�K��A�,�������g�$�:<R�L>�������~��X��w4T@L�;���ߍuzj�IT�ф1Y^²�"T���R썷�GYC�eV;�Ä�32���9��,��t�&���\/���޿�����S4���b�sV�/UZ���k4��u��Z� uv��bc3��Bpʿi\�E�G�_R%X�O�EP��ʜ��<�Y7��A��hr�@72��$��*�Z�������+1�2�H�E�_R	�T��g97����+�C.�#��G�F�Uj<EᏳ��'�&i�/g��Fp�"�4����K��y�˘�e-?�,����Sc�&��w%Ɏ�H�>����tNrB��J����U}�f�+F��7hS�~l9l�R����&���a�p�0�=(��e�w�ϣ[�p�E��G��s���T�J�Q�#9SNF�>��/'m�����I�⸗>��F�ઋ�c��A64s�X�~��f��8w����_Fhy~EpI�3� � �������Cr60�m��!Yܞ�w������!ׂ��N�ͱn
[FIx���'���Y�Ĉ��!r�����Pމ� ot��l�eD��+���h�T:it���S��� B����V��B�9�2Sg�f�yw�O<�������2䞯�;f���Rȑ���q��R�3T�_z�0S/����4�䞳�b� �{\�E2~�%M��W=���T�Rmެ�_�U1	�ɀ�Ѐ�`�7FP�a����"�?��`|͟2L�2���gT|�2����9|�Xn����M�Dvql���
���q�z�p��F�q�i��z%_���\�z*��^����Ϙ^^L�Lr/!�~�]ۯޡ�G��x:��k�G�~��ݥ����R���XOL���V�X��s �,��'9bN������p@�"%���b&�S���Q��Q��"������.)�ɑ,�C�Kt����WPյ���� ƪ��yEQ�_���v�e�ǡ���]nf�{,t�M�_!��H�l�
�Y�;�-���'ǫ%Kt��%�ml)��r{�U��j�ߖ�#d��d��U��ý1��k����x\�)���-����I���z������t�x6C�W�Z	!O����E`$ٽLyt��[��Ӱ���?C
_���y=��ƘƋ�_*Nӿ�bGG�IZu(R��k��bc���IN˵�7�E�*ߜ��Ş	��6����P�w�а.[�t�S$�s
l��祡�>7?���Rc�I�^���(ƀ�'2��ߌ�U�Bj���F����A�9��bά�-tǊ�j@u�v�E�1"�0�n(�O�CN��M�[�C(2I��s����z��Y
BA@Iz�-�a����8��)���LO�P��v�m~�LDv�L�}�W�]�?k�����
�Ԑ���5�s~B��#P�T� s�PXks��F/`�����B���8Xl(���"�n��a�A���35�A�(W���`�S����Qq��9ۧ��MJ�ؖ0��sC?ɕ-�d"L�i�T9�<��1>؋aGR�<��w�*dVT]R�����.{'F�y��d1NV.}���%G���W
����M����}�_�'f�������=� "�%�7�`�uq���[T��m�X�Q!�]l��f�2{Y8Q�'�K�a��J��$hnܻ�,g7ᑦ=]F���
��%-���JPBe+���G�]�i�J���hN�)�E��������^Τ��}9����\�����!�p��N�
�I�p����j���tMx��_�����z�����RW��#���n-ƏT�0�٠m�5P��qX�!�Щ*�}���̓���B�nY���K�����~Y[Wx:&�3եt)-��T<��B�wH[$HH:��G��MlI��
�VSTl����9hUaI�''��2�����h��)�.�j�L�Y��-a�
�W�Ƹ��.�miˈ���^����.�൹;lg������,`��I,K��Aw�P���QC����Zg(҉x��zY���*�C��/r2�}��b�l�E�{'
:i�w�'qa���PP��:i4�Z�Y�@��k0�DvWe��T��	��7:�$UK�N�b��^1,:8�Ф�_���2���me�u��9�F���u�$ L��S`�n��p"7'�R�L{c�9�P���~�f�	Q(�e���L��r�+�7�!aqǣ!1��p�LI��Q�P�u5��#���9���,ؕ�z� �=���I����R:Bdwe�8��V ��q�0LF}�)�?W�FI��� �G;����V�0�
ez�l.o�!Z�'u�}3�ƮS'�rNgu����J���*�?���[����!�Y!4��g�p��b�D�C��-2������Oiz,9L8|��]��ط.^��\�I�
4�VyT���ޯ`M�Ե�:��̀°^����?X�6��vE1Cx�4s�n�NZƔ�n.����4�}��B��&��V��/m�1��1dN��9�
��|���zVF���maq[��{����ݜr��0�����5Y ��*���p�
���Ѭ���eG����3R�V�R�[��z&5�W�Lk�����Rr�b���j)���ٓ�h�sf��u���@��~|���k�2&[lzŋ��p�Ռ� ��[�8G��D���J�?{4�Ç^����"�;���~���w`a��s0�St>N9�mU�Z��z�/hpe���)�ҽ¿0�� ���q�n6�$Xr�Y�_�f^�+�r߆��՜TN��Yy��+��So�(z(�����Y}D���c�1_}�&�YvOz����c:���w{3�����L��P�����3x�=i$yw�VZ���3��Į����WY,�^5���ه`i�� �;�������`��m$L�̜��L����ͷ�/c(�<@�E��s����)9�Df�O�-��{���X'��2��(��]��?�m,��Ȑ��h�]~��& g��lf�ԏQ��3�-�����=��R��@�����a�ܯw�ֽ-Nf	��f{����Y>0Qp��fE���|�� ��'��ɂ��� W�U
�Х����I*!C-�_���4��W�!	c'��
��J������C����Q�G�1^ߴM���2�Gf*�B�{&C��CVe��]e�B�bV�?TE�5�ߵx�s��1 �p!���w:��aK߁y-m��(>�۲��:�3�FY��#�4o< ��������q�u��y��m�Q)�oU�f�f��Z���9hOߛB\P	 _�AI���E�����Z�U�Qqz�GY
�c,��,���lB��O���kQ-g�yT��^G�Uj�l�2R8�Z"����z"i����pi+�cHp՘��yݤ�(p���+d
#{шJ[�r1�{����E�G�3�!iG�mk�?+'ԛ'$�԰z4c�������))5��n�L��9�z���+�ӚhZ�Z���q�S��`k]}o�o*�A���)_����s)�,�	A�	��]�m>�	�$��`�JF,"t��\V�g�&m� x���u[�6�7H����i�h�cOD �uXj����g�JY�_��0̆6fR�������ū����9����E�@&�\[�vƉ�Q���^�� >[zR묟���]z���p3�sF5�JR���x���n���q�E,:)+"ꔏ,��p���6��++���S�L��Kv!��X��CQ�!��ʕ���qcڱ|�|� �)��!��������L��bM��2s���-A&�)��}��kN�`���&��Fm�>al(�d([U~���h�>��FT�g�7U�3�M~�� P�FU�������M�1����[�B��ُ��2���Y�'���Q����Z:fjQ�.�Wq�~�t�����ѠL��VI�!�FBb�s��Uw���c9�]|���@������޷IUl�^V	u��b�4ͨN$8#�,��>X�������1>N��!�@Hi�'��g2n���!�j~L!*rdz�J)|��@�uT᚝���^GQ����Eq���e4�}�(��>�aB��y隝�[�ᕥ���^e�ȏLRb�U�LL��v]��z���<��1�8J�AE�!���`��p�?Hq~�G'p>� ���C)J���;010�\osp�����W#'{�RiX:��.HO��Jͯ�l��vk5d�T}���SkN%RM�D/O�e~�R�v�m��D*m���u��VQn"ݦ|N_[���<���W =�Ӕ��l*��폴Ah�O��Y�nì���0�Sn;�����C��tZ�~�ƞ^-�im;�y+�b(m�G6\�[k��v��|�D$�N׷�����D(>�~�����^�RV�]q��n ��ڍ��ʌ>��v4�Р�䳠^�J��%GSּ���x;\���i��\���iz9����@ 1���:j�m��q�U�G��h�IG�ܪT]ѫJWf�M�S쎣hR�^	��ߏ��+:�*/Y������D8�����V6�1�ؑb���rь�kC����B������H,=.Dms��(.��
�v��v��J�^
�F������� �/��W�>_Id��j�p]�A�xVs�7���l��V:���	3rNt����N�;���o�I��V�_��(_��s0y��'��65sL�V�F��ϊ�G ���X��{�L���o��F�׭\�:?�v���� 8-��Y�c�
C��{�s +Z�����w�hL�$m������aӄ��wq/�ܐ�h ��V�U��I#�
�!�G���5Ƥ�JqeUr\�L��#�#CV�i�Bd, �͔}�;A��Y���"���m�bجs�����4T�5��e�ozD�ʹ�k��27��c�:�v�"�֙�v�v��>7��Q��#�Qsї:e�OH�y���TMY\aI�v{p�rK�V����c����w��Ub�ٲA3�_�$h���\���`l���`c!��n:i%��e�9d�{��}�o�m�?��F�A�)��|W߹	�H��[�T�$;Ƙ��y9.���,�5+)��-V3i�I:Ε�.��0��s�䫦~e��8N= x+�$�in�Kj����"D�?Y�;�2�M�a�?��Xp�*e�3�0�2�2�JP��'x��T����抓�y�Hm�>�"�=�\��Xg+w!�%=���u5��>���`��V���f[�YK����{�����z�(�?�`|������')a| ���	�aQ4������ ;��?��у�\N��'�`�u�t�ee,-;�~=�f���W{Y�y���r]9�,P����e�8�*s�k�3C�jia"[m@��&�����>}�Hf-�VI���0���7���%���<�b-��H���N.i* ��\���>��Z�c虛�X܀I�([�@olWcnİ��*C���"��B�"耄t�uG� ^Bt~����*ŦTWmB�;�2�i��ݶ�z��ኂ:�4a����I<5��G�k)���Z��֬�}3����	Z����..eJ]��<�q�ND�be�.�-M�I��0�w�PM�k%��-"���y�nM�K�l)��e��c����I�R!}�_�('��"�E@��3��8m��������)�㋔�Xc��-��p�D�ɣ�HHg�û�G��ʯ��`����:~�A�_��&��{�� Ͼt���'!ݻ_b�?�v�.�4�m%8p�3%8)li�%�x`\m���\t��;��53�G�o��F���6�	8��G���BrNt Cʸ��"32�R�+�=��8���.z}�_�����������{��B��FE@_H�yW$5�g0l��� s��۵eo2d��>����
٪#�Lo��e�
�c |�*=s�X{=ՙ^NJ�)c�|���	�޻��e�;װתrZkS����O��r��z��͏�@ܯ(�4�K��I	"?���=|���J�I=S�\�rȵ������t�7����^��"�֝f�����yj7Ҍ����
-4�Y����S>s��c��Lq��>ز�e�5B�B��pI�2��H�)��4>Q���*��H;�D�p=o���]�O���E>Ux��>��K~y�C��5Q�\}��mقə��VwO��(�H��m:��|��ێX{�De�ɜ܋��V�yEч�0q�]S5~y��i˳�����<ʎ�!Q}��ʤ�"gT�'i;�H��f�7���w=�Մ`�xI-�l�^�J4痚�������)J���6q�O"�6fAٙ�V`��?�ޑfA�V��� ������-�z�4��{l� ;/o?��E]��X�)L�C����&�Ug�St��Sk�q��}D��4��)mC䮗�� �$u��._����0�L��a&�@+M��:1QD �z��$憘��Q�Mt��v��d޹�,�t�+����۔����N] y�!�@׫�I��fI�8�"�l���skb1I����>�o��)tx�"yzO���� E��>��k�yT���w\�oD_Q�̱[6���M5!�?��0Zo���vl�
�Ǎ���lejGQ�;�p��sz���0z�YH�>������U��c��b��{�)V���\  :w�MJ����J��)�l�����֑3{$t} y4��n��'H?�f�zk��}3����dA�)�c�;}'��,9�r�@e2�r�:O�@H�5��� ��k8LO��҄�+��^a�S�ǫ`��/x�)�Ȁ�oo!a�iM��뽴qg�~9�������W�����)�z-r�Ipv/�4�W��"t�5I��d~�*�J'E�4�	��, l�F���p��|�-�N�����[ ����k���
��P�d����E��KmLD`BE��C\��LXm�5a���̽x�5jx�v"��?L�I��R�iF ���G��?&�F����S�M��9S,�	� ��@G�j��������4���1-�!DU��}و�����Pz�Ȏ�TE���1�<x-X��+mC���h�9l�A�����O�`M��J�.������R���p��k��ȹ���k���-�YO�Q�4!�t�����C�81G\�Y�Iy�n��C������V�8<w5�}����D �E�1ut?0FW7�%(;AP�xK������`��1�E�G�o\�r�h�G�blm-pR.�4$1�yֶ��5���~CGw`ӑ���P�wF���>�2��y:ӚYise�}�H.�D0 F�x��}�h'Z	��U�X$���0iX��4Sp���}�8e��@4���A���.{��<;�wX��T.~�k���BWCm�=IBn�x��M�h�R����{C�[������ �
��%~ ��n�g��lݠ+yw���� <�Ӊ��%��I6��XM"<P�mV����nw� q�/2E�=�'U��O������@��OSt(�;�~p�1[�yi��%_�[߰6�^�>��U�!ݤ.z=�̬r�3Z�_�M[�w�c(�)=o���ȫ£��ݥ��ߑ�~F<���g>�'|oY�g�ҧի��6��' Rŷ�6d��J���ޔ��ea�A��K�����Һ}��G�Z�x2�M�$��}7��#Z��.�K1/�?��9�o�w:A��`8�T$�g�_�U/��4�q%H���2��D��:����f���MT���p7���g̝
�t'�EjN}4������E�}�mC��uR�,��c�fZ�Bq�.���u&Rk ���0�N8/�^{ą=�Z���/`�,K<�cv���Ѝ�t�&9�%&�-�}��LaP�C�v:-��x�~A_�D:�����?9��4n/zH�|�a�k���
��3z�0bC����+��NyNA]Vi��[����
�T���I�:Ck��aW�U�?��3�*b�Y�Mx�W�Le!K����������)����yӹ'���a�V�J#��hh)����b�#ƍ��5��}r��)0�[���%|�l�*e�9��y���3��v0FtC �J�2�7i/���޳���f�F���!�^a�mA�l��eg�Y?X#�ỽk� G��s�y�8��n��~��l �M/�<&['�xm�E� �}-�1�U���e�� A� w�ݝg;�J!��T��v�4�gt$QJ��̿�yF�y�j'%���ۗ�h��"���Iԑ�T�)#����,d�/rf�_�a���X��s�_��5-Q��9��+|�6���1ͽ��[�_�$��I32T�dc��6͕D�4%٦W�ZM�ߏ�c51�Q��&�H�ނT8�`�I���-����/�j��:�ݴ���1��g~X�Q�M�WT�y��gh�"��L��,�LI�o��ڀ)A���!�i��8�&�R&�������ևϮ@��VuB|�����#Li�J�<iQ��J1ܣYR�(����j΁-���"]���\ ��v�y�wg0$)jM�s\Kl|ӗNpI�\G���G7z��]�ٸ�CXt>c�M�������:�>a7q[g@%w*Y��(Q�ӽ��ҽ�VT�t-�ΰY�V7���/5��
��9*qX9��@��;Q�cdSgR��E�6�q�&J�Լ�Щ�!%�>�.���?�5������C}���U�	���A�:��[�\6o�n�\��L�M!�x�~$���"��<5n-��ѿ�#��0���R4�9t�}Y=�@l���y���%x�h!�_�A�a���*`�CV��,ׇHM�����X=A�7��|M~AWJ�B�͕F$ˣ.��M���q�]�q%A^�a.qx�d�o���Ru��R�3�/� �8Ĝ�W��L���P�Ę��N�q���ܩ-ɩD�"�zb�Xo\1�(;����,	aV�y�������9���td�gв?l�kW��ޝ��,���^�	ىl0���.��OS׵'�_�����pLZa�@P��Ԑݶ�i�jYW+C�%�̈́��B�~�tC�"��!����!}�g)�8Lb���zU���x�F^ݳ;�CS	V��o2A��+�9��i���L��($�^z�ɿ�}���d>c�0��xC�Tb$D.zt:6�����<LY�Tu�
�U���uw2~�o�Dd��0��nM]�{��!X�n+�K{���N�)��e��l昼1����i�{��W�&{0�-J#�0���G��Cy��/�م�_G�����}�yKe��O��f�'9
xg��֚�v����s� �f���<q6� v�8�ݲ%��ꪮ�E�����xǽ�|��{RHW����Ե#[J�+�+O���y�M�[�O��ǀ��P�#��h�Z�P���iT1���7,?Y,��Y����-��^�%�&F�s�������u�9��L�-ݳ(�w����ꕲhd``��zM[��Hzu*֥���/�e���hKc����>ӛ�S�{S0�}-�Ӽ}!�PK-��>����0s��^HԤ��:3>���/n7G�����z��F	}��
Ҋ>؅+v�nj��GN���"�E�<�[��Z�m{�n� �S���q�N�Z��t=�~p�/4Lm|�7��Jnw��~��NXu�b���f���ẇ5w c���3�o�b�2bMc����Cxq�@"<2������0(y�%l_�oZY��ӡa3�X����Ӛ�C
�s�kh<�F%�w�X+]��-�h�0�ymg�^Ծ�tsѠ�t���2�n�ۂ�08[���r�Rq����beO*%�l�<�a�έa�t�9�M7}���$4ͫB/��ƄH�1N�",��+}8�����F#���S�����`���R^�ב4]�8åH�}��1�ߗ+����\��D���+�$�L1��|�(1 -�>h?x�Ab%�x._G�l��_�e�tl)���$Ɓ����ه�>Je��u�9+�U+g�o��k-e�������^�l��Pf0[��~q�p���d�8Y��y��n9k�|���B tqk������}[3�m�/9��Z�܂Q�R��Z��T� ��Pn}P�l��~�= ��A�&s�:�#{'���3q���7�TCb��b	m�c��0$��)!��5��7��E���O��у�m��K�k!�L�F�i]CH�>��e�隫���t�L8��8
��7�*�O��H�� S�X�����Z�H����ֆ��;4ɴ}��_(&�尊�L�t4w$�W#J�����*��/X+d�������fK�ٞ������/�Z�R�K��|�9Ш���aO3,�dھh��*&p%6�a4j�f��4���*S^�r\��A�}�),v�K7�_X����W��`1x��_�+M�E'�Hm ʯ�Q�%�'C�(񪱷���H"sĶ��_����j�'�7C��l��曜��,�I�Cт][Ў��Q%V~��c�3�V~"�[��=��ϯ}X�Vu��1����z�7�?O���5�~�������{�_=����B���>뫔P����mo��f_��=��<̾�w��C��=���e�/.���,#R]������E)��|cx�g
R�Jt^��-�9Goa���H�֊1Pz%{|�=�A#2��*pw)ѷ�{2��ZzC���>���C+���V�5n�v�<�(���J}�{|��y��,M�/_z$Ab#?&y�{-���:W������dm${d��:�ʧ����o���_�Q�������T��w�����f�8��*�ܹ<���*�a��}��xa�k4�lԳr�pb#�18[V-�͜�rF��b��D�����s`�?�I��br�n|FX�ʩx�2a��b�(�פ��j:rP�N�F�k�6��j#���m9)���/�
׀��!�ō���`���O.m�x��N"�@\�q������<�LV����)�I��5��|��oZ��yN�nI��Q��[n�Z?���k>�|\�9�PG\��8. �x�>�g;孲hH�2���IR�g�Q<U�ףR�g��2gqX�h��(}x��Q�yg�����-*�cm�9j�f���E_�k�Lx���t#c2s\R �ٗ���S�Nø����\�;����mT�g���}�F��@n!E~�+dcqI�f�0~�`�5#ʿ4O9"Z�zj�t�h
���{�A#�;��*���%�NL��-g�_�{I��C�����2a�<4f���ϸR�J��D���������V�J�+��-�Z{��ې��[��|�������u;�h�5<�\�$_��J]~S&�GM����"u�P�
��~@c��v�-s ��a��p[��P>��mЌ P��1��G:1����WW)f����1��W��V͈�y���O�gd#�ư8P�Ә��
�7�Po��Z�0K�9w�+�RO5��-�G{H��9�F�&W;x�ź���P^��yF�H��H�5㘚�TՁ��¶���U�����e���� ���]�g�E�du/L���b+���*9��U^o�C���W`;�xl�#Q�
�!�~�z�?�=��Ԧ{=CXa8'+���a2m?���rPw��ٌ�!�\�O�e�*��-�Z�Ǡ+��^�>_��bA�p�w7:P���h*~ܩq�}}>�����~�KJąX�����j�!�x>9#_�I�f�4�w�\Ix�*Z���xM>tL3ݠ����yw}�X�o(/t�X0(V�$��s�f��Z�w�pE�θ�Dq�Fq>��?5 r*M@n����y-�ʠ��F�v�^5#n�]��8�h�U�K$ôe\үG�v�3���q`k�,���\�Ϗ�&I-��������P��h���N����J ����JO�\ܕ������EK���LX��B$�؆������M��g���&�w�}�J3"�
q��N�������R^3��V�"�36Z�{��9q,����6��*��͵���Jb�̨����;�19W�e|	8ETCC����f��OQ�+[R�;��L��BՈ�|yu[~"�AO$�u��
T�%K#���7���9��&��7�@b���
b^�k$(%�<���ya�$��F3��͕�v8#�{dI�1+ѧib�'b���;0��Hݵ� $`EEJd��a���9�Ѯ�T��a�HO&���8Zw�8� }}ɝ��� .�nFe�
��'U+�NN���ř�n2wU��y{QK����#���J����r3b�P�q%,՜�^*���e}(�b�?��b^�n�(8c���,��!I�~�x�A�m(�c��V��r�]����B'�w9�6�r��}�U֌��潚B��w����;�T�����7�ҧ
���{��f-��IYwU�u�KRA�Q|���1KG8�q��9��X\Q�^x��Tt ��[��7��u%�����L}9lA-�}�l�WM�)��\��̆�ɰ�1��|da�d2�3���;ՎX�B&���s�KL�1��T�z�Z�Y�Z���-p���L��I:T�r��w@�o�-qzt�-�zeq�p���`I}u�l�[�|<~���sRP��I����|ɸ�I�vm�B�����t��f�
��J_���$ȉw��i���nA�U�D�}�]I���Z��G� ��;�6KC�h��&ƈ&���$4��dC�b�<)a�h��(���?뻍~VV�9@�p�/̖�I)��;�Hf��)>��bU�Ai������̝N�y�ҤY���tTY�$��O�q�����pfzb�c�^:���]�~v$5Dl�"C��R�h����C&�" �O��&�vk�����3���p��Av����8� ���ǎ eZ�5��g���p���踒�V���#�GH��{9�4�X��:��'@�������R�����u>���I�}Ǚ� �;T����0tTah�(QS��B<�(RY��{X�%a�U|Eܖ|���"g��g���>�8�5d�}{n�I���&AkZg,""�����MT<Hd�e���cbʷFᆆ��J��IA	��ߦ?;��f��7������q,0���!��&�}^����%�Y[�����%F�:�,4h��Q��-�)~��8���EE�1�z\�����&�b�ݸڃ.��"_��P���#9�Y������9�^ַ5|���D��[L@�P���zT��"/#�RϩU��A�����E�y���g\6�cz:�M-�M�a�h`�S��&������
�+e�W��<ٔϝɯ�s������!k7�9�a�3�P*V^RNk��Z]B���p��͋��O�`��l�ZG٧;uM"9=��K��j�BY.��\F��j�F3g�:9�����CR�HE���!t�ZZH%�[=!`���xZB�\�o�Ey>�����Q Q�42\�Y�	�D(�qɯ�ȥב՛A�B"��Ж�DP��tJ��a��J�'7A�w��T0b�?�Tet���a`�z�´2%C+��С����]p�\RC�'OwT���8/Wj��>��6�>�O��u_C/&��=�"��=�0o�nיz���1�l�C���/�T�4��O3,c���xD��V�]+��1"����q�
#�"��kիww�ZH�G�}�6"��Hqb#ua�x����قj֟�b�2X�m���>Li�e�D2�9�Ql}�|�A����-/�}*}�}�J��6KL
�ih���k�mSt�,SkRs�(/�\Nn�כr<vx�_��>�v�%��� y��ˆ��L3;.��=��{7������D<����YJ(��(} Ǐ�H+䬗BZ���_# ��vg��5���