��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ���������	���u�hώ�lvNH��3�z��$�m���)k�\�礇��Q͂E��,v���"yԝ�+v\�!������M6D?Gƕ7��^�$�w�(�E|��z3Rp�PMv�0�Y�n�0��yOp�i@+��5]��p�޽�h�/�@������l�ݥv�^��~h
�87��]��!A�~���jūG,��VF�.�<1Z��.wH��o_�,7^�p���!���y��5���+9U_�V��+������s�H6�e'^��K��6*����ѿ�x^�p����g>� ,IWWU}�nCo�U��U~۩��׾�yYg[L-��S���#�kg��A58��� ��/m�W�S_�:/�G�Gk:�5;e�#2���)ᙉ։��+���6�>αiE�y|�"�k�9yp#�(s�:'�e�M���Q�M2O[���՟��QqiM���sɼ;� H���4u~L��+��4�P������g(���lG4/��w/y��K]��`��Z�%b�FVVW�Sɏ!O���'�����L����q<ɿXhN����,r�r���l��xv�E5zs$� �-uJ��1����NE4�up�2"�Et�(Zd����'_ǚ�9Pg��'b�;S��1C��]�$�7wJy�4��Չ`����=�@%>"n׈�?ƶM���6��5�)��BK�ĤU��M#��6_r?-Du���b�Ee��.n�vYNէV8-HVn$��}���>�v~X��i�4�/sÏ�U�������Y|[u؋S8G	��e��;^��yk�[�7��Uw�Y��j���PX���4Lǎ�e�*�6�ni%:!k*��Š�%��D_F���阩��g|�)��I�/�c�t.\s5�s3>P��t�y|Н1+��'"̇2�D���|Hթ*Z B�*L;tYώ�-ʍ�I�mԇ�,��{ep���3�RW�w�<���u+p��~.'�Z��^�Y�m��P�-ʤT��?̧�9�1]G4~��p�J���%�L�,-!��lc�9�'���k��a� t��̝���93�i`�����5ŋH�9d�^�hoj����/�M��g�D����(V�e �g��>7.⟃�A���Pg��w �~������2�S+˳qO��z�S�����d'�_���T��Y����`�6gMUPs�L�M�)O#@i��CDhV⻈�!D5�5$�����|�"�e��+�r*�@�=�w���&ĎѲQkn2l�Sb)&�HTx%@(��F�	�v��Ւ�q��b��4��K�cy�}�)����%u�& Ts���1�����0g�]Ȋ�x��>������̊��$���~�Ti>��M���]�:��sXR�v��W���k�:�3���0l�2K#-E�K�,k�u�	���K�o�G�J�8Iۇ��ifrNT+f�:90��]䊷�����>=z/�6I�d��
�m���(���}�fp���qw�'�P�Ha0.�~޳��|�k��/E�_u鴂2Oӓ���<W����@l3�%�/r��?�&��Ug��C�Nݤ�";���Z2�?�O�0�B�'�0B<�΍�R���0���J#N? �S+���C�{T��Ty���ȫ��:�
ݬsfv}�!g�E�֣�U���y,��\�����b�;
��)QYr���gd�p�V���_|z���X��(�6��Z�iH,�t�{�s�m�XZ�P��U�>��.���+�!�J��t���_�A��:x��a��Ui6��I��k�,;;$؀��u�+�R/KM��ڑ�����t!z�9�FĖ������ojP=� L�%��Ρ�p���DBuч���$�׾�uMf{Hܟ��C0O�6��\�6홎؍�:����;va�R�)�����m���3��r� :�u��a���C���*�
$�#/�r&�d�/�+�b�p������ר�,�O��(U|�4���ԡ�T!S�-[���ܮ�4�g�LՑjE��\��DY[�kT��A6���L}kff\���	6�u|����%Cu�8 0�G�Rѭ(�$"K��%���-��u�Y�"y%?"�~h���;�O������~Ǣgb�<��'Su�ޗ�Opǭ�(ZT���}����(Ac��a�f'p��PR�����ߓD�� ��o��?ԋ�O�p��~fE�s�T��JQ�w?	���80�N����!���<S���%�Q��<v��W¾j�U�RD l� �oH�ڙ~��|	c��� ʷ��ZF�����f"J�_��Q;H�wDHGU��M�����i�6c��6yR���,�m:ul�`���d����ե&n/�MXY���JLA������~�4>6{����b����l�(7I��9,��@䷶��ʥ���;�AQ���4�v ��5b����,����rT	��(5�Fƅ5H/�۩,���V�#���L�J�����$�fb���&�js�Q��1�,�����jCVC�'���B�~iU@�����P����o!�/G@��u�T�w�v�2F��v`�|;{d�S�d7��3�(�
{��sP�a��x:�8o8�����@^��ME��1ۉ�{N��%T�,���6�c	?e�Ȩk�y`�czA�P���0��sb� ��]�Y?"�K	���sk�SUhK Jjș�FbA�9����>�g%^�_n������ ��U+��[;�ѣ$����G�Q$�q"�Or}p�ɔ����Ry��ڣ�����#@5���'�v�F��E�ů�!U�\�f�Y��6P�mw���.�r��p5��},Yp���m}L�:�z|F�NX#3��-�GA���"����0X�8��B��hH�{��HT|�zeSZ�P��N9O ��E���r�"`~[$�h��`�M�X�U)��zʫ?�#2ꡬ��=�aP����{�73���t��TӰ���ԕ�ց/��$� �$(�nڲXiLo�0p�ڞ��h�W�\��T�B��<쉯W�.�S9u�ڋX�d��X:��kW?~?��;wGe��эQTȶmhAъ��S�a7L�B�i�\,܀��Л����غmdqX"m���&U���4B"�g2�������\��f;i��B��=:�*��7�&~���]z����7�[I%�:aǱl��^Q$����̾¹�}���[����B�$@�X�������>=b�<�p�d%'�t9��Q3��9���qt��e�+0�yп�3̃�O��EJ~s��6��,��c�C��=fHeBjL`���G� $J��Ur�S��Ti�0��:�~�S!��Z���kŦ��p��F�YV
��[q�R����k��@%f9�����X���^.�f$��Z{:(|��3�r%�a����ɍٕ��eQ�J4��B���9��K_�%C&��-V����1,�\"=�����;��(�Η����C���r�U��x�д���S��HV\rk��m��C<�	���~��"���>?֤���Ԓ���ֿlM�T7�(N^ ��l�qnIt�jA`5"��/'�|�1A{IK���>�l#&p�2R�:0��b��|�/��v��_��������s�*a?^�bj@�o׀�z&ɢ_�\}X� G�d�c��Z]�ğ����H�1m@Q�)�!�m(R�`�7yT�WH�m��� (�1]D�#T��]����bs���ם���wۿ?��4�X+Wu4=͙Τ�VI��~�u9*�����V��_�>�N~,�R�|a��9bR���`�2���
Z௿�ec x	����~���z��;bim�hO<�̛�J�-�a�?�կ�[�/OC �� �-�c��|����3è�����\��vd���B�&F�����0电� �/L��͝bY5���%��;o�����ͦ�:����.�Cq�{t�ИD�O:E�?SB�)6p4�N1�F�/s�X���*�rk�M�#C
�(^��(�R~ߔIR!ԫf�H%b$[ WΦ��ݝx��Wi��/lMY��~)&W��̨B�$! <�'�XAC��91S������%_�	G�v$>�zb���!3L�ZM_r�I�������lW0�?�`��.T�I�%�����\m�%�~�[w�	���蹜H�ᛍ[P�c�/#ִ6X���%�X�&尶��Kƨ��Z�ϛ -�Y��j��gc��,7�b|"ł��U�d[��)�M��#{xW�9n%PR�+;��wD�(Ɔ�L[��Y��gS�ONS�ŗ����؏'�hΩ�����
Lo����y� �~�"��Z;��j�uO:0�P!3��q�M�V�%�	\��T������t��r�o��*���2�#��x�j-��C�[� �%4� �\c4���nu��`XA�{�ʧ�S�+��I��0{n"`���9�??:�:sq��lWm�K�^K�T����UKt�C*d�Q�r����`�����.�p:�+^o�1CoL-����p��}&�2�gSj�w�%7m7��1P��}Dwa��WC0�怔���T�C6l�k��b_n���2]Iz��F�f�`�2�^��37.�B\4��X��,��=�ҹ�F�ymkz��}��0�[،�)�7�y���=?$�������R֩�{�Q���D&��=T�� 
���Ӈ�b� _3�2y�t���ϯt��@.��٢�'���O�J�����pJ[��'�d��Yx�'��MT+��-{?�X<׾��A~<�TƼ+T����;K\�b����,����F8Ӎ"��"��?%f�m,��{e?$�7��x����PL�r+�^�@�2H3X�;��.���O�<�����
�u����ι�H	,�lLX�ϣ�AQ����5�z�<f�:q`�)P�"q�ia1F�\��-u������>�IbV`�C�{�5[L�2pSg�]�S���q6)�o��������O3o4�Ȏ�[ٺ U7fz��� ^��H)L���+�ll�l�'��~>�U��	�����o=������A�P��z��!��hQ��A�Υ��_�,w>Ke�ޜ�g>7»�[f_��^n���iD��=2q���B�����*�v��"���j^͔9
��p=��#����и���m<��E@��Y���uV
�ge����MȦka��RWT-4�����^L�.���گ�qF����G挙����P�sV��֩ziU�?S�Hr�a�9
�|�Qg�c�ǢU�hߖ��M��P6w�_�ř_pT@B��p���ӃkN51��O@]�!��:���!����CvΝ��p�S��\Aㅧ�����հ�&�}�m�2�Y9�nE~�" ��+J�=�3W�_Ԝ�A�(��*u�[®ϩ"x��ݾ{,��f��UG�g����5�H�(p��ۧ%�҄��� ��C)%�n��f�Oy���lϺ�㑥\���d��F�#��q3��s�Q���U`嚄F菠��4%�*�׳x�ݾ����>�u(�vۃ^�=߽˕0�S����ĝD���p`<����+��QeT�6�<#���V���u�ac�B���(�Lr���&�ĘK�!<.�j�c�X����g��	���>��C8�����{��zcv����[��W�p���v顜��,*�#bI���`�FC,�:{`��g6R}]&@�sf���r�M�� x�d],;�mOΈp}D�%^���3I��kA�����J1�w�2�43h9�m�#d�\�Rr�8�%�(��R�A��m�MX����	�#�!� �;���k�x���"+�2а{���'Gq�.��=� 妅�OZ���󣭽|酑�+m!��U@(��"q#"z�6�&����8.�������D(��t\�����%�{U�.}��Ԛ��Ke��p�1����o�<���9��z���}��D;A��V?1̿G��A��9��*�1~p���6���)o��3���������P�l���,��!_T�zp�i�S��)�Ze�
��Lu�q5D����4�g��-6��?�A|���7�ߕ��#�#ڈ�w�����~�Z>��íӶ����5�1i��@3��*���#I��["Ϧ�Q�B������ENe?����&�R!?}��b����x+v�����s"�%�#MrQ��6�֘�!^$�����)XNs�~� ���Ǯ�@�{ʘ#�GB�%�8ZiSP��	���=��.5q�a%a�e�'�bȨ�#C����E}J� ����-yd�&�Aّ;ġ"(���^`����������=WaP8��
�`.Ҍ̭OF�ׇ�	�����	�b��,a���ŐP��b�R@�����HUᕙ*����O(�Ļo��$����|�6����uo�+�K\.����1��	�Ц���\�8Z�LY5F=�/P%���l{Gf�Nl���M�
�(�ֽ �#s昄�c@�>���ĥS[����)�W1Xa�x�e*1:�[���'��c����@ɦ�m-��D��G������q�B��*�jQUeU W�uM[�:G�b�f��g����,��fb�8Q7�hD�%�v��F���l��\�PC���� ^��~Y܁��2�s���|'Ӌ�Ic}zD@�$�����q=����w�d$�Q3�Ȗ}�v/Y�
�wա(Nm����a�1���M��.L�A��W{ob�2���Hx��#Bu���t�r%`�m.�����L�ؐ�׶ڞ�����8'aNl�X��5���fΑ��F�_�H���m�(GKt_L��[�f���Q�6z��t8$����;��/��Ub~�,WZy���g:�*1S�F�5��z�����"�$����"6�V�<_�5�����Hͮb���6�9	$5��v緒����Ã�� `GL���N�����X\�/R1�\�ghr�����OnF�'X�����S��ρ;*t��[B�yW��mvvM�k��P͇�@�,G���Bܷ�HU���ދ�5�Ъ�ӈ��#vE�N���D
�.��Lw2=<��E�{�X�8P��nK�li�p��dW5�g&&�gڙ%{L9����w�nJV��"F-&P?�Y�\�͈�O��̍}���5Sw #��o��2��Z�W�v���$����>�JY��w< 5<��9n"���]�rގ4v�2̩��!�w`Ȧ����mV��#������(���V8��S���-��A��%��ae�t\>�RG	��R{��\6��m���yء!]R�}0��y,G�9Z�W��$�#&j�i�~�͞/�[y�S}�s=��\]��j�k�9ƨ��9	� B���B	�Qk�)NM���K�����x	���t�,!*���T&�[Lďo0����T��(RGf~S5�f�l.�)���K�#�b�ǟYo-�>�b����;hn6岴�.����>�ƥ~�UN��y�@-�翨0.��;��#kא3LK&���
�R�k���;E��@��|�
 ��V��I׆=��]���:N^;�F�k��&���̵`���9�k�*�*�{,=�1�jS&��Hܐ�ah�ŀ�M�@d�S����ۏނ`oT�>��Ō�0�q����|�-ZCo�b��
񂹩q���G�R)f�G�!�"�W�}H�@m�BM΁}�9uKu�Y>�ſ����D���D�����l6|�ꏔ�$y{�{����4m��i��j]�Z��_�qr�%[h�􇕍�٪�g�ܞ���JD���0SRB������|����]ױ��Z����QP����X%��OHL��I��L]����%`ŝ�[=�I��t%��bv�h�I_5����h�Z��XPp>���X�߸�HY�T2aHI�յyV>ʰ+�9y�Q��r�r�K_�k[H>���BJ�?$��7m��P
+Ŕ��t��g;�RZ�,���b�}Q���&�}�ء�W������R���a
-Pz�D6���t~ە_������#���yd���m�s#�)[�dg,Xam�x�����WةX!�dCo8�/���h�(�u�U�ݙ�r���߿�_�J����e	M %0k�աg�km�{�mE�P��	^Ƹ���1�@���X�Qwt�F|�z�.Z��Щh��E1@�����V�{ءۏo�<iu��v��@R���S̛(Ĩ_ӥ�0���g���m;��G�����!��v�E�#}��<�z��#Jv�Z�Y���I�&U
����q�Lm<���,�[h�R�r�AK�]N�I��9�t,@�=J�`/��a�W!?�q X�%P��'.��:���Ui3�ar�����]'�Bs�����E���-�@T�������J��6��$�^p�P�"n0@�������� FF�J3O�.d]�$[<Ũ"Tz�J^�`�n`��fm���X�SaJ5C�hn��Y#�s=��re\�kr���?1a]+�ƾ~����|���C�Tt=-	���/�Sj¤�G�A���(ah���$1ۨ�1!3����N���2`��~�������e�H�wA�����Q�S����#��+t��'�K4��a=�1!��?U���\�#F���_�o?9eߐ��7j½zC)����u$]�5�Y]`L�ړ�����L�A}�G�B7dX���x�iG��d��a�3�`��*��]�jc.U1����(�/�)�!�$@۩tɧ�D?blj4�N2��ej��#Y�r9����|g���d�F���s�-I��(��q �A��B?01��Toڮ/���1k�>0�Z��b^����M���k��}qg(h�ӷք���!�D������8��r����-
�� �Ka����6�3X��R`/Y��MD���ΉKw��N�H��Z�)lw��kO�|7���y�>��|A=��v��O�{'���<�:3s<��.o��Ue��]B*e���b���l��]�����\eO�3l����r:z�
)6σe����� �D�]%���N�R��,��1��bf���\$Ѻ�����~�1e�p2��>�s~|�"&)zC�!�&Hx����}���	?0�:�U�9���>���+�/P���+)���E8���|�Rj؆�KL�U�TҒdd`#q������jk�B�K���͕��)�{F����(G����u]�,ިΛ?v ��TSc������/��0���
:%���u�9o��{��v�M�P�Ƣo���B��F[S`��ir����.���Ð�0i�4C���g����Q0ZM������j@��s�U׍�}}뻼�k���*��X��n7��P�I y�ą�f9�c)]>e�� e��P	yYP��u,_�M�B�.4	t�L���f�O�WJS�G�j��i��;.�,�:p�(�����ARdK�3yI#s�D���B�ɥo�B[nĭP������C�C1Z�y�u/]V���^���f	�-尮�EQ��
���w�߸���;XU{�Ub@}OX���U�
K��C���$B�;�!�>���1�W���l��_��tM�A�EjG����d�4Cu�d���P���tӦH3s�<�ަm���x`ֻJs-j��x$=@
Ѻd�9�/�3�?WǅY��MN�*��f�
�<u�ܪn�⃖sU��� ��"`4������ �\�H�i��d��b��$؀���}�qR�J�ִ�|�W-��B��%U�� �c��[$�\��Z�-�bf���$!�������a�n/W�rz���Ҿ�B]�*�&���ϊ79��e��>�M���3�~x�^2�RkM5z-�-�V��=k��n�p��,=�]lڒ��n���Sq��oQ�az(:�=U0������Ο��u�"�6��_������A�+]'�~�����B0��+��)Ig��;Dzra��h�k
*��'݈�"��d�{Tbr�#�;[�I���A����ľ4Lf>�\���;2"r�l�p�.���������v[훘ǘ��J�q; [$7�sC���\ �rZ����K�0R�HY����^Xz�Nx�W�Ll�x|Ⱥ��WD5�,;#=���. ��,�!���b<܋qN��&Dk���4b0�]W"ڭ�L�b����.����Vv��Y!0.H�̉�'�H��m'��|͚M�׋	sc�kvlN�0�_CAt 
$�W�(�lȈ��m-D�d�+�q^,���֫���k���P��߲ ݶ?g�F��;�Xh��6Vŵ ���H��([��mw-	k�_\hU�k�VVq��u0�J�Y����h� ^f�%��c���<a"cl�_9G̜�������P)�&�W|a���Ec���NPX��!)$@��*�ӄD��������8�xv&�@!�9���(5������!��:�ze3���{D�;1ra���� VВdbnQF��G�Y�LH ��az�j]�K��x�0j;{]yu���L�#��g��D��]�����5
'Z���>
���c���~�����eӓ�������_9�÷�����p`�O]n�]�g��5�|�"B2����bD��M���(�h.��1w�=����nN"��!�?ۏ�k\l����-Ja��? ����Hۡ���'C�����箨p;���>_���f�4Xv�½�r6,�e0����Ak���?T1�	HG}�|�)5ۅ�R������²�h�tZ^yƻ'�t\�;���l�Z8sb���T�4G2�ԢNk#�4�EB[��7�M��Dw6�z������w��ԛvz�}.O�w��i_�n����-��za�(����L�	�×� �����θz�ԨX��[9E~$�q��;�:w�D��ͨ�oN�K�\�H���'�<|���S8�`����zG����]A�M˽�����i]n�7�f�P\fGY2�6w��.�`��<ɏ��Tl�E�cS�,��u`Zc�y��~�bC���oe�}׿��A�wWr�C��Z5�����T5}u�P�L0��ۑ�2H����4
�vb�E+W��{V]r�b��Ď��T�Kn�0��@y�!�k#7�o��ZG>�ZWǕY�<�8u�V�ʌ�c�R"�X2��~�$[�R�o��ލ険�w��6i6p�u�:^���ƭ�fa�bgك��f����|;կ�]��V�d��v�(E/~d�)4Ɓ�`�Ds�L۴/���h�Js7㷹��Qw���W���x���ۼ�!=?��@���9������6����B���&-Ls��:M�g!Y�e�I��9c���ٸ�Dɾ�G"��U�_��5T�\����2,j���b�a��T�m��{r�:��uG}m����ʳu6�I��k �2J�!�m��?����(����i��U�e�xe��1��Y��`n)m��<�va��zc����Z6p ����Q�0��zI?�r����b7B�F�����hoN5��1Ճ�����෸��aAm{;��W���]�ZA�X
|��O�
6ڇ+��>Uw(��+4y�-}��T����j:���9._�ǫz���E�S�?^dC �vj?&):9` :�y`�"K���TO�KS7�k�9�n��k
2g͝[]G�]�O)O/��������w��g��N]8;�%"���ⲝCXC�ځ��8f�C�|(��ܜg�t9�n��)�x�QF'��s��C���'����E��ص<�Y��$���X	F/�������@��\�:�xK��$8`N�/�荿s�6�4����1�� ��9��q�>�6:,,��j����-�]Mk��~�����c�0��x�v�^�b�����Pqh&O7�!�ʆ�N�f��6�>tWR����e=X���>t�\��� &��$��7���֤�/(��:�MA"Os��~�2u %���uv�p��Q�}i7���e9��i󺴭]��ȶ��������]�=t;���J7T@��x�8;�*�CV?���j��a�{��ȧr��e��ˮ�Y����!��u��ͯ~�)�
7~K�/�W�I>��E�I���a������6>�/3|Q�j���V�v !��=�J��n� ��tsh���O!�R�^��v��/G��b��!PG�~��\'dY�r>F%?�ՆmIb��R�'�O(U�������?�h��	�\ߣ�A����?�-�A?�6i>ttQ�%���p�8q���
���_�%vXa���[�ʚ����,vU�L��6#�����E�&}��]��N�
:���oG�Y����u�vv�,�9y��>��+��Bx�,+mG2��ݖ�i��qZ]��&6f��w��q~�Ȳ�ޒ\����\s�3�^�����Yi��ًcph�C�R� a��5�x��}>����ș��1z�d��%Z�ţ%ɧca���{�o^s�?by�x�`i{�� ����|�mk�5KP T��T���1F���u(��ǰ;�b�y\�2I�k�{������u?5ܘ�-����W)�ĥA
���t>ݷ���:qZ<j�z�.=^ǰ�>��
����t=�_0)j�9�?����7�=Ӛ#?%o=�F,�P��R�S5�d,N:C�Ѝ��4��h�Y5�j�'k ���	%��ω���{r@w�F��N�!9ø/�6n�OI�w	���^T� ����X8�BȢ��|
��Ol�+ì���� �����Θ
������2 �S�f�1��I��8hypB�\�1�d,^��i�8��抵��U�2ͼ
�~��*"���8T�m
I��Ծ)����Ԟ�X^��r�1o��6���iF(�� d�
'j��8� �x��4ȴk⍅
8t�m�@�dn��6����	��KB�pWQ}9�46�M�ޫ\���k��Th`��,;�VFri9C��r4!lq��ﵜL��|T�^�رr�]��P'D6H&M�����[� j��Q�����k�$��#X����P�Z8�� �9i]��TlCs����\3�v��A�V�WB�;�� �1������
�v�L�r!��ؠ�&Dh��҉���g�z8C2b�C4-�)i-��1).�S|gQ|!�7�r���ſC�ǭ��J��4˜���@QU�� Gk�^Ԉo���#�Pt�������F�/df�,��.ݛmOY��~���0��)K�9H�g�?Uk�[+�Ĺg��/�k�yE�P�&Rl�K�d����p^���U����!dTh� ęF���w�g�3Wj���F�%.s:{����,�?��]<H,-�$���ȟvr,��%����[`���Zga���&��i0��3�ݲ�k�]���I.n�u��H�С%lVܭ��g�05y�3��w�����{���#el�<g3�ܰWV��a�O9~
�(��-CJ%ϵ>͖\F'��
>9±P&ۉ E歴d�Έ埘mnC�F�x�R�n,���Č�����!7�/���3/�!�D�����z�В�H�x`? �>q��܍���p�����f�ʏq�J�h�M鉛�Rtq��I�$DE�P�Ws���\|u[D��T1$L�=���
R�g������?��N�����/�:9�� c����� 
%q���. (���U���iG.�P���gj"�/=g��F{c-�Wɔ��0B
��⽧�0��(|*�q��L��X�l7�:���(7u:>�g�����==�������r��y�H�P�����KD���������gNV�>� P�� /;���_�`iã��"��Yɐ�ʑ�ƍ-����J8���-��T��`�vd��i�.�g*S���@���H(�t��I����I���}+oy�U(�~ϻ���O���h �2
��4 
�P�JE�	�����Ԯ�5f�{^��i�`��>�s:v�7H�
��D�3	7+Zc�%�O�J�J�2�)
|�-!9<+����DD�Qk�#�2?NJ���u�՞گ��?���Z��R-�d�A����"Pԃ$3o��8�s����Gj��-,Aiv({Av}\�����5��|�i??��OSm�Nc�v��$�� �g�Z9�A�������T����#��䡬��Wd�,F��a�^t�h�W���1Ȗ{�F��A�  E��{����J�h�s�������x�s�55�R3��|o�5�6�Jфw]=c֝v}՟�i�]�F"%�4d"�B\���<i<�Ґ)��ǃљ,�z86�����7;J�b�.���`��~�p�� ��d��'�2:�-[�ʓ.��a��>��r'<��p�(��c���M��2l7�dN/�CFc��Wa���N�����+}YQ����Ӷ���C�*5�8��s��=��Vl��V��蓼�s���D*����Rz�y�' �z�#` jU��'��+aOA����χ���קɛ����gqI�3�D0�d	~��{�k�a�C�:�?>����}���Ȼ�yx�1��-!`���V���=2���i�@f������3w,�)��)@Z���^���(?O����'��EUg6%�y����HыjU<���[S�O��ڝ��1�k�j<UU����e��=��w��M��<
[X���nm����!/Q��b��ec�d��Z]�����]_�F�Q�·W���'�x;�O��yԌ ����ȇ�u$��բ�%�L�_}?�/�5����]/��P��G:���"Q��3�!�N��.w�)Yy��Od[�ht;�-,90ռ[�����$t��Fj�p�`ڲ��H\�6�=��t�T7s.)ʙP=}���o^�,FAQ�jсrրBgJ������wQ&��28%"ZK%�l��3;�IFB���l�������|M�t�[S��$7dt�s(k���{�RK�;��������A���`;Ŗn@�A/;}�K�fɳ��`X�����,�|@�zR�cU�Fs8�ގ��:���}��}w��Ѧ�',k�0N���<f1]���i�6�w�xlb�
o>}����+.9���~<N_�W|P+�~���q^����a.�ش�D�T �Jf[kuju�Kޫ��4�a��ui�$�������A�V�kM�M�&��O1�2O���&Yv]��޶ߣ4X�M�A(�4:������'�K�U�Bu���P��@��=ҷa��Q��i����6�,[��A
	��)/2k�+�J��#�䶓�N�1���O$�ؐX��}6p浴�萤�$��f��q}���}a�#��Q�s]-�t㿵r�>���q) '@�;9��)6n|��rٸG����?�����dt��%�f�q�����7k�^0���:�+���E���n�������*�h��|��,3�����X�O9�4/��:E9���&Q`�@&���t��0<������O-Ro��ɤ���k�78�������� ӷr۲P��O�u���5�-6�S����360uN{]����q{����vìF-��_)�{��ǀ�x=�V8�?f`�x��O�����ڢ���SdC�7l�"� ^s��-�TqP�T�l�E�����'��ҰfM���o���%0�Hl�7�B�7�L;0�E�đCc��,M�XP�+�FqxX�#��.�b���V?�Hk���f�ue��vju���7��C�"۬�>d��v�%:_� ��]m��
zl�'�-���3�t2HXj�E����&mۆۧ�9�[�0�M�2`��d���=C/�աƠ'r�}�z6t燔�dM�v�Y��� W����xG��c��[K��D6�����w���~ٯI@�E�,�R
�z�3��B�u)oh߳��)oU�?:+Me a�T׉��>���7�/`������@�?p�B��WH� ��*S��a2�*mw�:�/�����bb�#d�P�YA$���r���M3b�5���6h��v����9y���ֻUH���)��1�+�S�b�/�mG9R^���3�tc73i��4�V��J�
O�&JRR��Kݹ�>���Ghrp�MH��E���.��Y�0;ԧ��7�'ѫ��[rj���B)]g�w�:�.�ꁎ��r�X�}7f���t����A�b����-��T�he_�|@s"JI�!Gg���y��q�qs��j�9� BTF�G�q�G�%� �]d�ѽP��ƫ�A�W6-5��Æ�, F�eD����͘�>"i_���P�g�|?�.IH^d�6	���.���;����T�x��@���g��Ϭ%��C_�A=l���p�m�����TeLZ҉?G�lA,�C�	��f�]��n������͒&�*���ǰ�_�;u�����J��C�/���h2�@� F��E.5�B\E4����Lcvp=~3��0���FNk�g�Vm�N�
~�Z�I��S�����:��qBA���~���Oؑ7,{A��W��b�TH��"?��?:�`}\aB����TM����9X���3f�-��3�{�����N���y�7=�GX��%~}(��@�0`V��n5�^�ƥ$�0��\��s��lC��c�(������/�EM�'� �Q5+���A�w�wgOx엛��J����U� �z��V��/PA�	� ��K�p?��*��������l����ԁ7(U�P��os�Zwc71^s?[�}NK�Q r^�9���4O�(�1�q�\�10�+n���0�zVb�v&Qq�5j�?�Ф��1'����T�#�0��]�\����g)Q�����Z�A0�]r{��IsX���!�b)4�h��H[Y԰d�u=���hpn�T��Z�~�?��+F0)��EM/��̾�L�s�T���P�?n�� T�
ܮ5��6?�U����%��'m���	�V��}kQ�ez_�G�b(�Xd.��;�#�
�]ܼ��^7OcM���1Q���ٵee^�'����2�#(�$��߂��H�i��<hיj���'O&d�"��;Κ�gڣ=$#ܡ�ر�pٵ�_Nϣ.~�e=n	ӝ�F�	�}S�O;�;��ɬbN��_�!���Z�5g�$U�0��L{α�b)`��Sҙ��ǎ�;�O�q��gĀm���n��IR2n���IR��Q�����|����8������Z��=�P�s=�w��p%N��,Iq��c���P����c�H�M�[�X�_�#q�Q/�v�d�A��%��(aY{�4������ANc�$�}�,	T�5���	�Hr��J��ږ�gn��WL�����Q}����{��������uL��> ӧ1��+���0�d�!�g� H��XF�V��!R���w�Qq��zk>��8���)��j���*LD����0�I)�g��-���=�T���A1̍N���#(L9O�7ӡ����O��Qv��`���F�y0F��7w|e�;^>kR�皗�L�u���	���}<�a�^;��7�A��j�C?N������H�*3��=k ��^='~8g�B���P�n���}��Kw���1֚�`:zI�|�e4��i�s�݈�g��g�/i2ȶ6ǔw��~��;���l%[P�J�a�Ǧr����J܀ȝ��T�۵�_�4^/YQL\LYDT��H��$d �E��,��ɿ)���'G��&h��"�����n��&��,1U��V�����G<{���ó2�Q��,Lգ&�A�	*���$��S͵�xKwt�����ZnD݀6�wN�9� ]�,Ը��T�T�Byk4�lvh�WыU�`MϨ��+�C��G����g��:��Ku�"׹�r�mX�W��$��������2���si��57��S��m��L�0wdt�Rai*Q>��=���	�Â�p���`�ԙ'��$�E�?r�2`okb�q<.��9P�tR�CR����'Jɿ]���U`m�Iӭ�����YF��2�h5L�����J�:U��}b
�}�f���Ϛ��ğ��	X� �b=�	�;���P1;Ï�ֶ����<�W�' ��cM&�˘c;�`UA+J�B�v����OY��SItD�n����x=
���O����hS<�F�㸧���?�B�K�s��i:�p�/��D��@�Y!�����Ǩ�8��}�6���#���'�@� �Bj���&��-���)�F�w�$���z�4Qo��a��|�X�>ry��ʠ5�{:,�!����J�`H�n��0Nu�E�,�:?�-Y;�}��3����u8�rFd#<.�R�p�q�U�Ȇ���5�}�Xv�f��q 3|��ոZm ��4�^Q��Y{���{!��@#�}	�\��>q51;�Hgh��=$CÊ<��q'��/PP��̽*��#/����g�gG���A�oL���6�=�:��YS½�[��;m�LAh��Ty��H��'���݅=u�^����4�D�66�VB̞]Y��<nAsyUhGVy��a�2x9�p�0�З��OxF=�.(8��=J{g�F/*'���\�J���Y�\Gp��V������#x[9 �cY�k"u0+F:�^@l���#����݂�b��y�4M���"��7G�q�6��ً3B��6��c�����)���������3X٨1a`�Y�c��"E�&�L_�P/B=&NРշ�*��ׄ�2l.��n ֐��#�"�k�N�ۘ��W�4%�����('!�\� �X�w��"�֗!�X�-�u��* � ����
6�.��3n~��|����ܸ��]
.Wp�N���F��G�g��S�J�P��%�a���Ͷ캇���t�,/����?��-�u5�h�]�L��Ck��!�ɽ�yA�=ݐB��D�J %��*R�����H�a��g#�U��Zn���V��]��;�y�K�*��+'�^)�e =HF��Y0!�#]|�K��
旲��v��=hp�/:$�������2�u���rZb���_��SC�y�P�ce^����~윆�^{_�1���ʖ�Be�Ahc��VxLx�8��E߯V�m�fU�?�6�F���J5������Ǻ`�쿂6��ю�S�@��14o3XtE���Wp�uP�R�SiK���D�M �����x�������
���N�q�`���*6қ<o0_�(��~ �&�{Hw4Jg�Y����q��G��n��ww&�}�;���D�2��
�=���N�#����Q��o�ـOr���� ����	�Ձ}���4�Z\��j��lnT�����FG%�$7z��	�vn1�U�]9�:]����/�S��W���Nxq���Q����L&����+c��/4UU�&<;����U���!*��U��,8�f�ߪv�d��	T���D�:.��� ϸ��)��r�(��M�Aa�[���?�V��0f%��ڞ9r��ļPkuHI���9qLI�zKR#=@�2�Z��)��3��쟵�6���4m~T�#K(��P˽�x[>�t���lY I
g40�7ǻoo��D*?؈f't�YM���D�^�9�_�Ä�#�Λfo�w���;E���ќܦ��4��Qi�����ZJ*��	��?;z�&�����[�J�C7���0u��X@�Dϓ��l�!��k7p �i����ځ�
\=�[,��$�-�mlE���|94[���I�/�2}!�$���н�m��`5S#O��p�9�h��uY�Ɩ[N�����(j��m@����%��:��:eM��`lI���+��I�N��(&���`� y?��[ǘF�V�2���NDE\���p��a���#t��F�����*�HwM)�����mot��JG P��&˼ìÛ�}��,���V�hjS[A���B����H�������UL� &̢�q���aI�$p�98'�R�똬�GG2Q�f�[�����DJ���Os��@�:�E}}xE����LKG�C�#oXʐ�2t�Zw�����Z��`�~֗�!�`@w��j�pO�t&ܭF#s��s�꣣��X����W��}S秀���wS�z�V���Q��z��@u����;�e�IC`�-w&�@�8���<O,�*y�l\]oA��>Ou��S��tS@��q׫5s��<9�ط�{�=����I�!G�Q(,��v8�\�l��l�@�R�)��A��� �����!`��@M���M�I��2��3� �i��{�]CK�
l�{V+9��Ra�r̵����!�J�('<�t�y\�K�-����>2�>v'u*�a���Cl[Z�L@�<&Q����``�e�q�VpQ]�]������~����HNV���j,��:#6o���82e�줠�KV6�8�f�,�eI�Ϛ����E����:��N�Q ��7IK��,w�p�۾=N��8�[��6�㧍�8:KiͿV%e���>����Ux��г�&�`<=�RP�A`G�6�p6J�a��5k��.��?q�7[2����X�����Vt=���t�p��Q��Y�|l��k��Q*w����DFǕm�_��!e]d��U45�[ׁ6|M����D�<Tz��Q��� �o	��.x']p�4/�`/T��gfL�7�<��J�@�r�/�/�o
�xcՀŘ�b�u�)�"#;�Û��e�x��������J��ʷ�ǩ\�[�����C��A��8O����<D�ʣw��2�gż~��2�5z�Bj�� �� ۅ�^)� �#oovW���P/26>�����f$�T��A�R���́�������~Kr������^����S����K�J�Bj.80+��Ee<����ogm31V��� ��	w�i��uQ�~�$&����1E#�6����O�Fި3���Z��W���I�}v��`f+MB��'#1�z1<ؠ;�M��R�͎�ֶg����*E�`�F��̉$=o�ן*&�:� �7�QǷ�._N|0�-sdN'@'�"��A�tE�9/!��,�j��n�a��D��
�ʥJ��Pn� �>�.X�Բ2K����Eս䊞j�ltLc��s�����Uw"S�����K]��7�������\/bd ���HH��L����>�M����s�J=�i�L|\u�솓�&�N$zŎǍ�Q�r��g8���nZ�� ��On�4��,r���Ѫ@��qV�����w
�	�>;�KH�1x�����Hؑm�%>g�c׃iz`�Ti�m���d�x���c�Dݹ�Nca	��Us�)�	����^�o�Ǽ z�� ����m�]��_w�9����h"��.	���QU�^+�s����)��4�q�'8c�&��*�}�S_�$�!�p�k"h�+�@̀k%wN]�'pk�;:[8�H���ukg�f�������#4H�x���$�)ibkE��_0�v�8
����-��F��eG�p�d���]D5����������'����/�.ҷz��ʊ7�SV���<Õm�QV�|?�2�5���^Ȇ�yIU��F'�M��v���%�o?�5z��}�`��8�؂���SԆ[
�nz�*u��^����~�o+�D��� ����5��8��B_�{ q��֑o�2	姞f��\-Ú�dV��Җ�O���4k[O!�,U���Ɛ�>)�>�S�B�p:jO3��1�*NMqXu%S�#{���dYd�#RH�ᕠ^d�Å��|�T�}?fPa8�uE`:U�Kǈ��O(x��n.�J�f��ѿ]���Z�D3��4�#k�k=�t��]��쓵g�W%q��%�G ?�c�R#�Zh����J�]ԚG�S�e�g��JY��a!�^��AܣJ��ZU�P�f����䲨�;�S���r��%�sy(!�5~6��d��-pD��ا�K��J��L����#�Ǽ
�AVt�D�=��Pq��'BP���J!}���@��=;\P���>�fʬ����v6ݎq�(�@a�q٩�ϳb݄��ൕ.x�%����2�0��0��|ԕv��&�һ�2ۯ��H�-�!���s4
���GW�S����]5vɦ���5N����r���D-XF�T�=f���#��ˆWa���W)V�l��@��D�����$���Es�K�ç��������ʬ��n�~(�����7�U��*I�9����;J:5�M7'yZQ��W�a�	����3W����G"���R|�&�h�T��.��*��X;����,N?��#RH��VE���CqU=�Dt�e��2o��1B��_��,�Q�2�}�!Y*y�͍>��D{�LS�7� _xB_;�Pyӊ&O�w]6c�\ǕP}��H	U��=��qC��ό�97����������3��+�.X�v�b��$��/9n�|e����d�0s����� ��R�S�@I��N�7���QcT!E�����4��y3��]��-s5�6� L�d�L+kX-���{��S4����0��4�]��I[o@��%|O�kJH"���iһ/���E����V����x��N�|^�
˷dU���T���O0�x���I<�U�6��9��[ᐁ�$��m�R3N�pNk'�v�`�����.�O>P3�B��DM^�����<���#�7�)j@U��K��卿�!YJ���m��/BӧK\@ �GH���֒���{��Pm h��)�+�<�VQQ[��o�GZ~�ا:b�׻c��
r�Ʌ����ӗ�J'��I:2<����=��	�C9�i瓯PH �v\[�1q��u{SS�Ʀ��!�654���-9M�	ɂ:����w�����	~	�}g��K >��mcsW�y�����w����%�.Ɛ39gb�m���Y��=����*,�!#���W����=���;��� �#�K�np�A���78��ZnZI���`�X\˶_z��}�Ǌ��h�0\���/��w���T�ל��[�X���N8";�l?����y�&�8D�y��<�P�E(`�:�`mE������O�T0�)oWr��>�C\?���=瑙��su(�ğV��K���"��\�S0�%÷ObA��|��$��`�5y|��%7*Q��hl��$X!{��ŉ4��M��U'RK�RT�S���U[g4��Y;~ȏ���e��$R�/��J�܊��D�����꒑��� �(���-�AL�������
�!�s�<سF�T�3�~n�r��%�C�/�:�_�z?��"��&�W��YV�|R��P�h�(Qg̬��rS<t�}��.Q�#;π�0_. Ob���Wd5�C`�"bI�Z���du�������{����w�o^i���xOξ�Dd�OT��,�߼[QCF�\���\�8�a��t�~� �e&%!	��E6 p[q�῟SV�N�[�����;b.(���Ћ�"(:���� m����$��p����H.E�pf���b�E�L���CD��Q��S&�� ��g�B����vu����"���hO�n?^����&J�@�yW&E���(�Х�B�1��;�_����߰y�W��
�tF�EU��l�����S.���:����������%n�^!.9jS�v~5���\S�f��Hχ�oM�z
�Z��/'O�!.	{J ;����nK��z#f��F�W�3��lx<��U��O��4�Q��}�����
z����y�&T}o��$OH��L�z-s�%���]UvNN�[��K�L�9�	
-���Ī��>�M�ť���)��������� N�p��SQ��.S�a�� Ν��Z��njǵ�`̾�gp1����nYZ�#�NH��I��T�6u���R)��@)F�b�w�:�g;{��y�"�����P�2�UF
��gP%�����/���iL�`�@���v1(Q�أu�����y������d�+}*�C��Phy�i�,���r��(_�VҰv}�m]+�������nU���.d����b��DhP3�nv�<@T���O��T���x�S8�]~rm���S�e��W>P���9�둁��i������!#�I�$��������WrW����8Є3"B�>���� o[������M_g���2<c�An���]�>̄�	���c]�NH��K�-�������*�K��8'�Hƫ����h&Ϫr��V������c�,ς�̾=40`�2��,=M懼�1��z��܋2����άC��XIa�QN��*=���_Q�u2B�2zIj ��R�m�[Rp�@.ڷ9�|�������\pcF�?@�2��R�$?=��s��C�P8L��4hc�5,nS�k���ǰ���Q֐M��a�K6������J[��1G�rQ�%�`�&��WH���(�`�������brJ{a(����'��h5V.��J<7�wL�d+��-͓�p�#��>� K/0�=d�]��4e�^ҁ�q�r�B_����n=M��
�-�b�Ń��u��;
�����51�|e�M�aTl[�KQ�N	/2�p��Q��U�2KS�!V��[V�0fg^�U&�Z<M�"n���+��s�S�r�ZG#�;<�����t�"�eH�Ԇ6�`z��`yТ]X�d8"���ߙ�@4<�,����h���kM01ȣi��}tR�8�+
��E���������h����|��I���x?��5�W�aS��DUo*]׈ �F�Q��ﾕ�Zy�X�W/0y{���p`ؘ��Su��dI�0a�ű��̝N�f(+�iȥ������8�m�qܠ Ǻ��NO/U��u	�Ɨ�$��Y�J1���7��~���}8`�=��E	���&�$]g�/�:���  �\�[�FHN�sM��ˆ7����p�&�¿=E�Mh�c�/��j���h_FMc!<t���L8I�4�cǵ��e��3�x��G5��;��FZ���o�,���MF���1:R�޴͒mSg'�@��#���+�d��즾�cr0�R���3��;I[��d�xWM� oT���.8��j�}
�oM5?�����y4��mg��c]��0p��d�;��ҋP��U�uz*���WM��G�T�q�n#�^Dt�9�'��Z5¹��3�oGW�Ŷq>|-m�IFO"	�鼍$�<�N?���t���Ա��7"���Z�gV��1'XU�5�Z�}��C�^�m����2]��I�P�6�Q,n�97�`6�S)��_��������?�}𫲡�H�V��!��tL��B�0jf�4�9�C;q;�F1�����Rڵi��2�L*>M#�N8�?���P��4[�Է��M���e3~g��s�S��24��%��-���Эc�������c�9��������ȍ�Q&%���=v tq�f����oa�<��,FG�7*%=~�@���w��2��B��E̤��Qe�`�{#�o��>�e�>�����B��պ["(_���0�tӱ��_>�D�Wjú��Y֐��=̤�$�;)0�-t�@���Z�2H�*婆K��.~������ގ��]�s�Q{�zݳ�=
frG�
�l�.�T�Pz�Mq64DIb�D]l���	�?-�E�G��8 �:4�9�qz�x�G�FN�=H7#�V�h
�{{���v�u O�.}і�Q��2-�W��#qW"��3�_J*�fw؂��*�nBY
��?����>,b�f����<N(UTg�G;;�����Ё	ۈ��Hۡ�q隺�]����q6f�Fx���ڬ�~���6������ �ݻ3H�Rxq�a*����Y`[6�"}�m"bz�A�\b_n��l��Xj����3�]xk<]��V�a�_�4Ni�ޮ8�����]�~j�_Iɹ�帛���������L �c/�;�c�Ѵ�[�S:�yN��h�_�����q�4�e�7�e<0�3W��54����T(Њŕdڟ�����O��k&��d�v������>��؆�O��,th�mō�ڲM>OԢ�}#B�\�)1�<�]4�9�.��sZ5�H��W@�%M�0ϲ�����#�ҵ���H�l�d?�]t�7���4+�����bo�1�^WX��%�3,1�@��L  d{��ws�H��	��>,yy�A��b>xK;ň�~��|]�	Yi�H+0�OM���*��ӧb��=ts�ս>;+���֍hx�6�F4t��N���� .K681xM7��v�zb��Mt�J�������|��������b$�m2r�������ΊOV���Ԫxn.P�k#�\][�W�!���@-`�Z��vetO.�Q�M;q���?�%���JZ�WB�e�m@��1�����q�����v,����_��;?ҧ�v9�k[�1��3~nc�Ŗ?|q~V�)P��g\�C3^4FxUZ�� ,�4DKu;m8�a�`f��A<X�['H�e_	�Wtӫ�,����|!cπ�Q��m�sU3�S���p;j��Y�f�Ү���lx��[puV+��%�o���Y����G���L�wb!=�k�L�Q���>@����ph'�.T�'AVb�Hv���L�P�w L�ԅ�)���6q��@	w�F�������^)2����Uҵ��k$$4��.���c"�>��Q���A��9�/����J�(l�a YH�x?J��uݢ�� ��R,�g`����|gF��6�)V��g0MO5�/����S�L��@��-�f=��̹�ݬ�y��$�ӣ�On�O�*�ZS6\5���.�r��
�����lz?�>��[�`B�W(75WL0�5p�x(�2zX�3]3�4ݲ�%�"�b�f�`9)Ikq�<��P��ܻ^x��g�:܋]���]�٢��z��Co;�%
�==`�@���P����$P��Ft�
�,�K����9e���(K��#7 � LQ��`�Ǫ�9���2��pz�������xF�B=:��sE���Զ\'I��ih׹ca]l8��HU*�4���'̜=n.���P�[yvyp;��%p�\��t��<#W�	J:�u�.����Xw�q���jB��8�$��䳀
Yx�P�S��]�	�$���|���&E�0v���?�`�F�z@�Y��K��_�@a��|R��c��&���ÙIk���e�݀��d�XԯD�Um�偶�	�i9a��r�v�^=�?^z�����\��l-׫ΰ�:��%���qj�>*�+78?�G��C�W�������$��};:�MfWtK%R9-�5$������۶F��(�s�wݖ�/S���D	7%��r\=��v�8B]V�c�캪�ѕ hy���22�	$�_X�$c�%O��ܩ9��?��LTY����Ն��G^��\����BQ���+D}�5o�O'�؆	�S���J�V&N�MС�ş��� C��|���R�7��
�˴%�u��C.�LW��??�X�.�J����