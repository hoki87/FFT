��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ���������|���sA\Ѓ�e��-��6�A�ȋx�HXA�A����~s{����P:b�� 7����Õ/F�*���f�1�fn��cWkt������
5v��Na�7��l��z�|	���/"��x[��V����μ�*��09[����Vc"�\3�#v�;��}�>d �wqv�˵W���Y��}�3�����-z��-���2�1��!&��d�3N�Ub��4UR@�2��Z�_eɮ!'��EA�I�o��%Fa�����0b���@�E�K��@�ʙ��7Qk��\7�2p�X�V��x��%�E�y��.���<X�e���ڍ}4}L߹En�#�1i�G|��܇�����'�*��}*�/@�6}91�+�Bɒ`y�C�	LDŨ�y6� �\t�q���O=���)�W���Ρ����@�罓:_fzVs~P�+B�.�[��R6(�M�@ 6�7tH]|T�opV�`ԩ��mWֽa�9-�Ș���Z/܎��~�-.~�cPE��M)�V���	��A�&�^|(C�����I�4.|��)7c�R��z�b�m#���ć�z�~tE�HȤ�u�=\w ߴ
��I=�4~��e�_�2��
sN�Ĝ��[���{*�3��2���B�7�3$\t���䧾�X�e��
r'�$T/��ի�'�cB��nY����骖�Y�������|���˩�l��FFX]{4Sh��8g�&l�%�<��Ⱥ�οb��p~'s @�*zX+���ks|B��.��������Ra��>�m��V��w�u~Ń����c'���	�o��s�W�	��%y�p�_v���+�u��� r�ǣ�����K1�W�_ir�Q95���a8�"27�G��$]����L��no�:>Ǚ�E5��[5Z5V	��l�W��X�M��E�����^7�W�2V�+� ^�F�0f�'q�269���'ObN T.Ż����X�����	ؚ����&η����Ehl
�3�c���Ð������ɕeބ�;2;:��KE܁o��\xYu�}ɲ�ll��Ö��pO�_N�:���� �A����8)��iA�W&ogɲ���c�,����<�7�.r�ϟ(~��y9/�M�w?-�;
ۂ���j�y��_h����T��+Q`�w-k�i���c�شN��q����X^챞�u�"�$5�_��1I������~̩?�3!���k��Ž�0h�4g�e�@Q�:�M�ĩ�j�G�KJʴ˕@3z�Ja/d�dkB��>��ة�~��ۖ�E��Bq�"��ђ�0B�k�MPd*��E'Ax�t���C�����6P�*n%i"�l�;YiF+��ѩ�j�D�U�/9jum�,�-&v}��?��-�Tyʙ1�r-M��l�+&�٬e�15��̟�yπח�V����Hs0 >עw{y���Tx����[����YM��V%P�ب@�1u��6>��a `}�!pB�En|