��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#�����~H�����pl�Um�v:��L��Q����;�~��?U�b����1�w���`� �2����:S���Bq��6w*��v����m��<�,E�H����,�b�M��1>k�^��&�SV%�n��b77� ��������m?��8��O�07�����v����-��Z�h�-"�f����v�Lk��em.������~A+@$���V�����z�K�Ex�;Q�2���Ij0�P~�ZR[�J�>��As6�a�!9�D0��c7�w�䔋G���ITwߦ�8k��i\˧�Ǚ��3|�İ^?��g!��
&�GCW��'W=+4�E!X�m���,0b�f"����h��D�z*�s;C�w ��j�4�������]eB�壟�������9<sc�+W#ټ��){���{~	r�T�y�٢s��`j����P��M]��H�.�����1�ҫd;����C�y3g�.E�ChvT�JE�W���xQ�(^�N��|/��ڳ�*���R'~�>1[�f�@7�!h! �j��O���6�@Z���u��8Vo����x�ֻM:�>�9T��Z�CORw��;5�\�R^� � ���{�C/�p�����xw��ʈy��C�=���8�E�{j��٠��z�H��t�Ԙ�e݊�y.V��@��vxɺ������B�Oi$��E�����,yqe4>�NP��C�Kj�/ T��9Ð%�E%0K�s���q��IݻB�!"�R�����n�}�>�4,_<
V1\���|�E�8����_��S~ū,��\�Z�/\��mWt��Ko���:��V�Kh��D�l�ͪ/����}��9�5f����w�`�E�qW���!UR�N����n���BiҸV�*��%mE1���#��.f̵([���,��Q�M�`�i�{�s�=A���}� յ�I�/�/����f���/��q/��`���(54&N'	���2���9���&�Im��X�)<���R�~��C�F&PDv=HK����٥�}��B��>����fH��Ȃ<�{�`��*dB���ղ]ε*�.�.8M����:=��a�MLC�HU�4�=���S���{�,�XgT�m�]_���l� C v�������G〤v��B���|�xt�Z��x�5�Ŧ�#e�h�HV�^����4����R=��_4��gF�	;i�7��-/T:e�g����t���93�q�|�P�j�C��	�	��ZO�I�b�sqw�'��/O���w������k���(�څ���=�e7�=7���?�d
�?WBI|$�.�M�\`zv���c)�w+pe~@���UT��I���RI�ʺ\��E��3�l0�F.v0<v|�:�B�d8���_7t��V�07��T��c/4��K�W�����dH�ν�����$�Y" �$�ْڣ�Nk�7 �����l��i��|�q�]�ٵM�Ap���=ќ�Ĕ |)C�����I�1}����J��Y��$�y�o�pv�x��Xz.>'��r���_�t���p�p��%�(�&Qg=��%��q�n<EH }}y܅V `��C�����V�Z���ٺ��*�`ǉ�}7#+��Tfeq&\���Ij3�	��@ky,�F�³hD�)ts�Sy�� �j碙�>@�?x��)����]��]�<��`D݇��5����$!Խ����qWv��f�5jb�eE#���[��58!�Gd��فK�f@b�Ywv��.����m�<���h����&~�VM��\��`
b\?�K*���PM�ZG-K�0D'w =jb�v�1�<�A�r:K�;��I�eT�mF�?(� ���d*�j��.z�n���ѢP�9��7s)#x+����1��<<rf'
ܧ�T�u�=�X'.ۥ��Vz�Q�LxO԰{�L4%x%�
#�n����o!�l�mZuv�(�lf�A�����n�	NĮ"��g]�3e�:ñ�������;����Z��ӆ��t)zW��Ty	5`���J}�n�ѵ%�	��;���~3ڠK���l�����ε�_�.I饇M�e�����0;�:f�b<B��l�����-)�f�;/ڱ�������ˆ⸟B�r�֔�z
��[�V�t�gϟWߘBq���n��̖����@��H��k�w�T;�iH��}�у=�~?��ڝ*5௝�3S|� �kxyai�,9!�,�i^hwx	����H�'r��)����Te����_MbRL�?��b<�-�m\�:�涋wɕ��D@�3L�kH�����#���Uh�8p'U���V�3�(zgJ�	�s�;�����g��阥_�	Oy(��gx}�/R�+{�%m�	dF�`3Gqm�/P�Eₘ�Yҩ��ғt�M1{[]��!\o]�\}��贞��R4���;6��w&�9�<0������J|�F��J�k'�@���r��7����� ��C��@_s��֍����N�~`���1����t܉Wǧ�p[*�[Vf��t~����Ȣ�5�ҍ�W�!���y�X`�\��|CA�£������=�sN��,�0�+���-���
�Q`ǝ��q�%Y�Bk+b~�Q�[�]�B�6���]���S����r���q��Q��'�:��ˑ)�����))��������}K\���X��9�{���N�Έ�y�L[�����ךL���G�ã�Ji�;��������JT���7M���82�&�,��m%�j����;+�����v�D�=�O�ƒ�Xw�Q�X(�⪡ϓ�-<V�r���T{�Q�ͳ��G�A�;\w��mHj���O�8�>�6�����Hn���/��`����@V91�a3^V�{�FQ����j̂�?�!V׊�:x4#���aH�5�5c�V���8=�g��5�b�z~�t��9��@��l\�<�� �d��F��=A��2b��L!�:H��H��s����$�.Z��:��=��A�n>��"p|�Ҳ� �SȅG���N/]<s����U�xMq�%HTf���C}޲㖛AX!w%6� U��+"��|X���;}`����η(�v��Cf=!�v����2����u1�19@Q�8�Y0���˝�Y�9%Ӣ�OA�=}~ǣ0�2m�Ǒ�jE����US�Ƽ���D��JkĖ�G�{��C���#/�ca�����H��/��I�axOx�C��I5`����FG�_���
�ث%|���׌pl'��* �K7��'R���6*�sՒ7������UuG�џ&Ҳ�;vZ6��![��3�җ���mĦr���?�ę��P]�̠��A|�x�QԹf'��#�T] w����{�������Ja�iLF���~~N��h��O�zy���j���; u�c�����:�I�'�Nz�ܷ��;,�˜���ࢎ��gE��:��ɴ�f���-)��m��#6�>5@E�g���,U�Xd�LB�7k�~�~��BE��]��"�M��j���@�� S�W�����`�}L�qC��~�%ݢex�u�A��{/l�=B�k8ʆ�g�]���9>>R�՝���3��M��ލ��V��=��۞�����fO
aszV���;4jd�S�����D���/1��E��$m�cH>i���Dg�d�*�[�P!�/Y:8��|'�3�x9�_���(��H����,�5 �A�螉-:�·�^��KY����kM�՝�U�?�P�z�3G���K��SoJ��� Í�D�{����L�|�JuCw���;�
ӥT��f<����'X�Ly�����y��>t�#ɅqCgŉ�լpM����YL�̔��	��oi^��/���|ϐ9MD񪿮��z�{�ܲ	�+�E��\!�AJl.�ɓa�J�,Lt��j�[zM�"`��(���^9o����O�`�+n��J�i0D�a�#���I&�Xܧ�0t��u�P�G��Sr��z��K�6����(g�S�D₠�I6:���ycϲ%��0��\&N�������{n�-�E#,���v��"\2���S6�S�1*4�p��'�ۇ��@�a73DL9��o,,���]�3);�Ro-%/���]�e�]��؄�Nz�@�]nݟPc�]y)-�F(����-�l��k������[�ҍU����g�����]��gw^�x��.#2lhd$I�n�r�� ��3�2�^��@����r�َ�#��u��WU�,�<]060�oCԊ����Q�7?� ib҆iVek.�L�6��~�MP#4��'����%��>��Ϗ���L��{,%������1H5��3��<IZ��Zr�7�P�z�8nd_COg���������(�}~�	��Q�`�>8��ٻ9)P�w� 3�
���zHOeF~\�ETP>�8�����p�["w�r�>l	ۯ �j�Qa	��$�O�ŘM�� ��t��KK_�d0�|}�9���q��9*���U�}h�_�=Xl���}1.�:.��ӱdx�}�����] u\���f��9{�&���(��~�^�l��o�7)O�.���A�;��01�{��P�	����CM�*t�D#�" 
�3��1��� `���x��\,U���X��v�"WG�d�����~��%X�(�\~��N��~��G�*E@x.���w֏z�`Ӻ�~�&b<��	�J���[����5k	��oiXJC�n�e�v�=I�/C�uĶ�p���N�x��(x,����/d��nEA,k ���e�@��3�*)�u�/��F�e�]7�ט���^��ϝ��O�̺C���ق����(HE����Rw#��Y���xU�l�eu�� �q�t�:�i�ɇ�0y�|������Q�D�.��ٕC����`��d��X���hR��v+�=#�^����|�+c�Ѝ((p1�B�X�h,�8F���������7��l����y���͇rՄ<�F>Q���;����AJf %|� ���b%��P1�q������C�ӹ���4H��Dp��(b�$_�?���]̀p���Ď���C�3>��m:���T�'��~:�߾���Z��\A����ȜsG�x \^��i��RC]a]P1_Y�ҁX���9vH��x����5�͇�׈�R�oǭ���$AM�z�������.J�b����e@�J�Y���\�:�0h�"-<��Q�pR3�~��%�,��zy�Fvչ3�9(��e��5�o���?���u��vmp�'�0��|�V7V���"+�Y4�+�ڱ+�L<Q����k9jE]Յ[M���㝃��t�$��*^��)��7:��>�޻��[L��E}{���<�z��(��\!g�:SsK�AFcK��l&:�a	!��)�qB����kǉ���@dOքd�o&ߡ�N�c���h�F��!���-j�2�Z&��3�?��!�iabd���9>���8c?3�'/�Wi����#�'7��5����N>�����Y������>�$3[e0��d����6\x.�=�G�Ɯ��Կ��%Rz���u_���ߴ��rM��[�CV�*=LF���D�a@�zAkQ��1�K��b�e�-<*�����w�ю8�:�r)�o��F1\�f�u+PR_�G���ͯ���?V�{a�;h�"���|�Z�&b�B��O�0���j]��2��y-�=8[ȶi�o3	>�I�>�$t?�k���1�ꂡ��.��<��1�y D�y���9�IoOC�s��E��ڸ��Ω[�hNpxk�7ܢ�b1�>�5P#�1�K�a�T/j5R\�� ecE����6�����ݩ+�VLAZ b�=��fQ�KcFP���U�IĴ�Rk������hR�)�t��:�a�q��x̨^f��S�0������$j��� �	���3�;҇�,�M=CH}]i<T�\��$
�ʳ�9�}���5�J}j�X*�Bٗ4�M���=cL�ҹP�U����)�h%�`��<��� N���2ʞ�E����0,c����z���#{�f�B"�5�&gq�\s�*t���h�e�Y$aT@�8�J��j:���-��^��|	���q����^���Bfx72�#J�����e@k�S�u��������@���7�ƚ��{�,�Ik�9^��ãԽW>)�� �J;���t� H� z� nڞ�>Z�2���V�9�5B�PuE	B�q5�Lቩ�	r�̈�Ϝxg�zx���,�kn�Hp�,��;B��醉���FZVݏ�~!�	�K�u�fA�-�����L�Z���(0RiB�݂$Q��'��a=WWi� �/��������#~%�Jy�N��d\G�ntjp�A��t�k2O����P��,�@Ơ8ȃZ�0"�HY��3��߾G2R"����E.$gDti�:�������TZ�� �mK�������!嵢rնn�6��E����0<dY�I�9$nĢcu��{Y�M�K|'���疿�S71E�y�K`�,v��z�JȰ�tJu��a�X!_��5[�)?��D�1|����˜���(��-�L,(;���9��|��~X����ʢS�Ht�����؂,�����aզ����i4��!�A�_}�Iz�ԟ?\W��]n��5ʍ0)5��EFb�5n쿅�OH����dbgF���F\����ȗ��{F/�.!ψ�~����G�7Pݶ�����qx�%%@����N��J��������\=�b�$��G��F��0�d����I� �2O�#p�䘒
=�m
o�N�[� A��7t8�
(�}k�0>L��miУ�'�}.�B� c��{A0!Ve�ь�-��<q:�8�tW"v"sӬ�S���H�b�����|��~/qN^x��X_��j]^��h�a�y|��?|��LW�DPb���~���ۄ���*Z��N��#��!Qe��w�2�U��BV�5�6�:�R�S�{�ψz(
�Rj�-�2�����\{���Uh�YS���`�]6�ݙ`�����3-�=yԏaD[��.��$��,��-+>�d��&]���$3bS�6"�H�t��
��_%��J�Uk�rqr��!�� 
�����c��ol���@�h�|r���̪��i�5�J�\�I�8�*�� �����ö0�_�*z36yy# FDR���8E0:���m�Nh*E�/:����W�dp�6�ev83���T�����o\����;�/���W�-�;&L.�s�吣�1��yM2,t��i����w�����$$[�^��}�+bJ�N�㢲'�F�x��\�����%"N�,4Lx�2�4��G�$���{(G�y �_�fwv��@<�{H��;'?F.y�m�h�y�ҥJ���,4���Wgqg���w�	#tX�����������vB)J,z���P~����[N����)����<�8wMI#��p���`��(wh43�P3T]��C# C��I�c%FM���ќ($1RZ�(�"����/ n)�!��i��	?������I��{<����#�T�R��vDn}S��Df �D�=!�-�f��Y�@�d��H��C$	K$�!�|���h�� h��H���Cp��_ᠽ�م�wqp ӹ�u�hwԎ�C�)Zj����iT�Q�� �k�`�t�Ө�je�Ͼ�p�e6�ת���,�gR��^��Gd� P G���,tݵ{@4���q��638�_��k�>�#JlF!����X��߲ ;���W7���D59?�j6�a'ĵa-����A�bŮ �T+�IQ ˯ذ;�?Hy��G��찈��c!�G�Ԋ�țO��9�V��7��\��B��V��i�a��f�^���O�2�q׾�e� �,�;�[�h$\�E�YN����Ƴ���S�w���M,�9�n���Wl�0߾>����_P�,,�G�y3RQ�n'cM�G��_��dHO�N�TJn���]�Id�hq�&��x{ g{�S����D��Oa��b.&ccu%���YT��r='� <��mxC���?�؅�:�>ϑ]����@Z2��̝�s^����q�<}�)*���.T֤+��$�����9��<�j6���;����t�@β�|���+#Lzw��c�@��-��eW�֘Zӌ�@��N�D���;�� _?ھ�!��&7��-iM�ՊN�F��CCT�dIA��33�ĺ�oH���g%^P4���*�֪����=u] ژ��^�)5r���ʒN��ȸ�ןe�g�|�^����a���/��0�[*���^�?[�oG�8���4V�"��P���@K̠����r��C�N�P �h���NkK��� ��lh�wq���NlI�d[�c���M���4�"S9l3 Yk҉��C] ��Wt�W���d�.f�R������:��Q,z���
 �)�����B�d�E�#��H�t>�A��&�N���J�y�2h��qB?¨�m��)2�r�y%�x!X�D��b��3���$*�^�!�I��Ts)\�K�
��]6��tZCML�%#�E"h�<$�|�::���`��#����@���.͒x?7�yLk�44M\J�;�P���E�R�qg�~S�:�HE �@7�I�<h�oB�ڈЃ�aWw��� ���z������.[��7̳���*O[Fc<F�X�4e�����f��	*��C�����C�ǧ�y�����̀��Ao��zHMG��E�K��_S�H��Zf�'�3g�˓��2�O 9�c�oNe;F����v(n�I�<Ox�t0��>��Ȳ�*��р��>!�����'����'�/!�h����M��M�E���o�ql��~ W;1_k#�w�aGv������ⳡ��B�%��YUR�j���N�]��䷁�G����,a½��$���������F+9"�� �����U�$7�3��`.F
��$�BTi"�Uۼ��NWM�LF����P��:��~mI#�#��Q�p�@�b�{(R�)V�n42%�Y]���� �d�͆��J:�h*X#�y�� +&6�����G�nο����S/�r�߯4��Q����Z�+��P��3F�g�+������ʥA���KJ@�iT�_N��#��^��R2�V����Mc�L+p���-����ûM6� ����z:`�p�"ƍpS�T�cK��»�Z����G���}<z�ѫ�&��A�`����ĴIv�d� �-��hu�/?;�K�J�Ob�:�k�7���G�28#}�����$Ъ{?����)�����{闶#K�����a,����>B�f��N���A����� gl?�1�6��C:��e��NX�e�
�8�wt��8;��(3��K���p=���!"4�!��p+Y�^����A�px�Z����3U�>��l�-p_��Å*?s�ǼĮ�&�"�j��S��V�?�i9�{�4��Z&1nI^?�~앛د�g��Y�Óg=�%���$;�Se�"=F���?���)��_t1��k �<��\���z�� ��ʍ]h<� S�_��3� |3&|����_/X�7���xr����'��?ɌF��]pe
둡��k��_�����l���,��A����o�{����iGD����fEh�@C5�p�Ȋs	s��f�X̰PD�;���a; ��"�o���X�4#}4�,��H���V�1D8ǭ�,a�K�e�-��.^�(.a!K�� -�r{���3��<�����(be�Q�w�W��1���y����N��59n�u{���A��X�w_F��Yw^�N5�� ĕ9=|�N��)��;=M��>�A/�sf*���ѡPMԞ��ȓh� ���K����NU`�Q�<)��ޤ~�x��Ipi��B��3ť���(?��&����ڀ�!7�^:��)ξ�-�:h�pΟ���?`'�N������p�Q�^�T(���sМ��řG��,�ñ�I�u
�֐��_k����J
Zy-�.��$��?�ZDD& g�!�b�D�i��b�-�bt�9��}TT��WףM�-e�=�SK*��)P�{u�T����1k'�n�Y�I_HFQ�=!�c
�s����g����P�	FI=tWhB�G�Ȉ闋K�k�_t�2⋝
�dfǘ��L�e�Vrm0���9z���n{�1$��*�a��S��1�19�5`�e�("�5e/�����a���ee*4*I�(�x�E#���z�B��'���$m�w��U�Sj	�q7[�����%�ܵy�b��?mt<f ��p��j>�a��	��"q�׿��f]-��!~���U�IM��@��\47�D(�nF@7��w�h���տYW�D�[��j;nHe�	�'|XV6Xa�fm��\HZ*^��U	
�] �k��dށ��d8#{.zI�f�G��dG��ЍQ���&���i`���1^�vb)���X��h��Ҭ�X �Iq�Q���v�Z �/vYg��v���>���Ebl�R���Z���菉G�6� f��`}��:�6�$�[yM���3�[��q����BJ!=6����(+�����TKlZ�[@]Ҳ�Y|u���m��G���XSR+��gyy�s�x�"-���$"�G�]�����	[�� /�f�Ǡ�!��6;Ʈc+qʹg��Z����8V)�(�r5�?�_�z�	�%T�C����NJ�˦�4j����C S�{Xw��8M}R8��Ȟh2z@}G2�9��$���S�x_�m����z,!�A�>�r�a�.��!7��j�<w0�j��Gj,��F�lF�w�QS�3I(%D&�ųZ��x@�!!Mz&��o��Z�ș������L��, 2��5	�A�j�:=������Ym���tl	G����hp�($0	��d�H�H�SV'������Y�l0-���� ų�f���8�h�q�\�8^"7���I���s��-|VG ������8�-젍(uqW s|B¶�V�`ql�n*[dZLK��[�d�L�\��-�:�����R��h���- +\�+�f:Wz�~�%<Pp���;e�����O+�Y��6���@$D�; x:� ����.���*�bԨ8l:=w�m�s� ��nä��(P��G4��s���_�1P͆��y��/��%���ӻk�ה�T��1��)^l���D���EJ�<�ῼ�+�o��b} ,���frY�޼ �������ٍ$���y�ĕ�W��ܾV��s�z�:���va��y�L+�v-�SI�:�*�@����O$?RAa��&Q�W�BQ�	�Z	��S$wҰ�ًP���!����|k������a�7�n+�%�&�U<�V�m�}6:�u���9F��ϊ5 ʹ<hW�������ՊL�@��sv�"IX ���U�2f��&�'���;�K�}��z� 0���G�c����oĖȲ�ŕm��1�;- q6V���k��r��s�|5�,�
?��j�k8?�ܭ�Hd�`0i3!���	{͔�7��v��he6�N�֌�����a�ڗ�BDֆ+<�D�dj���v��̤� TpctL��	�s"��K��h��ʹ��_��9�r6I˱{� �rt;�B�%p t{����`�ޛ��7�qr�~��r$5��M��_xg2��7�-rQf�g4����;*���/�;��	��㪖Q��:~
��"��R?���K��S�S�3A	[�3d�͋ׄww`����,ϰ�f���u1�gj���y���JE�Q_O00�[�h�n8J�3fX����F�'��7CҎ���&C�6f{B,N����`O�c�	���ꓟ�U'L=����sE�����0�vtS�G�$���O�%�I��
�SLC3L����j�e�G�����`JFl�������f9^�6����Du������N�j0�l�� ���hk�P,^�r���j-�a,�E<Jo�n2~�vU�n����i����;�X>H�t�9�}٬dVK'S�8pssqΓ�!�܂�B,i>��aK�!�Aq��.��9���#�`�/���a�P)�,��C.�>����=�)�Jq{�T��m�.�E�qGU��Kؔg��;��N�(�P3���;�!�$&�^��)t$�S� nZ��DX��0���=�Մ�N�����=NC�`^��K�����%+Y){��l��x�����Q={�t�(v�$b=<�	E��ɴ��kL����f��_�߭e#���!�Oz�GBai�d9sߛ����:�p���p��F�֠a�
�j-�q~�A�+eƱT���=�Tַ �wU:��_�2v-���O�4�� ��~
Z�����1�D	3� x$Gx�<���'�a��9�6h�r@�U���XvZ\I�-�f-I�a0J cg����n��H��Ũ��V�<DW�|�3Y�:�̀�G�58A=�d��$�a��H�4��!�M��-��+���M��-�?�?[����Q�;#SB^�(j�B,Ѯ7y��=0�7q\�&�ɓ%h���/���{%��-͒l�����H�
�X��L��+����~��^ �b�`�h�o�q^���n!����cj@s��SD\ޡU�A w��
�(�T��x�4p�<�X�g�ȏ� �9���
�kؙ������Ȥ~�A���8�b	w�R����{�<��e(l�ʭ|���Dl�߾?�H�l���ڐ{�L������H#�G'�@��li��ߝ��g�!q��g?�U�xDF�q��D�1����]�HT� s�a���xh[G{�ȭ/�t�����hn#��/X�CL��]�
�H�XC�C՟����y��Χ�q����O�w#h��z�ޘ���Ϣ�G�(onk͇A�v u���^94��Ͳ�,�
�wd_]�Z2��&����f��_�-�8�I�������n��Q뭔��c���Ub�,�by}4P����y�Ppa�鄝�m�V�X�a�	�Y`
"C⫻V*yߟ¹��na�hD�C���!�r���P������#yS�؇�˹���4ނ\y:&=��C8�J�˹�:�%���mPT�*uM.D���F�F[��+ �YSS���Aݢ-��Q�ֵ`C�ұo����B-A�w��a�������|�*���Ǫ�+�Uڑ�/��d�I\~AJ~��נVb���r���w؝�5��Kn-=�%�%�}�b��=Z�m$��90�
������ˌ������<ꆞza����(:���v�q��lT믳��@B#�1eu%q�N>�sD>�vRYA4q,��8`�7��1�Ee�@��y'�Y�9���Q ��j�C�}o�����6� ����p4��<$�̚T�9Qkp�����b$�3f*
L_�K��������a`���2*��Ơ�y"䅆?C���n�!���]}z�������V#fl�H����D|y���n��4�3p�ե��P�[ʌ�i�sߓN8��H��l�(ء���1�y-��ia�eҬ;�+�wpI��t�*p�~���.�e
��Sv��W�S� �����`<�g�oŸzm��4&����K��o�!��Q���b�^��͠�U�����F%�-�_��u�죻۸�@���h��,OT��V��i��|v����Eb�c	*���	L:�Nލ�m�� {���r�y����K�������)��Բm�<R�#	+�l��M�C%���'�(�uU�PE�b��1b��)��yR�j��o8�w}�+}8�G�U!,�b3)D�U��v���,>5�Ax�P��`a�����}�n��K��3��Њ;2k�L�k	^N]��O�"���r͓|�%B��)$�#0��j��C��7J�S�:�ǦSK�na���Q���	54ܛc�{�Hbj�)e�	���8�]jkB�����R�wLg�r��Ĝ\�h����>�#�K��żwTR�<�c|��2�-�S+Ѿ�<�X[�7t����?����;��p���!lE���^j�<���C�֧a�̙�@����b]5����醳p��=m�#��O��;�K+IK!c�r k������)����w1�P���z��⌎O����bs,`�1����P%�\��� ���&a� M̋T�@K�m��r��q�K���C��4H1gD
���˕Wh������o�$�bt3O�F`c�Ь��d��k���+p?=���4�\��ga�<Foi"���>�ҝGτ�����n��(J�0��T�r|���x�?�h�����f~�̎���@���\�(^�Λ�D����W�G�7� �?����)���Zz�����^C�4J���/G���9�bdz�ӰQ؝�)Ks�6j*����6QS��k&��XR�Wf��o� �o9TC�%%�?���;�/�%�a��`�e��E���-��Y?�ؐL��e��|�*Ʉ�> ���{Ko�ZP�˺cw�ahɌ���G9i�/���vP���9��<yi5d+�h�Q/����N�ը��=�>Y�v{�r�,b�0��j���,	.αV�7HN�b�4H�2f9��� ��\@�*h�S}� ��O0�Hv	�a��P{�&���P}3A�m�<?q�D|���x���F�?]�^M�ڑ��
·1�8�P^�����s�m+�*���v�x�%��b�=Lh�,:��X������O��[�ၵ�|o5Ƭ!I�vk#v3$������Qe�_���
d�ʎR������}$�#�:�V�+y�S}�tc�a���fk��z��>����j�L�NfAFA�IϓV����H�~S� w���I��daB��Ͽ���!��f��/�:5�Ŵo,9�tέy�K1|	J9��x�����r���B�MJ��E���<���T�Zu�K���,Tő�j�g3Q��,�Q+G^T������!�Rta�e8EA9G�Y{U�F��à�g���e'�OO��|i�{8��@��o"�o5��huWZn���S��"�J5���xX��ڤ�>+Kn�I��LY�ש<�v��}n�{�5��k�A%��H�F!5�)
��y;g�/�(� �7j�M{c}A-J��}�WL�֌����V�عH>���6nTJ�:Q�]O�lh.6�䙄�� �[QjKB�%��cyD(��L����q�	~:�qW]8�B�����f��U�WwL�E�}�|�t�r?���aij"n���[YF��.5�K���ф��R����/�eHo����p%%��?Bi��ފ�Oz�X$ķL�F[� 	��r��<h�χ朎*6kN��ط�|�#��%��E*u
�
䁺-��cGO�R2�(��c1�DO��e���n�J�0ܓ�.��9��ߢ^��i�t�E LЮЮ"��9HN�S�Q��Ǎ�4�0o��kt������u�.|��-�7N���(�b݄N0�� ��Q_ӗ��i�@[#���6�h�_�r�k�A��2�)������u���F�uL�ғ�KΗI�aU�]!+`MU�x�� lG�xh�H��=�sĭ�(��,A;�,/��:S��n�"|i�[(^(����ׄ||�~+��4j�)i�4�ZD���c�"\؏Gd���h����U9��� �tcW �IV�e�b��:y}<)��ͮ�i���s��o(r,s"s*\����2��O�|�dcs|8�W�_�;1W)&��5��f��A
K�Ape��h,tw�H�E䋛�oq+�7��(|�5�bW���Zh��.���R�M����)��x�����zL���D��j����6ٸ�
�w�63�.�o3-}ﳗ}�:�1b�nD�����P��o���H<��SB��Vx}�$��R/r���t�I���C���,{�O�L���	�>�j E�љ$M���b�P��;S5����>6�씒Bub��M�,u{.
�i!DX�?!�ȃ�]�/}�g�=�Y"�'$Qɩ���� �Q�Ǝ&pT����ۮ�KT�D��j#���Q
��O�9�L6�3�W���9��Az�猞�@� O�#B�;�O��N�{�2|t2l ��.1�oo9X=l��:���	�j79�9���t2W���d���tK�g��;����v�f��݃���u��FA��$nĪ,�T.8['�����\a7�a�m���c�J�i_s�lc�		�����3���1�bTA�7��N�fo�|�� ?�Qt�� T�=ǌ�"s5S@��޷�������]x}�~DS�ږ���2��sl�c�{�=����|J�c}9�R�/r#�K+�\z���|5��T'�E$
�<qg#��m�eV�M� e��E�7�BJnA�#����֌�cC�a��%*P�q���n�l�VTl:2��]~m-8�5��}���E�؀����a�3�BlQq8�(�b~��V{��<-z&�z�p�U�qJK�M��X��g�r>v*2Yە������XC����No�YM͗�~jy�
�<g��B��_V�`/Vpa7Ƅ�jQX�HH���-���A�{M �����${��@I�-z�����*�K��[���T�Y0� �;��OG���-A;��;RI����d׹�Y��"��{�LR#��%�ø��kԀt�D	����)�xъ˯����u���a{w�n;��p�����bH#�S�y������oӀ���>�]� �έL��� SV�z�yd@IWp7�8[�D���Z%K��g%R���Dn���/g�V���,{�M"�NM_�ܲ�H�R��5&�v��Z@1D�U��R�g���{���_3��7�U��DC`����e��fj^��)55_�S��2�.�5��q���m�������������:��$�`�?-^�]o��d0*�shRT�`����=��P��Y�ѡ�ZUJ����G*-��K%�Z_�y�샯��.E�����}�>��4�NCX��~��r���.��1�|V|�Ym�&�Ɂ��岻m�ʶ;������^���8+%�b%z�c����|n���@��ʻ����I�P��c�KM㝏���+�w�N���6P6��T ����S��?��Z��NŰ�PiX��V��u�
�����D���~�U)`j����Pǵ�>c,k"������u�}��
����f,�Ң(,!���).�S��J�ppօ�6��u�)	U��n���x�V}g\�|	�g(���q��&�H�<�-��n�����j���ں��(r�`���*��p��}e.㧙��|�:��c���NR��"8�u������;���x�E�0,��$朹>Ui2>�5nx*$���s�X{E��}�:��ڗi*��"I}V[�{me�)=.$�]����"q�wh�J�m:&4��d��0']��*81��}�&�Z�F����8a��������~;[>^w�,8�7�msr�şt��O�d�8	)<�pjQA(�/�_.��)�ڹ-�,\�!��Ҵ����_�`�z�3T�f+���$� �PZ�JĘ������]��Y������V����
�����`hN?�sڷ�]�.���%�X�͚�cz�t�陗Nv�l�&�R��ҵ9=<]*b����f�C*�
��jy:+t團E��+®�4_� L�+� ռŁnYQ��i��G!k��Ӷ�q�a�)e���(󞍅�X�. �ԘN���MaL�T��mޫ��+u܏�3H��K]�yqR�Ͱ�n(Y��׬�`�:��>��G�52���F�I�i��e�T��+���v�vMآ���w^+�D���>��ڕ��,���Ln�n�Y�4�aƸ�g6IۖQY	�����=�3u,������<��~�ݭ���G�tb��?�~�+�i�%\dOji�!5�����?�GS�^�>����y� U���<�$e���LP������Y�n@S���*.���u��̺��������Q��p�3V���XnP�A��D?}�
D���UVbH��;Aj�2�"�툝�E�E�c��a펌)UĎFڡ�	�	�k��~ǅ�_�hX�&ʫ�]�@Fy�%=�����yXCa(:V�c&����en|}聇Qdk��v�8Jr1��Ȭ]VҾch��x0M��En(�(<�9�ȵx���4�ͅ�3F�����.��x�I���xb��7��(y��cY����p�@�/[l~Z�)�s�w�:捡vm7�c��7kqq*�S�0�}I[J+Tp�8HG��Dv2�&�g��V��F��q�Gؿ>,w��W������-���S-��b������cV���T-���w��f���i�=�i2��j05*�J���B�2}9do=���U`$8�j��T�2�k��t鳣}�o�x�^�N0������{͕��4��q�rD��_��ӛo�q?�1j��������p�Ҷ���0��'�޳ �r�x�VOc�$���� �ҷ����9�,ۖW�/x2(��O/|�ӆ�~��]��-�լm\m��\,�E~XvrDK �i�����(;L��6@G*t�1�� ���t�`�S�����:>�yX�ޑx�5Z.�BPq�Q�u����^��@$��I��2m2�X/�(x�#�9�ֲ0Ф;�[��Id}!�Y��>�����i��P���$#�����_]�����˧�+�@�0�����R�KTm�hu��Vߠ�?�r0�3,X�i0LF&-��'�������)����){�#���P��T�S.,���U�F�r:��6�����_ ~�����DZb�\%>P�]�H��r�4�]ޕ���/���K燥�� u�-���Ӫ��T+�Z��{�8��E=��fV�C� ����ڋ��0v���� 63�6z�=̧�ƌ-92�:�ɵ����<�UU-�(�Z�]�� �$�v��\�5s4 �� �a}�g�ƶPֲ?&�D
�g��$���87p$�w�KPJ����\��:�
��䣲�f���ɵ\�wc�D��=G���o�rC����\#��fx�O�e��^�.@L�.c�@]־�#J'G
��?Nn|+&��-Do:�4K�_� 981Qmw��z"�R;����1$�%����x���h��S��3R��N�re�r��q�ZCn��K��q��
�������_T �^Țy7��+m��zx)����|��ESmIns�%���D@�ղ[:�;�\ĺ���>�
���5��w,��=$ǏZ����*.�M�մ�dμ�� �o��מ�P�#�a̑�@V�1��S��F�w"FY�e|��z"��XS��
�ͮ����VT�T�ڻ5�;\�KYl�b���Ȍ43dm�ϫT��x�Yn��t1����y�-	��Sc֟�fvZ�LQɜGg���X���?t$�[�8�ϙ�rw�z�:�e��ษ"�����ڬ�d�Z�R���\����������uRdfަ!u�R���3);|�^8ř��2|�=Ν�e�<�*:�W͚�hv�R>��9 E��Թ�=>V�~��OmH�&�m��uW�%t�>E'��sִ�JhZ�Mr��^���n�~��ђ�hb�"�>7�^�r`���R�.��8Ӆ�i<��&a��8Ӷ[%:4y���ᯡ	Z��#�߻��u���BV2�B5+\�u~1�P�]���1X�R�H�i3[�>�pL?�S���^M/1p�P�8�_`2/�N�D����T4�����;�p�0��:�$x�\A���,A8I;��� ��Rq��1/LHR��]$���$C�Ϊi�-
�u#liզ�z���_V�r+���0����T&"y&����b/ ?��𑺠y��Oȱ��.��z����m��~u��q��"t�'��r���Uܩ�G#N�=��v�_���(�RqxmH��V�P�
�V���#ܒ�5������@c�@?�1�`�� liyap��~i��Ԕ0�7�3�#�?u��vG{�^T�y�v�T�}��	�uXl��G�ɬ�U��n��]AU����4Q�v�������b~|-̗��9��G����m�����򕦚^���e�a=^��0�l�@��1"|^R��j���J�4G&3E��$8������ư�9�*8��R:���ĊIk ��,�g'�?��{6�<pr E�O o88�"��n2�8�QzԒT�܏��Nվ�ܴ����ۡ��0��j+R$�'8x�Ӧi�b��0�T�7Z`�Z��k"@�H���� ��b�� � ����[�sj9���Gr�$xx@[U��_�|�@�A�{9�����r6ٻ*�8���r�A(�ց���kU���ʨ'Du*=�}�Sq���Q��WS^�t��05��1�	RKEa��w�+��mZ���v�\�pQ!a���VrL��6�D�K�ʆ£)s�#z����W��$7N爎����1��B��\���(y���+�=%���I5��\�#L�xE��z�4���"s�&tx�"U�c-���>堼�s����2��a^��NԘ���C��c���&��o9Sc���юc��i��1(k�a��>�
��C�H|*c n9E��s���/+#G?��^�o��(L�	�%�{*�t�\U,��?.��7jCr5u����'��s����ɾ!�M����;?a��&�

��@�O���'�+�ع���`��N�O(,���A{+�@W��d�{��"i`�p[�s?�p��Q=�sqT6b�NU���g?�����"�}��c�:rF��s��>;M3�Q�$��	OP$�w��3�]T9ؑqͅ.�'��ޖ`1�o٢�|��&~�H������z���=:�N��<�.Nd;��5�=�|lxq{������.�OP�Xgr��27���Bq��2���!�R�
�a�X��g/��N�Np�7L�Z��9�.��b���ꙿWǩ<���rq��_�5+�ΩB�\�P��SW��_�)�lĆ^CA��vfV*}~6KY��
�(ѝ�t-�% �>*�z9��1cSe��"�ږ�^�����`�-!�`�!o>�)z�Z^^�<d��A=��*N�Gt"��)�V;<[�Vb2�b��E+����*I6>�	H�X���a
_Ȃכm&�O`����>T_n/+K���TXv���"�h�ٍ�n���˪�Ts�=���W�K3&~z��3�S�?�+Ġ���#��lKpۧR�O�i�Ƌ5�:��j�{�}j�������s�}�F	�d��_I��枚��C���#�,��FCS�eJE8��kЖ�4%����֐WI�oR�n�-Sv5K��Ov;� �R�Dj� 9��RZIG����q�JB8�p��;�2B~nCE���F�*T&�,������;S�1�:b3=����M�v͙��ݖ��3;�30�Ddl�Ϡ�O}�R����2=�W>B�'�!N���Р�U���S�V�2���/kO����?Ďm��(���22��~���w��K)>��G��y�A�����j@h�^%����d>bG����M�v&A����;��b�zw��K?��vX[~�p�����ʟΈ�Tclm4�o?ycGűvK����<�%���:�ķb��1�IY�rf(f��Y;�o��"ZR��f�5�u�.t�b�����9�W[��t��x����A��&�-�U@���J�m��n���L��r���7����5���t�$Ӄ�o�j��r4��Zf�(W���`ǒx��[���u}�,fs��(�g봝�I�l-Q\����I n���C��IM_�t%�6�<3!�q�X�.����7k�Yd���9B�ہG���I,#`:rm%Y0����O{��:�~��	ł-�3�Ҝ�]���nA���������
t2�$9���sVR`I���d$� ���Z�`	f��K�6W����D�V+�����@Qǰ��d׮�b�-�)�V\sB%�V���M�Y绖�N�<�X��x�1,(���);�Z�Cǋ��;�o��{�=��h?u�z����]���9	� ��g(I�4R��>�v#9s֨1�m5ڡ���|�C�*�~��_,���}C����O]l&zj������P�̋L+
���N�"T������kۦB�*sc�9'���#U��/�>C�!�u1�`��JX@���|��������.�%���O�(!e��\��A/�7�[O��(�����h�>2(<���T�_��X��M'0kP�B��v�ʋY_r��'� fϷ���4@��7��&�,�dr���6���$.[�$�.�i�ޗ/6�v!�.H��.�������7!$�K����q��vd�;�bG�"��{*]_5%�jfm1DWf���9��Y4���+�4��j�N�>^���&q��ڄ��˦���l�!t�k51i߉~;sM�1ݨ� ��Se�mep��x�X��XV�B�m��9�w���h�d�UT@�dO,����,*��kzl4]�J�3|`�~cWw�P;K�[��w��;Q���&�$"����j9�9�����h]A�S�2?�������E�:�E-L)��?�fc/	T�d� Ÿ#�ufcn��8��+k9�b����0�������o΍U�e�h�{���h��#�?c'�E{���n�Γ��
9ׁ5�1����YŴ3���L�ςG�R�Z�����m�4i*���b�����"t ��w�aJ����;�B�}�
P��ߑ:4* �jw� ˓�F�'��1�d|���XN���H/D��bvX.���U�����Rް,���(���6X��C[�<�W��t�GI��3��af��=�뇚��j�(��ޅTL��r�2mX�F3��Z�)���u;ĚuY\���x���h}~t���4*�׳"�^�ڻ��tV
&�Q����Vu���F�Ĵ�� �뒙��e���@3A��	�	�wY�t�-Tuܜ�E���1U�)�\O1�F�jA(��c
7�ȣ|�Jl;�ߕ�E*-��[��/:޳�����f���-D�
�;@���p��j��� ��4�
b0v�>7�j�ҫ��?�wt����}�	��B�G,I��P���2�A����N�(l`��}�a����Ͳ[5'����֩��w��de|b���'����ke	�ʫ��W@EIc�nŉ���t��/��U�mC�����?������Ԭe>��-���ܳ�L���M�>�b[�o��[�a��|W�-ߊ�4b��6i޼?��x7�kY��)G��\&1/�������`<_�B��`ة���B%� �ޕ�I�^��5��/��1]IX�t�O���NDB�.���N���GV����۰d-6�7ϑ��i�����lc ;e�}����F�a�#��{�����uHp���� ͞_h�,�!'5
Bp%hq�Ƿ"9!�j��%�B��twOq}�9���W8���9~\g]��A)��yR�=�DV9༺�C�m��6���Yn�Rou�O9��MxK�7��soVn	Z���g���{��S���K*k욏4t�N�9���4#@��g�x�\uN����w}�b�hOCi��(��Z��%X�`��f	$��yZ���H�yx,I�?�
$���۞:��I?A�{k��K.-����sy�U��_�btp�� f/�n�b
[�Ћ��K1�^?�rENbN[ip�Lŷ� |W���#}�=a	8�6������"���ٽ�Z0M�Q��ϻ���2��Q�̯��-��k�@��Z{ J>N�	d�jF�tx8��;�dLށ�h�_�M`�G��Sc�6[$)�p�{r��)e#5��W�����`�?���bYX��T1D���p�<���6�X4�zHxH��Y<m��L�Pop�U��Zɴ2��i�,�Ĉ��fcW�iSZ�3+��
�:.��^��>��4I�i�N���>w˷~��Y����ߏ���Nb�zC�9r0�z.�k`�����!����2Ǭd��V<�X�##�8������֦;fR�C����ѱ�!�t{Df���rqYf��~zۓ��s�!����ớxռ��K+\��)���:5�N�!2��]��{nװ��y�ȉ69������0ǡ�V>�@�N���l|V��Mf�����:@�y�EU��1598�z׋������Q{�s!���>k�~Y���
�h x��o������/΃3B7�$1�B�Ju�eNq�5C7W�4'��P�U�%����;ev3Gt7��/� ��iu��˂��FY�.��'�����{��ʗ'��م�۷DzU`;:��h��F�JF� �WDk����@DA�x��^�����zbz,G�	ǩi(�v1���+܉��ϭQ�M�Ba�{�ޒ&�M6L�h5bU�"�ZJ��u1hc�����|�4,�\���mF�\���!�%T�����ݵPS*~Vn�
�V�A�����A�R��k��P��sz���t�)�f��)=*I��,,��?\�� �E��SB���������\O.6v�lM�9k7��{׸Ji�4�η6�{~�������D����)���a��]���S����p���S1l�L�P/��`�}�K������Y��k��2��Ii��ٰ�v]B�,�	Y�$�_�t�RwA���P�=���6w~��0�q��i/��N���	r��=?pC�kM�* 
 ��W�BлT��X�?�`ׅ� N�J�� :�.=p���@L��ۮ枏�`�Y"@8Ń�L�D=�����y�?R�D����5�Jjv�3!���O6��y}}�yL�38ɀ��$q�"2��Z�T��{�����mvgۻe�-�
�H�~����5���@D�s�����V��sz�q�S�\[o�k���I�M�4�ز��O��	ߜ�
�ؼC�{�sd��}��R�"�t�n=_ͦ#{I3!c�\~��k�rM�` �������rBV���).�?�5⻮��W�:f�F�W�3���3��RT�_��m�Fj�uc��8N�v���7;}�?����fv��o�
�	G�7�_�Q�I�j�=�k��]7�z罒HW�1���5�4N�n�9H�1H:=w���[cs/�'3s L�pj�3\�Qwz��a�$�u��?�q\'�_N��׉��[{����^1�H���s��&�Rz�	6 ���4���#�m3�:�jri������ϔ\���̟*�}��rv+�j�u^�}�9*KX�DQ���DH�oS�Ĕ����1q8���)h�kh���f�\������s���gvIe&1#���a����bu�[ ����zQ�w~i���Ut�Z�8S�O�ŤBr��E�Ϻ���/D��݋醕�|5�Hr���ڗ���X�0��U���Od�N��d=�XFQ���ţ�}�+hͬ�`
�����`��H=�u�����:wkB%�Dg��o[[����g�?2T���(p�:%!����?ƙZ���0i�%BTF˄����,�I$.�X��#��Kz��+?�w�hs��zO�R��Z}>� M�B��$לq��t^�����:��srf����Y�a7�j��)�Ab��&@��q�0#
�ԇ��E��)���AX�e�[�1�T0�)("%��:�0��f�� �Bp� E�d
_�Πb�cQSr���������XX��ӹ����mT}beh�����QY�Z��2�m�h"���;AL� �"�e	��k���O���x����">;u�H���:˙�"̇�3��a%b�#�^.;a&��U�v�;Zjp����38ڠ�1����;�]�6�d|�3���_b�w�c\��Sf�T������E��g�Ěy��.�(���<`(�}'|3`�8�x�ܸ���zҥ�v�=m�?k���:0���#�1/���2��0�b�?[�\,ϠQZ��-�<��V%Q�i,3���B�.w�	�sP���O���֡��n8-/c�B_�H�� �]0���xAp���ʯEE^��g��+�ѱFF�+_k�j�$ciPbC�j�r?#�o���\M����Ů��?_�BR
��p�6�5A��e]lɆ&��e��N����2(�������j��|�l��^�k��fݩK�YT�����B��	¬hc�Da��e�%!��q����?J|�� hW��ۢ��Fw�ȵ�����ZYX�g(V�T�q�/{F �nWx��wo�R��b.q��ם��������y�c�y�CO�_ ����a�r8_"�9�s�
�o�5�����7�hp��8������L"|?�4\-䉣K׿�Z5�� ����<�
�I�W}4�v7����.�,�W�ЇڷV��F�衽�9	�7?�ya��")0S\��a��X{T#�ef�@.�'�7"� ��I�l1��k��)V����3���Z�'??]䦱�{Bióp���TFi���>�>�9�f����s�K�QSG�6�7-�-G���M"sL���ȫ\gο㹢\葽�j�&�)��蛱�z�ӧ]%;y3�_g��}�0���m���.��F�	Q<�dFy���'}f�N4�U���^>��k����i����0������z<
m���_��5�|y�������[�k�/�����j�U����˞?s��Ѣ�{�/��oz)����ʛ:s�!��F�i����*���y�
�S��!p5Sj���eE&�k)y�R�B�:��{g�Uj����A�� �0�&�fo�@�m�*�x�a���8�����hU��j��.����Uٺ���>3���0���:G9�-U҅�p��I1Ͷ�����W變��4�q]a]V'j�;\��}O���s�7���f�D�1��VB�������,�ԏ|�}h,%Bg���L�o�OwY�i���y+�_�F� !c�G?����.3ށ��^��9i�[-}*��+��ɶ��<�Ds����vZ�?��b���ߨj�ǩO����HF�A2�����h���;�/�8��q��FYAR#�֊��Q�6Ov��l�ͦk|Q���.p�_|Y��;�]�KYh^R2���N��	{+�^Q&�2V��T�\S$C%ȇ6m�h�Ϛ��C��q�����<��ꌯ�1MTND��!N�W7���hG������g���&"©{hD�i0�#+�kD1����٩͗��Q�{�Mh |˿�Ke�i+�T�տ��P�]�T�_�?���Xeox���Mcn�$^u�����$��ъ�)��K=ߵ]��f0�Q3��t,���X�����hm�h�C�Y����D�)g"��\7Ib$;,�%N1���[�M���A���:+dc�HϚ��J�,�%��bH�QG�y
� ̝��7��;�H%�!Q	��p�l��J��o�?�O(ÄzP Xګk�k�;��p�S�!�c���fcugq�gT*�siv^=��[ ��v��	y�Kn���{^�`�xW"�yr�wbF���u:�8)�z��L�Fb`�V���mI�����G����h*,����n��`9`6K)b�V�Iw���+����TQ�>1ѻE��E.�U�?���xWE����n2�����tQf�to>��e���X�l����"L��dȠ�S~��������$K`��߫��Mq)ցI�n��H���'���]���&#�|!/�֒��e�. z{�z�2���9v�W��@۾��c%O�+T����G�O����{��x ӕ�T��M������\#��I���׸-�%���J��vؓ韧͚Ƃ���i�*6��=��)����m[��/�Ht���*Ea�X<�nK�=�rI��!6e4Ho����6Ce�f��X�T4���d��E2���	.�>H���L]�lr��o(��$�ەf{�zT��ӯ�j�-����B]����9O�.}h���Dd��.��i"M?�=����^y�܏��{M��qp�}T~��0�����+lDX-���c��%�*G>�:|������a�x��h�aG|�_V4σ}=�i���mZ����9��)��M�b����W���{����������#б�j����Z|�'Z.���EH�Ú��[H���҂�?AT�q�`�-З�?���ik�O�^��V"���"1W/��/�2/���[/<�-�+2?����r[�I��Q���R##�_��A�٤����<�����D?�W�T�����[�����i��H$&��]uR��q�H�ַӊ"y�$������k�4 W,�B�8�I������v}M!��uGpV`�0� ���&<Q"�QR�&Ƕ�c����R
��;�qw����cNI����Ͷ
]�c��{��
���h�>�$n��.���2����rA�Y1�v\��d��)��wXa�m��4�u[�Zf�\���D��Q�g�������ʱg	�;	P���	�G Y���dص�Iƨ�m+�_�v����C��R|#}x,gG�P��2��摧?�`l��pX\������<%��r����b�?��֦Pv^�n]���霏ȚhT0�>z�̪V�W{,ikA�$>�?8�U� �+ �(��"�1�@\7�Q�D�\r8ۡ=��x���#0
R^�%�>7����͝Ӈ����zy���&�kg:C^9gEvS#;D�\���5��;���)W�Z zs�R���[�5���n�k]w@�?.���H�m�xF<?�q�|��{���myb)z*��.����nJ�@���3\�)\V"~Lc��a��_���(���YΎ�LfN�
�%�a:�bEm	�+18ԉ_8#E@(,�V�*�*����-KM:�Q����_7F�EɃD�-
�xt<�]��-��Y!��e�1_s��錬,�!�}�z0.��:�Q�����- �35t���8��)a-��@Û��÷�M~W���t���""PD�����/e�	4}�\�/-���Ț\��̃�k�,f��_�?[;ժ*z3��T�Qt��RN�
�RQQ-Do��)�? z�))���C�*�A��ٻn�:�v��S������U���o#/��~ �������R��7Kjlwx2@ߥ��|��XM�����K���uXڕ+xp�Ba�g �5�J�{Rִc��nF5(!p��J9�?J۷+����<^�&�2e�r�=F�n5�:�N�>㸈����&�vO��i�ұM#S�drX��2U�1m6z	���
�g6	�kO�>S�=�þJ�VH�}�_�+%�z�6�4U�5��M!�`#�����ڢÄۛ��qo�fܙ�`��=;�<O��!O�R+Rsي�"9��Dt��D�w���Yd5Y�auzY0�4���-���iR+�$��J���'�������m�_�:���R�s���!v萴l�8C��qؘ�5�nB����j��w+�/����L�J�������{�&'�qŏ��3��G9��0���\�һdT�^�pɧ�P8�~D�c^``ɀ���E�fo(l�B5�V�v���O-���ב�պ����gF��nX���-�t�e,F��1�1c�[;zG�J��i��l3� %�'����Z�V�\�DF���so���p#�s�3�y��?�\vf���;aAˎ��K�a��kߌ*9�Ld����13L�*P�!$���j{>v��/�������m����+϶�a{�,ѥ�IX�R��/:�0� v�*��-8����5#�\��D�A�ˁ�^�r��gBF�G=��0<_�*PO�����X5k|m����"��h@��q/�Qvau�����[�&2�˱�]U,�?c$�Sc�Wh����9�R�����v�P�.�7Ԅ���_hTo/}�A�m�X��2�&�"�x���*�À��>M���VѴ�͕b%��$a�(P~�A����A�E&B[�~ɟ�ڳ��,\s�)���y�OT{AM�&�4&R��E�#s��עvФ���� ��1�%�>`!���ݰ�5�,���I��/�lV6��(D�a�����;�K��@��'�S���(V	��{���,�9Z(�M1����E˙��|��ɬ��c�^��:p,e�-oU$��u�Qx���4H�9,�2j�S���^�͜
!~a
-�T.��k������q��DAa� ��b+�"?����)��3�߰4���g�7X��>����3��UC��L��KJ[����M����Ѧ��5��Eh�O����8����u8��ĘQ-�k���z��Qi�5�Lx�͊���y�M<pԠ�f9>kp������c����� �a��>u�P���g�zU"�(�~֊��vRP�Y^�ߦ�0X�f׾mzA�K�.	'VS�+�}��!�	��l���Ta�c���=P	~Q���U3R��$5zχiᥗ�l9:5;P=Nm1<0e �kفjCg��j�~}��Cu&�_dPۡ���j�`|S����c��S�1��Õ�ts]�7��Ԥ���YFPU��R�Aɒ�?���`.��5��m�v~6�mգ�Һ5�mr�F�p'yWf�f"~�΅ײ���l%N��Kh&�"􆰭�s=�8���?�3�E�l�����|&h&��{��:V�<��^���L��cp�͖(Xls��(�������8�m\�:.qyK��&�Y~��X a����ER��P3X�hu��Ȥ�ܥa����
�[g�\�K,~tJ���d[��+�.��q
����R��w��iU��2�\Q����Q�+�p���Ԃ5F���М}�/��s�<�i��~����i}�;iG~�:���C$᝼7�ml�y�%�|�8O�4k1�
����VE#w�['	i'f�?\B�w����UL����&^F� �����Y����P���3��Q����s�D'�3�����'FP��U�8~:ؼ�ݒ�C֒{L�Τ���Y�5��ɢ{������
"�hr�Ƿ�44(�d�z�!�O/Hi����e�Mͩv�{C���P�J�(�����2�j��n�HK-,��,�T�b�x�is�?V^��d���M�fs����Q��h�t��^o�Y�FqZ�֐���[O�� e\��k��te\�Z������/�![U`u3LJ��L}�1��0�]�� ��Ȇ�@�m+�݊`-W�q|�ڪD������Q}�Յ���lF>#z:������Uƻz|@�	z����A����o=F�!(si���	M�}�r��[c���g���i@��sB9
����2���"W���bE˯����'��>\zܔ���	���
e+� C(~��v�8Z"���dC!�w!��#���8�G���E�*7s�HC�\?�8X����ǜ9r1�o�!�v���4_!}-K����Cz���+�|��C����]� ������}� ބ�jJm>&�`�y����N�!����?T�Z�V�J�/�]j:��C�a@��?��C[��LJ��5!qi�#�������h
�M"#�6#�g�Tf7���!��E`
P��m2Td�MIMy7C��xez���7x�`��j��H�]�e��oOU��È��ݰ�b8�7�00Bq�?�B��z����b*��jI�?pn�sMZ�d<2q+��_���kċ�.#cӜ����j`��ÍB�u
QC�p��n�o�c�����&.���<�S���w�� �5��ps�t'D�a:����������k�·�1��'Ǭ3|7����ʽ-&�}M�S,��}+pN�xʍ5 &P��!���:�ԫݙ�t��H$��Y�����3c�ĭ��$�8	p�H:����� d����i�f��Z��/�M�/k�mS�6��ê���M�w�9bh�Gx�\�~�D�EJ�m� ����	�g6F�K�#ì�6Es���^>�+��>{[yR�h��T��ɡ0BL?�;,>���s�$/��W��ȡKs�(8YD���X�V��Z��JR��x��7՗{O����#��9m�yt5_�[xR	�p��g���!q����5�s�3��Xo��	B?���e�o�		�aP�]'Ts��̜��[9��,|��g�-���>�@;b��ӨNNJ0y0�~�Dh��:�`�ޛ����k-�Ӱ�u�`�cd���r�3�Ւ"�B��06)���8�8ĕ�%Kr���I���B�(���eXv�� �� �6�N(o>�/��2������"�1��+g �X���'a���n�v���x�Ĥ�u���N����_\0V��k�h9�$�>��p�,=�e��A�X2�3���z��j�L��&��ȀI��\hz~eQ9XED3�oj(�Z�)�be��8��m�qI�{rvH�:�&?��K���	1\N��'bW"�ڤ�t�(�6�&i�1%�Bd䶘���Lh���°����$�.�3�}X�)q�L;j"�	�"p�i��h�+ݔ���#+��j��b�D�d|8pT ���y~z�,�T�;��D1�q�t��i�6ʞ�.�#�����=�'���(��Cǹ:?�J:�K� /("�F��]����#讄LF'纎�j��}��\x�%=>Z�|�����O�P{�a^
��>jh;w�W��)���B��mB�/��A(hP��Ӯ��������t�L(;[����k�r*Z�`<6�� ����4Bd�	Y��D���AU�.4�I���[�R|C�
cm�kL�]�I<P���m蛆Q0B�e�$�Y��v�:c����� )�_���G����5��[�r���K�,�\��Z�*�z�iƴLY�p�"r݄JdF��*�X]Ӻ-*�ǧ@E���.:K\+��*f�f����(%pt�f�
�G"?������r���@Y�ɩ}��	,;2��1E�"xb�y���~����)��5���.��c�������%ư���M`ܾ]�j����/x`��}�=�^&�Z�`���/��G�6�5x3��`:��x��h�Y��t<cZ�ga�e-�DX�����/Pn�3���0"��u�w�/_�rin����f+���;Q��4��<ܽ�I[�ޠli����R�V>��#����s_��r���y���)g���=,܎��l����hq��m��1�8Qy��v�(@Ƿpe��`��<=mv@���5{v2"�ZI�`H�6TB�.�C�T*�3��E�J��%X��.�QNU�z*п��гI�h'ٺ/����*_�{����U�[ �T)=lR|*B��h��i=�U1�[qNp��Dη���Z@��-�z@G����}J��W3"y.���&�r�aS ���7�$�L�C�����@aX��u@p�2�bpTkI
l��Ҍ�ɑ�jh8�q�
�6-	zt��b���d��P��r�����O�Y�� r�7lߏQ \� 6��0[r�A(�ʭʡ����N8�v�	W?��J&��X5�L��̒���]Cs�j�-�U&M���N�?��vVQ����T���{]�Y�`w��1��
�$鴯�Mc�+- F����L��o �O$RאVv�7�W���&G��uEl��-Vx�N�$���1 j��F|�,�b`1�.OИ�Ŭb#&3e��ʲr��9_�Lb��8(wj2���+����)��t�c	p�voeј-5U䊉��dV��`�-f�^�R���k���EPЁφ��TOe�p�)(�>���q����N�8�����D��M�Ek�'����t�Œ�(�H�~O�*<�(}�[��i "�R�h�����og&�1π�Pc+!TtZ�Uh�^��|>����B ����� �sG��v����9�B?�\�`���r9 �E��J�8&�Le1�.���c��XE�[X�� ^>�Q>Y��������5��|�jf�\��y�tPB�K.��۾Ւ,=�wXl�f�@h�4��ռf�Z��N����������iڜ�R��"l}c�2K�7�T�LR&�@i�w���s�s�i��G�2J�R���&G����1���u��
�9v�yv�/������-K/��J7j��*;���]jK|��WJٹ����Z-G���>4du0�r��H�"�lU�N���#�I����g�b`Ⱦ����c��h���l��Y"<��B�4�����t���0��7[�E}������O^q�M�Dv�\Z�����F�f�ڱK�tw_)��Er�zȽ�:&�~!s�|��f�6{�+�n���ߘ��7�mIU��� 
�r%�a��{AxM�6��܉���v��M���7V�w/��j�;���.պ��S-�:�
���W�B�����1��`f��Z�0�!4|dY�'Uѕ�R���}^�D�&�p0�c�+z*�hp�Ѩ>�sԊ�d�`��d%�B�P�"��Y 2G�T� �%�vY�ŮF`��PuI2�
�ʭ{����U��{��Y`/���;׀�r������P��W吘�"s��d���� ���]��H288ۥcp)>>�4�'���<�s�to.P�	�܂�l3l$�}0�R����vSBg�)��!ڋ��J����%;?�(<�Wk�tz6�Y5s}V�z�K��$#����-��#]�֐���mI^K�w�����=�&��yT�
����bx�;&���s�N��u_̫�1��G��m��}O��sw��pV�f�H0�liu��ELLWF���m�h�'�U?Z�G��|Cژ��Ni��_]^���%EQ8��ζ�~D[}��o�!�L�)�*:�&��09�Qlw��C�҅�W�8�q66 
��-lq�Owm�Ζ�fe0ޙg�y5�L���Y2^ת�>�;p����w��
r �͜f�9*��٥��2}���N����I��AR3��>Ʈ���ۯ�T6�gF\]�<��$
�`�yP�9����e����t�UM��.G�q��Eܲ��2XR�Y���:d-z`UT�zW��*1�7f�a6�з��奌���&�"n�fǉMP�٭�*(�E�� 7�����������:�k��qQ�(4���ȵ��a^c�6款�|.�����3W�O��m5���cU{��$���(d�&�?���� [�H@���5�+
���Y/�U��g9;io�0d�J/�Iĺ�KF�0@^�-I%\�=��=ߪm���N����Ɲ�Q��'ݖ#PtqG68��cG��o1���� ;W���M�7�I�յ3lĴ�xX9t�ꋼ?�4�M�?��Nf��s
��*��刭����_��نHGAzqd�����`����D��r�ᢥX�\}N9�"r[��6E�
 ��.%17����
С�I�U�b���C�-h;$a|��?�T�7>X<����q}JI)�è=�� .�[���'n��A�W�P����6% �����o�aw�� ��ޗ�z�o˾O}��DQA���Vh�U��1ķ���r�eol�����IP��EY)c���pd�V�r0�F��ܜe���vn-_����G�~�0k/pyz�G�K��xk�蜈 Y,��:3.���f���A?� �bj��IKCOI��堤xk��L&�>1< _7�0x3J�0٭D�Z̮�]�"�y��t�g���pwНU��v������*�h�#�������-��^�
96�۟��P��#�Ց ��JU%�����{�'�(Y>	��6n�v#"Φ߸/c�w�B�K�.�md�,�✡�������`Am,�Xr���J"Nv�j�.԰�6�̊DF��#vM�����w(���+UchW#�D�h�ű�WF�ļa��p0Nx(�Z��Y�OeDj��b71%l�AT�%�fZ=p:�S�4��)���]'P��17�I����z�z��VB���`r6��O:�:���	Z@/3"3�i�Z'�B�G^�kG�=��k<��	�f�Z�o3�s��75�@
���Na����UPu52p.�rH;��������]���E8ʦ���F��&O0<��K��I<9$+8�)���(B(m���Y��9.}7�&�S3W�sd����o%R�n�hϛ�z�=�ȣg�PM�P�өj��uZ�A�OJ)Eeh�d��L�r&g���)����;�h�i����s�mpziJ�.墷?ѕ9�$�!d��TD��N�2�Sb2��h2�~��B�2*���B���1�nN�Xd�E����]|�����{������	��.�.���,u��~h���D�QZ����?*1�+��hy�m�d|Ӓ\iW�6'���h��I���>l���ُ�v��fX�5�F��]�U�5���"��"�^H�(C�S1O�X�*��X�y΢:�j����jv��t[�Daz�/�L�3�Y�(б�12}Y����n��!jڞaj�W	�p��V�������{�m��f� ̺iZ]ڑ7�}ǯe�|OV6���^
Ц��+��D��˯ٙ��I��'c����Xm3�kE��I�6��w�V�Ax�ͤ�i����^�=�D����8fA=���0(�n����==�O���_@�ۯe��dxU `��Z3�)x�(ꄊ�K���o�+��<VePSplP�L&N\�ЙW��;7~���֘�	 ��0�APF���3�B���9�[���J����+9�/�Mr�ݎ�i��ǧ&HS��(�#�%��0��X��[�<��|���Y�Y@�����x_Y@�ᰕ��c!���x���[��ahai��]�#$D�L���&6�e���b��U��ß.;�<2��ICr��C�7�-������"� ��'��YYLf�'^f7�����B���H}�@��2=Gc�������qBa	$����WȎ�����B�W%��KR�3��\v"��FJ�QK�@9�f�K�.4��l���X����cIc�c��Z���]ޅx�fҷ�B' �1W�y��`*.=��J��P�����]��m��o.ߍ><�Nt�~ԹX��7�Ofh�x[�b�H�{�F�;�;r[���k��,����1�Xq�#�/�x��y�4p��!�t)�IқZC�(���|��'�IP'�R�3<m�:���4Z����~(�a5��*s��l�r�h�$�j9�R��"z�3�8.��:��Św.08UQ?���ɘ�-@Ө}��ލ=�������ۨ�H�3&cA:�p�Ѧ�)���3�A\�W&S��K'fq0��^9�\�5Ԧ�ְ[}�g�z�]����zZ����v؊/hZihGa�<r�	�h�~�`wIhU#Oֲ� �#ϧ5f��ҋx���F��lj���u�h�si�9���� Sg	�r�7{�`�u�����X��s��9-s��|r~�@��w�*H�5��rP�9��6�KB� �Q�_�` C��?ӊ�q��J���߫��!��dzj/�)���dfVC�v��A���]^��Fx�]�Ed���Dw�-�"�%p 5��ƈ&\�2af	�1v�[S[Ѱ���IȠ�t� k 7ߚV�ϣ�j�0���Wx�#��{c�m��8Mȇڡ���e��� �ьG��~<@�B,��S�`���ӆc ��#��N��F옘Nl�����?�`}�����ׄi��D����"_bQ����EoO	*�¢,�轻�A��O�I�NoS�Td$"�#�L�JS��v1�^Wzh�\T��D�H���ŧ�5���L�K�(��6�����$�{���lٰ1�)�8巡dk�y`�ÚA<��}�tlIU�y�V��L��k'���M ��o�ּ�-�g����;�����x�G�l�I���dx|ĀP�W������xi�$]��!;�	�޿53
uF���� ����M�H ���Ee�N?#�R�}"/�/J��3t���g�xg!���+���OT[7�O�W��//����yp�}�[
�~�x��C���G�Q�j���S��U�&������㛽s���R�"��d��4X��/���@o8N�+\�O�i�&�b�/ƽؠ�m��꠳�w�eZ����m�捳�|1�]#�C}���Yk�CܷO�,����C�rq�b�����6�g.�~���K�>'��[?m�b��_m���c�^�wW�y�i��}��	31ܵ�=�֖ �4o���c��v��A(�>`����m�y���;k�S8=�θ�O�ӽ��U�\����d��<��]���q-?��Beg��Ȳ�FF��=U�"��C�6�E�{������ŗWA̿���W���|���Irn[�p�~-������A���u�jN�#�.*�7�,����bohm~ ��C���J�c�P��̄��0 	�K��kYK߅Qr ?��O�P�oۻ�vn�X@[`��G;;@V�_jͧ׸�o[�2�W�+.�� �����xE5��6� �N/�E�Wt"�N�W9=���nί7K�9⧄݄�0�hh�&h�F+�j��������_�{��2d?��Z���Б;��ZR޶)@����T�s��tj��Iu�!��#L����:g`�:{+�����"ڡ�
!��]��%g_$��/��u�lw�QĢ�1�/|?�̓�����av�ّ��Z$#%��*V����|��25�c�6(���+�5�\�k���+�R�%W��)wH�F�RF�%��C�?��������z���f{�TK��хɮqH��>gÈb��.�\lJ��}~��X�RA�	��0y}z;�FNa�c�v����|4�\ՃU�-pS��p�2߇�"�
�����#��=�CH�Xy�[,!<sh}�u!9��,w\��p�*堖�A��LJ{��k]��4�w�#�#j�%B�3�?��(����e9�=+��KfJ-�|$���+ Y�I�߇Vǌ9����m���Afť 2I�-��+���ƽP�h�@oH�,n}F9ט1�M]��BukT��g��!d"0��m�M��UU4����i�RM/�>v�ݷ�?����Y���?Qː �����o��#�L��?����z�Wj�����$�vB����W���]}���4�]��1+���9��z�7Y���j��L�wybm:..�b/��G�yZ�L$����'���'Z-�"zk��{���/66�ڒz��C� K~�K)!�[��VP;�Ҋ�������F"1=&�Jb�~�"@%�D g猀CK(�w��c�܋c�;]�#`�i�6�Y��:����KV�څ��i�M�Ԏ�Z�L��h�n�m���)GA���E���!��z���L�/
t,��&�H���[͝����WV�U5'���C�f���n�N���Ja��H��Óy���[����Ȥ���=|j3J�0�+�ϓ��Z;�z|��fc��VK�����Ǩ��A��E�o����#brꄇ���j��ӯ�	@c,LV p�ws���/�N.>��6��ѓ��j�ӞH5X�9�6Ƭ?�t& (����"n��N%w����y;{Fl�<vK�R9�|@�۸.� *_���߶�7��`�84����.�c&���]T����\��z�N�Ӏ�܄�C&�7�S���#+(R?Ǚ����x)|h���'��xp���3��I�1ioY�K��PΫ��w�aOQxD`f���D���w\|Fr:9��|+��O��]8ݏ#� �� lC��x��|y�rF-H�:^m����������;�s"o+��Xu��oJw����%'9�qBrZ�E���:�B�h{A�s�����;*T��_NX4:r��T��sq�>}j�#��?�@���i����ք��C��[�x��"O;��k�����R+�W{�^��d����%?O�m������ݠ28�q�&��j�Ч��MI؎w�b����}6�\�ҥ5ay��#���3'g��k��F
ڐ++O`c�~�s�;��ӄ��D�Ģ!�T��a��$IL.�bk&ݕ^�M�����z�%���������j5ɍ��m3r���=/�p���$��������4�I^@v�Ñ����,�Rk[��$`��̌�C|�H�"nJ�
�\��{UٛV�\�wL����C�(9� �3�}��= �h{���%QW�=-�a�ԗI?Ċҽd����������}�+�z:��K�}[�Bd*D�FN��*��#ľƵ[�>S<#�1}�+0���L<zݷG�*@&�0J`�c8t�|������-��և�E��%�Kf�����O�o}�%`G�D"�t�ev�(>=Ů�Q���'�9BQq�=��[=�a	�X `	)X�����/��7��o
�qX�����'�k��u�1<X��(��p�T),��)a#��+re�.���˂իۀ[���'�-��+ oc꫓blw�ɡ��#c��?�䫸�8�
up��[��g�e�C^岸me��V��R)M�r���=��7�܏\{����	G�g����G�y�=j�n���U@mц�织yM���L�P��A0����̅�F}���D�Ԑ�!7�rOR���*bc���g���·[@kv�n�����EG7|l?�J
��m���d/{3 ���A��MJ�������#�$4�?���?��L����ʭl�C�-f�_0��E����3�� &���.s���Ӌ�*<�,@�PV�&F���pb�L=8���+O�yu�@"���N����2P��u�b�@d��v��4X�c�C���v��p&�.Ve�w./mf�4�����q�c�cK�5U��[c��llb��N�V]��((��ܜG�@M���,KQڑ@,�#��Յ!p������Ց�����|,Cc��<욙�np*oLOt�D�`T0ѰK#�]�<������(e��{{EJ�����5�Ů��rZR�-��Z�7����N�������#�Ί&���g�v�.�tv�j���1,�tN��n)�K�c/t��(g��j)9Ilƽ��:��4�;%0�}�A|��,�JTM/��&G�]�	]j
�HXm��>�w�l������oy�����"��<������1K�r�q[�!� �N<�HJ�erS��^@��"��#f��a70C7�1�$���Hy����q�\9�|���U��zׯ�U!2�kC�n�x4>�`����[���|x��O��}��?K�=iC��r�u�`��E,XZ�n;�x6j��(��gI�휙�J�����ӫ='jйV���@�����)�)�[�>i �
��EVgJ�a�><�*�<%�q>jݭā����<�s=u�͏'�J8Z��"r3���Z$��j(�5�|djm�F�|H��?��w�I2
���u�/}��mZ�&�lNrC��{J��&��F��]�t�-������7�$��p(5vC@�3U6�[?����	'�����'p/e Q�`Dc���;��:���*o1�z}��dx7��jB�h�����ÊB�6s?PRb�Fh�WFXZ^���^�[����[5E S��ȍ��;%zy��}�@a
x|#?!�Ņ:�V�[�թ�UoٌG�kn
�y�h|�pP��jړ_kJpGi�sIf����S�j�M�Q`��Nq�'HV��oY��G���	�ą�����rX9�;��Sp/l��69D�dy��Ww*'5OŪ��l��GE�j{%���Px�Y�@��[���Z��r��H&U4(����޲N��O�ŗ���]a�K�+Ks�e�����1�=8\r������K��A��*<Z*4uS������5�V{�m�-�)��@��z$�c���y�[�~�@)�r�<���1&�z̡�&W X���죡[��I\҇E+�������z�s}B��J��j�GN���"��t犴��m�<�~%c�6i&Ef���VO�B҇�W�rږ�[%�v�wƯ>Ad��X�󥹈�6�\>Ѯ/���oK%�J����vP������e�V>
f�|8�u�d�O��0�,�q�����qawx�З��*(�S'w8g��jc��~:����Q��Ev~�nx�NW��u�pR��f�g���aY��ݮ��AZ9���]Řu��R�F[��QPW�kOR�(����US����jg�I{օ�9��eg��Z-`f=��EL�c�^��$'�RUW��XؓtV�NZ���S��NE�[L���/Y]�F1��o	�ɕ�"[������R�YX�E�7�N����Jx;�úb;�(���y�E�6��I��:D�D� )�*=�.1�`t��>��/�b䛴=v�� �]O&s ׈�iآ��c�ڶG���f:g���r�\+y�sD�>g0Jq�ۻL�3\m��$].Ýz0"5�#����ю�*A���w�;q[e��>$��Sc'�w������/��:���h�9�$�	AE"+�� �H+��N?�r�U;%�Z�����t>��6�
~D�h��悲���I�CT�c'{H�_XIp{�d�A�9*�,t�.�G�ZBcY�=f<3cp���U��+J'��ҷ�w��� �K�����s�`o�cr�����m����-���Nd�Т
���������j9�?m��e=n��l{\t��"��-��z���+��c�n�ߏU�]f���+X�EZ]�{	t�B���P�Y[M���;��&w�]�����Ͽ(l�u�����S���7a]`%8釱��Yu�=���i���{� 5�5[o�ъ[�����Vt���l��˸0̖s�C�+2�Z�A��ǆ�G���n�A^�0u�&1���9&¬u ��XJR�<����s5��9���S���4�����F�Cl��)6�S��Z�f&h�L�w�. 9����^�����2���M��"����_�<�*9p��w�zLv膥J@�ˑ2
0E�Wz�G��Ȩ��������B7i����	oI�'�rk2�$Ϣ��H��s"��$�#�-���i�Ir��	�b�f�a����zK�'lݮ�L�ٜ�V�&e3E�U+.���]�*6qS���l�k�W�W�&�8q�/?J�p6�~F���byoHLR&D����6����zNL6Qn�SѺ����zz��fp�P�>n��U��|������I���+�T�>��YRu,Z�-�����`�I��hF5B�l?6TT���}�6��^'4��I!a[q0�q�d�XȚp�i��鉑:�{$�� �U��H)ۚXfD��0R�t��G�ݵ�<��MV�J�ũ�i�G�i탖��� ����S'���Ԩff)(�<�+���\�q�b��K�pM����|��O���Q+h�C
]4Ce�@�
��(��"|JW{��`A�u��M�֜��̂g8�v(�DftZ4��h|�	�l�t[Pz!�\�4n�ᔺ����F�Dl/�{}n�:�����Ok��N��#x��X#.����	d��R& ˨�VB�[p�۷�M��CU.՗b8d�h���6��M�bDY66���`��Q�هu�w#�ϳO~��އ{�e˿�WRM����fC�B0l���G�[�� EFlptTo�܍�P���H�2��h}��۬�R߇�/���q����k�7����8kb ��c�ŏC���aq��-���ߠ�?\u�{���i� Kv���55ٯ���ߥ7Wv�̡�T��e�R�t�YS���\1��
�1���{ۤ�������%�v/~�[�؛o��a�dh�̉�݄��yk݈�#{�HO��j��Cބ�×��:�"�LQ����V�7�/��������8�
`��X���dV��F��pj"�E�,Rw�#DB�i�k�C�C�`��2��J�fZ[�!y�R��\d��(��n�,Wb��
��	�U	��HL��49�L G�c��s����5�D4}��_u7Õ�@ӽô~�U4�,�^>K3F�%B<��03�һd��������������-�,R�<\Kqu���IBN���V#�W�����m%���1�	@��'#�wb�K��SN�l.h �������Wd\�Ί�D��D���"���:)c/9��T�0h�� 2�a�<A�O�r�n�b�L����0T�xCv��5�U�������8rݳ�H�k`����w!Γ��`��&Ϝl>U6I7��.
��C��I��voV{�*��S6�s�������-@���L6m���t