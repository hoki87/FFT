��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ���������`z=�w�٠R�a��Ix2��6%|-\Mh~�.K��1ƾC.0_��9p��������3����)�(+<�k����?^yqKvc���9��j�Tm��O��
�9���e����G]$*H2=��@��^~|��-rٴK��75@Rz�L���{�����9gl�%�&��C��Ɯ�#�aM�yý�!�)՝a ?D�Q�i�Z�?��L�@�����y�_oB���(�ot��� %�^�)��H���rh��/=���R��(0DӰ:iPx?�pPQ��T� j�\iNs��.�u��88���{뭟r�h�Ɋ������]^;KժW7C���>���I5��с�����EmX�6�԰�}���\m����� V�C��Í��4 ���d�N��X�J��gg�nj�Ve�ax��/�����VḨ���D;��»�$��̎ �������S�Ro��\��Z�ȗ�b���@4R��&��9I2T߹��9���dH1o�L�snE��I3�bBn;�q�t(!�:�7н�̈.�`����Gy�p4�����4 S4��k|�I|x��g��~��x>B�1]�v�i my�I���!ܼ�z���)�{�zn����`
�w�9�����pb��G�����wa��3�ݩ��pJ����l���)@�v�����v,E�2�m0Ŭ	%�i�M/i%Ĝ��魬M�9�έk�2��`�p���c��M�_�v	S��Wly��="=�B��N�JA�5Z���n��膪��x��������.��$�R���u�`Nоd-'~�Iӎ���;�do!���{U�ݖ���IC}q�R������g��g�4�@��������V^ʩ&Jy�P����S&i#�������-���uo��7�]V�H�H�����[�p/������������k:�9���)��yB���"+5N�@PӪd:��t���cA�S���KD���67��1�j������ф���9M}�c ���b�x�:�<�'��I�S<v��6O�Y��2
���含�ܙ�8�ȬU�t�]��er���ݙ��_�q��y��M46��A�U������-Y��eDv~(;��z]-��l��~���:֒���^r�ɛkl�q�I �=�:w�,eW���5eT�<�YD-@a�z�����p�u��K�n�*�!�������G;���i�ђ"sE+�v��M���(�D\t\ہ��`�K5�i�b ����@���?fq����J]�̬?�z{, ����V�4k�N�h��k�Y6�xu�C�^��4�v2��WRK 5�<��}�IJ��`���رE�<g~����J����\��2Nns�1l��<���(V�C�/E����B�~���N�f��d��f ��V��w*��Y.��;Argh^<+7�V��+હ��0`��<R��!o���[U?K{Iػ�vVW�B��A9�-�yz��c�Z��z���������?_�<��1����i����J���	Tr��w�`�m@M�M*J=� ���������b�7��nT�mr���
w	|Ê���\P��q�:��8C=�Q��P���r����>�՘����?Q���_�(�I�n�m��r�|,�%�e�J�.�Y��3��L	�������ܑ��"����#��K�����\ٜ���:�.��^��ov���v��zМ�P�,J��1��	l�	�{DQ�e��8��d��LTw?X�+[�ů��A�5��1,_7�0���#J�q�h���D�;g&q�s�ɪo�Ġ��9ŻWLv2Ϲ�.�OOn��=ɾ�-�¹��-�Bk�'�q?�*�hh(Pk���W��{�St�\�:�9vd!Eo;}|J'60�}�8�S�]@(Yql��;�
 �ס����_}��<n�L�sZ�C^c�����G9�K	F$�������V����n)L��4��h�7s�M����g��8bM{�����ц~�b�G� �2�5$��O>П�Q�/�?I�+�3��ajc·�{R.nD��Tzp���ͫ<���[=���P������z�|;�˗"��5�G
I��D�<u,��=b�4eg7������é�<VYg���Ԁ���a,F�O���^�6Y;�� ���C�o�~�vs��;In��K��V�O�d	ǎG��:�r�[�o@��>o>�9\.����"z��&Y@jJ�����bu�[N<�.!ɬ�9�0�П6Aw�mi�[�Gʔ6��RDZS�Ns��o�F���妕3���\�-0-�mi�E̖۟�S��+}�}�]n���Y���*ir��SJHQ��u�^��B��ϸm�D��׫���*4(���(Z�;�� 8�)L&SB�d4�g������x�q������ 
�2*H�"���g/��.�g�;�b�vl5���c�����v�]�7SΘD�����W������=��qQL�q�qw�[��*|v(�V��ǹ�{2��SX�k�L�w�=�{ fz���^1*�I��KWY��]]��UpSW�?��
s�D���y)��=8�9%䄇D�O���FZ:�Xڇ�����C��ٷ�fČ&�3I�34�iu&g�g窭ס~�O����h�>À(�Zm�U^�L;��	&���Ï�I�Ŝ�A����λ�m �����Z����y��YxAǆ���[�1��S��Nz+�el��.�õ�RW0SWF�|��
TiV>��)�q�3[����	VM` �'����F����Za��W��V�C)%Uxny�%���T��s��Ȓ�<��҃�(_���)�.��9J�+���Bj��g����yB8�%�^`*�3�Ī���\�	�����Z|��'xbj��,�bp�x���V{u^|*дkڳ ��H^@��$�sZXZSg^�+B��+�zs�{�T�Z!�� �C�8�|���4��c�Py���o��c��3J���&������2��|�"
��
q?P���HV'��%}Z ��L��-1AU݆YHݙ��^�cʛ�U:��p"(��}v��+�uʣ�T\�h�2o~��~�!�N2��j{��2Ɲ�I��͹@������ܣ��J��y /u%͛`q�E�ƪ%,�^L�)o�h0'�}�Y�4�Kf�R��e�'��_WG�7��\.m�D��?��
�ԯ*,Rw�6]#\J%��P��}▵�ъ��S�F�>��@f�-�?�S�+A�u$�1o4�.��U�.p��,��������*4n�,4���s�`L�h�=$ �tf�����a���
�r�~����$b���6qp� Au���Jx�v��o��֕+�4Udb�T����5k�>G}��%=|� �"���r�'�������փ��-pEtj~Ǹ*�.����t��%�t�xY}7�rv��L�Mkώ���������3*l�z4�|�![��2~����g�BҚ�����Ɉ:u	g_�/{�Z?�������|ۺQ�j��b[��6h*�$I��l�ի��ߖ�wj�D�af���I��LD���B�:��B.j*�p�2b����p�\a����鶙�Z��l+n_��1cXu9Z�LR75b�-gD=}k����Yca������61�9|?��1�Sb���FQrH|��=���3�VIo��1e��$,��"�3��f3�A�$ޤE��*�,A#!T��\��j1�F�p@'���u����PZ{���%�P6���QnƤ�Z�ҍ�u���=��>���l��3�Ų���H9��d������"��	p+����-�й���á}� !G��8�(��L\�Xy��h�d�"~���Ѝh��w���}��x�Ɋ]�U�i����� =��-�&�0֌}B�������y[K��O�#��mn�ig�����K4��*��?ȁ@d�r�"z)?��R2Z{�+X��r��7ե��7F�������ZxQ�w�҂{/��	v-�P 芣^��ªݻq �����e���;I�u�
�����}��KE䂺��j�̼u;����e�oi�R/=9�uǟu��bt�p�9f��?���#s3�Q	��/�s��u�Z{/"Ғi-�*�A��J�S&%�