��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ����������=��o����W$qv��6�0�wYNR�>�u
��{AԎ��c�g���TCڶ��IF��rGl]1��[�qqa�'��������[�r��ԷM`��E�	e�Dt���B��fO2'�����R�����
�i�Sd"i%� �G�I��{� b_P�q�l�a�'�_4~1mc�_t����&u|S�%*EF�:��J��-I)�$�x����Jl�.��SI}{4��1a�`���%\yS8�(�e�,|)�Y��"ʨ�5��}r���ڠﲈ `�����'�􊚍�[�W (4�Ϣ�k�&pe]Ա~,���)��y�(�g,�w��s��xf�;U�\(z�Thڵ��ҿZ���Rd��s����"A�E�/$�w��RıEOp�F�Y�͘4/H�b�0��Q˜D�X
�E`���X`m�SEe�R��t���,�-��v���F�Zco�ߦ�k����H�#\C$�OT$rف�MP��<C7\N9 ��5'� .$����l��$�2�
_@�
��q��w��:d[]�&/MP�DG2Q=���c"�<4�ᡋ7M���s�u��J�߰�rL���I�;�m&��>�ۡ���v�<�m�t�h�W���5��|�{/
P�~�mqBE� �2r��8��|6H�	�:���YB����l��Էt��	@�����%��b+ְb���%� �qK/Y�]
3r(H.g���#S3g�^(�K7���J ��nOM�\0���\3 k30!7�`f���Ǎ6x)�an����|������9��$q���ӫ{�a�6��|I��$�pk]]�X��ŕ���k|x�Ht�5�B�G�&���A�`~��t�/���ė�l�ܷ�m!k��ʪ���}��=��Z{8l�L�A;�7�u��`�	Ǵ�.;�k|��r��aZ����5��0�-镃��2Y�qi���.?�	����Df��<JA� ��#���`A�o��/tΨR�����{{�v�̠>z�qВ��ΛBaAJZ�����a�3�:�QeE�:�"��V�W Y�U顺d&FU� D���� � G���G.|gC5�,$���~�Ÿ`#�$)�.#�q�⹳_Q�籡	}@�#x��y�� joQ�����c�N��!ݝE`��	�3L�3�7
��\�-F���ŪF9��_�_W�&�}i/�(�}�5[��,�$'�渓ǗZ���vM�_B������%��Z;�������U��b�
i�ތ�C K��ڽQ��/��X�:zz[4k��V��`�5��[6dYɑЌ8�Y�^�a�~��6����^?`�����Dh^
� ��v�\q>�i`���,0EadA�+#���i���e}M��ض�vOW�&f=���*� @W*׆��4Kb�'/ �%a.��Om��,�9���W�����yF�W8�,=Q�H(��ES�v�Z[�g�-�X�#j��!*y0zD�����J`�@F���XQH�����U�Pl���v\�v��gka��T�E�<��0��Y2���,,P(֒L�u������w
�� 	��7aJ�R��	�	[�: �בk�_dPq�t��RY�B�������$a�����="��4�����C��a�`Rg�,����!��i�GJﮊ����#a�y��"Y�-���O	׈�Lu�S.Y��(Ǘ�:����E"�A�K-�d�/Z�0A��6�}��.<�d����-(K]���1R�eg�\8%��� C�����$&�����ĉ��JNy%6"�x��n������ng�y|A��oдz�
T�(�ctT���@,�/�����-nTOC���x�j��Q�i:�0u�d�6����z���ǥ�x�d9 uw���q��) ����:�3���RXh\)qq��~%U}����g�d��.�>
��ٱ`t�Dٙ���OPn�Epu��z/DQ���ٝ�g��9�xn�k5� ���J �@�4a�(�C*^!'[��W޽�fZO��>��G�mi�u#5�������+oQ�9ś���6���TsѺXo��{�c���٣�k+� )������Y���&%����s�ᮭ��4!�G��|�Y}6-����d�M�P��T���q���6W�
!�3��xy�����d�u���c�Vw������,A�����.����"o�	$kZaCO�yG���PCkJխk���z����Cd2D�M[���_d�d::'I�)l�Z�"�3Sp�>���{�tЋp>�������~vJ��S��ߣ/��U��!��)�V�u�	{n���������'Ug�7�Xs]�k���E�("�~�ة�WP���-=���X��!c��=W�f��f��FH�I�}>�k�f�����c{3�*�"� 	9K2M���@�A'4�3�����x i0fPc�%>ߘ�pg�x�G���]�Q[��\��#���t'2D�)�b��\�#-+�w�(���P�s!�O�W�q)���r���t���+��J���ߊ�N�}��s��'��rۧj�q�ΫncQ?��.�ORM�~�/��9e���0��և��ݳx9���Ov�8��WP�7�Z>0p��v�
���8>���k�}�ȍ���h�����,�:�ӑU�a~n}�U�( hF����Ǵ�ս\�^&|$3������:51����Ø��W�h e��UP|	�X�7��ӷ=�S�͆	X��j�P���ס�b��|fu�]%�qF��"����/M�d|�	P��z3�������G�p�Q|�BWem�X�χˁI�\t���N��bk�X��&$ld��̈��{+�������b�)$DX�y��C�������a|w��A���^��2:i������>�4	(說4\��}%���Ps�zV�7�w^�-*�~*L'�Nhl4U�+��� �)P�QR���8�"?�K�Н$�8B��9�z��M�t̨��&�8���\�q��V�?
I!��'�<��x��.p�X�O2�(�-��o��J��V��^�*ꋳ��:ૻ�*U����Mo��=�[%��:H�7���)��wT�{@~��b��z��
N���W���p�Y��)�?�~��!�x��FlI���v�h�xT��nA�}�}�/Y;��.U���_���|�I�7)(<�0��,�줧�@X���3�<7n�:��u�u�|����o�!���%�*�Nq;�DƦ{ �J-N{h%f�����w��PeΨs( M�[�h�2�dZ~+l��Tz�-(x7ף#�#�r/y�R���bjiv�@�!�=H����N�89Y��]4~;���B�.Xz�l9HS2c�"������tj�vˇ���v��k\&�G�+KZ6��� ��8�;	�u�p��"Q¡W�5�ɂ�m�t�S���C�Ñ�K�a�l/\���Ń_�U�-�4� ��j0�,J���fQ�7&�͌�KeV":����tz�Ր�i�D`���q�����FAu9���_�$r�-T�hKf��D�r�!fH|E���3%P�oQ����=_�'�g2�p�I��}�Lz{}�l�X�
}H�؀|���u`��v�Q�̎F���2�{����[D@2׊<���֍f���@�0x, ��C�0�/��uM�f�����nM �`�貮 ,�!��H���-s{�����D}��%�Wy<�2��cX�_�1�}rÊ3L*/�m����w�@�T��ȈBW#��;����>��[vj<sȞY�l��C�nm�M����L�k�,Ҟ#%{�EQ�^Sʉ�L*�E�3h�6�`6S<�o�zu �]^CAj f�s�}9�����-��7� � �Ei��0)b�6e�{+��9�4K60$l�ЌȮ������t�)��颦�P��^Ԁ��
/��O�pb�_���ň}�^�V`By� qŐֽn�Z!a�#�Y������͔��<����}y�+F���0�KUW �����<E��q�+�`��ufS�
Y�l�Y+O ���V���a['�O9#�X(pQ�=�ш"JY-*P�4��+��!E ҩ ��n���5"�%�!=]��jn+�`�!$Y,[������jW��Uc�VJ �G���}�\��;�-�M����ڴ
���Ғ��b�6��C̤p��c4���bL%���rZf�k�A����.�UT%��ayF>�@��ssvFC�|��A�ro~��]�N��但㷝��?���Ԝ�̏,��Mm�xv�~��x����$3���.�g1������=a��>P\9���k�EI92 �^�qt�1�E���av ]��ٯ|���`��_C%�p��u�E$HdJ���-����Įꎑ�+�f����[���6�)��dRrQ��&37 n�@�BRZ�n6 ��	#�i)/�zp��jCX^����(��-*I&��qU�ЎJww���g���V���-$	 �#:�����!߳lK��Pi�SuZ=v�r2�{�� �����hn��}�������Uqs6�������cSn!���iW-���kk�;�wT]Vy�L͕�}�abK�^���V���0��>^=Y攼�J���'Q�ȕs���=�I,ɱ>�o��}Y����Xئ[x�U�2�+��<��y�� A��-���d�`����d�#�,W��G`5�Y�z౽����?���}�#y��V�+��w��)w**������i����%V���zq���������cHF��ǚ�;��&�"��l�|��e���Sf��N��0�|-���g�Hp��0�4I|9�?{T'(��J�C��*�ʠ����JB$�[X�uUQUnn�3�FGN�R���2�'��4$s=
lf����$XM�ڙע��1��,���F'{�h�9e��,���oB���R�����4Fj��d�j`���'C���Ռ��O :}3dS[
�N�:����_|�T�w�pPTֆfx�T��t�̓�%�&�)g�
/��"�"�N\���aZ�Je�f(]�(�Q�S��d�����L�B��qn,�ێ���Y�M���;�"q4#��1_C!G%r3�=�c���0sз�n����<0y'+�:��j~�Yd��߆Rq�FE'z��.�����T�:Fp	cW��T�H� ��gbm�J.�N���&���4T�>��_;�#f$6Mq4f9�o�j?e�.���q5UA"XÈ�x��-7�=��3V���]��!#��h�4wV#��9�۰|�l�Q� �Eo@x���V�c+iz�#8�|��m0\ohu��rN ��d��v��ȑ�'���5����}���3�0Ft�`/+ăO����i�~���ǩak���L�B�^q��M�Sv��Uh��8��D6֩� ���ʒS�'3p�x��B�ݗ0�b)��'��O��&ݷ�z�����ɟO�2w��$p�y�_���LA�<t��c��d��
���VR�.7���yn�|'\��<��=�죣��&H�5�+E����8��=/�դlB�:�"U´�.�K7X0>[�?!7�U�7߹�r�߭wy�X�ε׎�I&�UT�S�f[�ld��4p���.z%ğ�Q/k�|�����6���c:Aͩ}�B���3)�#5��BaS=)BK�V{�*o��R�RL1�kh,k��,�����0�/������c9���̛�����Y����o���m��jE/Nh�¸<`v�uV7�_f��)�֖fM&��6���6a���r�h���H���7[�
��P�C,�
��	�nk9xqg����d�p�"������M��qu����U0m�`+="�5X;݅��	�VS	�$��pg��|���n]x�	�e�ȍ]�C1��ۼic{�T��	c�m0v����4H�(��`8��t�Q�H�2���C��}}��V	�9;Դ��Y�r�E��N�dPS��ƚE�{7����r�%������H�s0:QKk='���U+�/�%��+�k�t��lGJ���qTg~;k��Df����ŉ�A�6z�g����FLh������qsp��6�V�Q�%�և"��j}f{s_��tN�6�]l��tVd�>�Q�!��0) �WK����2� �{�<��cA��m�-���4��қ45\������| �	6��D�4߁d���Ҁ�X�����Z��a��({�<����z6��ʼ	��L���j�c�*V)S��@gg��m��h�Eu�+�x;'�a �Cb��c��?����]f�\I?�mFr��r�~>"�!iޞϚ ��<c�X���WH4���&�V���M'�J���:�/�����Ϋ!�h�~��fײr��!����� �R0U�ݧ��0i-vL�	�zP\��"CZ��e�#��4|O��b7���Y^��x
L�d�,�� �m+�¹�笐;�����Rdۣ�
g�E�������=�����h�	��0M�Y���z��/ڴ�� fM��Q0H��N��3��@�4խn	��+aD.U��w �\0�Bj)��G�ύs�0e<��E�I�ț�_w�r�"����TSԠ y.7|�~��!����N�0� jrg�d0NL>Z���+S�6���5Z�?�g��H�8�u����x�d��*)!T�\��$�y�M=E�ѵ4��N�o���TZ���R�?��8�z]�y�97�e!�q��eC�4<]6i�kZiJT���H���o=��s��G/�\Aeu��l����T�]�.�q���4��9�d��R�O}�[�۫��Ա��ˇ*��Γ���5j�,�@�s���?��y?����dA˚��Ŏ=l]|��!���#$)1)\5ۋ��[�0d��f+�����ɐ�Q�_�����R��� �D�X ꕄ�Oj�x�������t������WsW����>˪�Cl��F]8)G�q,ÿ���@w׈{���3+/{@�OW��	#��K��2�ܫ��d�����'��]3�1��|�q��G���G�n�E�$̎�J�S	x��-X�ݡ��+Ώ�E���TB���gH���CEͥ6Wk��V��*b�C��#��t�$��#�79��Jכ-��Iwr|��R����)�6
_їw� mz�e^_��������V�4(�X�]r�d8�?l�oEy}�~N��m^�y w�j`UbK �\�^^js���3����MQ/������@�8���Z�g՘�HS�2�<�>�zW�2*|{�ޓ}Ԫ�y�6�!A�E�q�b��!����p�^1��	��<��&��u���Db���F�2ګD�'�Q�k�6>Uw�����0�B�6�(n0���N��������Z'�]�vT�sM�]����g#����)�L���o��$/g���O�^}�g����� lџR��$?i�(�뫢�}�����]z��Tg9	K�I��E0ߨ�����Gظ��b׽3�Q���I�<C����T���P�:�)~��t�]L����bE�<���`�D?���[����a3��Ѣ����J��`sQ�T���u@e�kST���	7q�{=0q6"(!Q=Ԛ��uG�\y�a���T_B!r�^��-*��d�D�S�+�ܳ�4��Q��=�˗e#8,���9TP M�? �� �~ln����t�2�d��~
�5&�UA�|�ǔ#���_����?&���J�Zol	4q�"�LJ�����_���1|�D\3��g�5�Eye��Qy�����܋D�믆Y�������?����m���]�V�{�X S��2�+��^�͵A�.E�n���97 �`پ�K��9��2�R_g���%C���8tb#�=	Y<���f�L�\��k�Q���a�(V �F4F�'����h�a��3@�z���򛝺�+7@\��b�_j�Ҷ&»�䧒M@t�9o��n.i��?D����銋�䆺E4��u�r�]�=0ީ�~O��=�4�� ���+�-��(�2�R�IEK��2���z'�h���c}��)���BC�ڒ�w��6]< �髤��n~.0 �c��Q��~��e�x��P׮M���@���|<.p	~Z鋪H#���iJ5b���?E�ꈩ��
YI��ś*D��R������MJJn�K*��n����f3�eO8ys FqeAF$eh5�	�z����w����eϫb!\֝��_#RK?�b(U6���У�0'��l�-�cJ���0%���li9lz�o=.�ӈ�%:�aX�WA�9ׄ��,��I	���g"m�9�aο֑��e!�au�P)�݈���'B8��]��hT﫮]�=�dz桌&�ơ��L�������I��QM�����ı!���R|�ݝ���~����ګC0���Җ  �d'bg;�U-{�-J �{m�b�v�m���?SثY�;B׎����O/�	��iv�i���tJ��
��Hwk���I��jlf��tv��P���i�K�=�4h�읮�������Y������i�V8�[n��Wj��dP�6�ߑf�wkbx��Z �?G0l�������7�"���Z�!�I& �~uqF�d1Z�OX���I��dN�=�����J㺬�3'_?�O�b��i��C[:�Z_�D��v���=j�&^��8��K�7�&yx���vP���L1˘)��W��Ժǳ��"~ʁڛ��Z�7g��[~�d�{���D�U����,�}��[������<�}aL����T�K�8�^;�2�o�-jT/��B�@�dj���u*Y�Sy�c�����[��tZ����}%��A�)�K��\��j��i7=>M0�S}�3���9����/�5o�&ec�O*JeS2G��P�Ku/�*��S�|'
�����N4���eRY�zY�Ƥ'�R5_�T0�T�eL��l��zIK�GJ<�s�9���	X�O�_<���U�[d��֚[�J��QMP����
�fB��v(+; o�̠>%k6'ܖpٸS�=+����+�R�*ٿ��c��,>w��=�Y��As֌KZ�Fm��2xr[!�V��!�k>�� �Id�!X����D�LZ\�+g��F�\�pUT��W��@ �2׿��U�>{//�D+�����b>�gJa�C�sb��⫋ ��c���/��3�8Pq�W����7�$���1�d)Y4fI����P�V�tŉ�ݑ�5�i�+�z��Z��s���Avw�� T=6I+�Л>rѧϰ�:���I�AU{�u�<�\�i�# nP�@D$�й�-}�u(g�`�@��k��a�P���<�t��L�Ë\}�z��j>F#�%��è�r��0P#B�A���4,l�I*5x��k��՟�p@�#�D�K�ŖJ^7�H<�����v0Rz��m;���}�T7�:8�7�d����)9���5.M�d[z����9o|�}$���>���Z��FV� N,�6�:����ǲp5L��[�>jl*�H�I�F1�1�/�-�8��\��N��2�>x[�}����>��31)5F�nX��+�Mr��oi�xbo���(Н��6����������
*��|ZuG���񁴸s R�Ç�XrDΜ+�w�a����t�>�yX�|-����M�i��>Kk�n7�57mu3k���Hw�Z��oS��,"�pȷ�*΅�`�/C���5H�����y�1+��r�/�����Y"vy�kn���8��9�*&���ƞDPmLT��-�6��x;�#U��&U@n����Z�*HLm�I��m0�ᝓ�:����+6)0�:�Oj�'���{y���(]�m^ܺ�J�〣����r���F\��9{��mky.j�R�w�����x�ƾ����:���W�p
#�g	�������{&��yV+�'8�>���JD�%��ͳ�S�ڣ��*LELkΡ���Z�J�ӌ��HzMM-��R�);Cl$k��ӭq�z&g�����OȆ/�#��N��5iׂM��wZ+� ��U�s��ǔ��L֨�y�Az��C�K����;��:�D~�7�y�\��cn����AIñ�3ei�ʐ���\ٟ\R�^��ؤa�8�r�PX��Ȧr��t]�i;^�yo%7��U�g>(Qވ�_1�B������5���J&D�CC��P��$~�~�p|d+��x�`Cy>���ܜ�-U|[?�9a(��c4ܼ�g)�v�r�/�(��]��������}Ÿ6swϋ� S� �6�xp�#r�nz�m%,y(M)/��2��\=�e�]����>z�*�7�fw���.��E]��ϫ�N�*���?����X�)3�1���&�u����N<Sy�^�VGX�@�&̡
���{�LJ�zUGQ#ь�ܐUD��EI����{ç�ڭ�J�=?�	�c}��j��-lHVGx�oـ��蔆��=<[kM/*�<*��l�����6E���Es��y�9z���u@�i\�?Xi��ʓ,�ذ:��s:'���A%�L���f��/�c>D�@��4(� ��郕o@P������x2>��'l2�E�,�ğ��'�k� �J�����9=_�X�P��6�C�"��%:��J�Y����[kN���I1��}/�B��l�}Y�|���b	B����֤�&���±����{k���2��E���򱱒�s��(Rr�$7��ʫ�����m�F�+
��QW��#��_c3�jˀ�G9t��Heԭ��N�]��Am g��g��קN5����D�;�ݬtk�(�3��b����E�~yT����YD���X[�0ݩ�j�0�4��4˾uh�~E��j�L�-d�'��]p�&o�U��语9}5�A؝�wǝfj�����b�a�('w����� �\�q5����(G���dn��3�����bN�Nfc�WE[�_��a�2iq<;7d�t�&���枘���ռu�5Z�a�$�l�\T��:�9�Z{$�d���wE֟�,:|]e
H#.z���ۤJ���a��u�E°T�b�Qm6�U�8��M~�ہ�:+d�ۯ��}���Ì�R$��:Q;�t{����$	"={�X9��}*xS�VX�#r���J�s6����§.�nJ-ƫ�I��o�'k�nۀd�A?����!�!99 ÇB\����QE����0��ۡb���b����S3:��:���hGD����X�§L�yNK��AmK>���.l�(�H	<��G�/�8�eaX�轓n(0*��7�N������ߌ�4tL3��Iu��Z��祧}f����VQ��B{���~=k<����^���y)&sQ��z��|��}Y�BJ�*"#/��=T��0��{�d�հ���e��T[�ů���	尙'���OxEa�p��Flu�8fV�0�ӑ�����{�����QC��wx�VU�ae�SX�Ї���z��-�A�ݘ�&�i��&R��n�B�3���b���.S^��fdװ�г>�Ε�Ձ���PD��Zu��m�lq���]7j���C�ւn��7����M}����7�Ĥ�3��#���8���Mv$&�mv�%=��{�)1��:~<J�������]�X�K��˨��Id�x��6<���~��7��F��Ӡܰ�$S`;�gx�.���d�x���F&���̢���'��呀"�N�6�Σ�n����ȫ�
zn!������"�H�aJ���zȠ�g,1=��Ӟ*�8E06~�� ,n�B�:�6m_�9�NxDG�<�3������{7�T\�5�m���LQ�~Qs�8Ya�]hJ\�u�y�WT��q'��V5���
]<�d�e�dJK����̹D��?�����/u8��:G����ՠ�f痧mn`��6�Ӌ�Y�z(u8���J��v`�U	��%�����ݣLX!T��ϳ�,�5<�rdߍQ�M�~�P j�';�EC�i�+Ę*�5��Tf�쬡Y#��x��Ř������`]�w/��7��]F�s%i�&��+���������k ڻUA�"g;� q~Q���#U�*2�,[0E�o�]?���y{�o��{z덳%3�	*L>ӱrS����R _dК|��x��8�Za��eD��_��P:,C,����9o���Ԡd���b5��`Zp���"���r�x�"x�~��;�q6��$N�aW���,./_Ժ���S�"l�������j�HCM�lQ�na�)���Ìli��nLV����[�dF%�u�����K���f��آU���z^mǥ��� �rLT:aH��^,�PL_�C�l�	!��
T|�%����0��G��'&�f6�Vl���� L&� qc���\߇�{3���7��ٵ[����P�W" O���J����wk���D��2�pK�o�9�l�:�񇐃�z��ע��Z.z��#P�D�FW?�k�؆"+ׯT��DQ_����~H2�1�A0�<I���Z�T\;�F��y�����~�Ob*���Ɗ��(��r�u�͉�1���?F�䛓�KT���v�~Ǳ)w���*۸A.���j�)��
HR|<��!�s����CT��-Ch����a���Ȭ��|Ud,�uT�h���"���N�@f����v��"m���ػUhdV)����m@A�ގ��I���3	���ʿ���z�?)U�v��u�6l �oPBRB>e}�G$�����|������i�+*gJ�*��*�@���)[1x�B !�?��a�
�2�YLpK���T�Pm!0��xc!� �����;�I=�&�i�gw. �\v�T5�y���U��� ��rC\Bh�஁�F&��b���$])���7f1S��^hX�o�����X�d�1{�=^+�7���@zF�$F�t�fvt�|T�R�����]&�#}f�����\5g ��WR�j�+�Lx�N�ī���~Z)���-���Av����(�zg�,��F�IK3'������.6(31I!�`ΐ���J���h��E���~� P�/U��K;$;oyr��2G���/�]���aUl��ͼ� �[���_���T�c��;R�X,�Z�{FO˞��6$��m]���ˡ�e����i�����m�4�/ԥU�;J5p��pÝ#��_��վ�6�M�c�+�����b�!_\���`�ht���L�j~��xW*FEB�BiP���9�J3kM�X��8�# ��_Ufqb�w�M|�� ��W����u��8�i��[�l�oޞW����_��}�*b�M �ٵ�ן��Eq��`{�H	��R�c���4>���NP�������V�ᄴcs?0M���kɅ3M�C�Ff�WFM�z��Yh�	6!��XnM�68���KPC�� ���O 8d�tD����d%~43*^l�O@~=��G��YU��+�vBa%+H��>� ��p��x���UaÙg6R���G?���c���BB�}��Fp˙�+�����:n�ٹ!�7Ѻ^#�q��'z�B?�_>�8y�a6{�oM����^ݺյi�Gꡂ�(���k��Y�����_4A�M�̴��L67������;�.+D ��?X�#g~�;� q���ce0���-%���{Kp���2�Þz��=��	�As���]�? ��8Q��<��Em�x9�!+P`ԟ����d�$�(*#v�Tf�C�tD�oC��dF������;ƊK�2uX[�������t�y�DY��u�j)�;�\\�dm�r��@��Q�gޝ>����_{,��YO�}]� ��Ͼw\�����{��:��a�&�R��o�^��׹5��]��Bas�E]������(+<�T�KcDFa���P��D�`�Yv��	��Ǔ6����v��q���Imٷ"#�*�v�5O�9\fP�xv&أ���:�O����U/�m������V�5��<嶹��ލ���,�rgf�A\�{�1@ܖK3���<�Q)؞6��^��?T� ��W"����!�������ƴ8�ENd�8t5��'��1x�A�tON�N bs�3'�:'l�����?���5#�4d���20�t/���X�m�P��uxuu�hӪ��[�\�r0��@���(�.�)��)?@4�l�Cd���AӋ�?��J�[NE�!�\�'!��L@ƨ̼�D�
7��=�m��^��#z�C����S-���)�����!�5*є�N�����ttn3������vHլ��=�nV`P:9{E����"�%�m(��|8U� "�6Co-�M�"BS�QNј���k�fZ)D��w]�E��r@Qۙ��U�����çR M�E�����@zc����|��B�X���5�F���pp�3)í�e|�՗|��V���;#	K�����/S� ���Y��C�l��4��ըNjk��+I��M)x-T%�ͧe������ ��h�n}�$���+�`��.>�$�p��j=I?��"�0I�1<���_��/z��嬫p�-a���ˇ0\�|��Au��&� !k:�Cu������#h_��朒�,7W���D����t�F2G����";P�!����U�fv�w�'Y�X��T�b�隼)���Ʀ�ne~��ɌZ��`�5B>��Jq�VA�9 �[wQv��t4S�����l3G)�e�E*�;a]�6)̀o���`�rT����p-�=�B�Q�=y�e&TH/{�e�%��u�K�Fi(%�3�h�q��F�
�B�����daWK���Z�j��<��s}�Wk�1 ��̘�\��7: )�*�[��	��N�2,�����]� L��݆uC��
�o�Z�z"����%����'z��M�lH��Z��&8Q�LM}f�Q/���|#Đ=ᛢ�BC%���b2�'1�	y�L�Ȁ��t�?�8�
cױ�������q��2�@�Ħ�D�3����0��U�^�q\N���ҧi�C�9�K�y�m^�����rgJ���4,�Z'�ΐFXjx����q֊q=���	�Un����41x3D���?���'��n<t�6E`e����U���U�`e�ͱ󩵜H���Q.[e���a�'ǁC����V�X��t�k%*Z�)&�G�My�N �ҭ���<J���q��9U� 2��X=�������-;��_\�\�'�t�"�'H�{9p;7�ͼ�^�2���J?-w7��[uU��'��a�%̬8n!��%o���s{j��R���ۯV�^U%���������������0�nJ�4!��D�o�P���遙�vz��Z����X�s�ͅc�W�P�ԡmu��q��7��i S��iR�"s8|$l�n�5�݉�7�"2ᩮn��~]�%��v�w�NH���UU���e�k���v!�:�ZP=0Fc k�eM��c��Hn�˂Xψq������fq \X]}6/)�$ҧ5L@���0�{�~�Y��2��2���] sP��7����s�#[�e.�V4��vid�l�N[6�(�o�+?3Fc �*�#�@{�5��6Uf5�A��L��D�z��BK�l�8t/�c#ɼo�jA���Ufv�D�B5or�"�[cCf��$�.�7����Ĭ�wV��*�*\���G��$*^��ɲ�xɱ}�-. ��^>�5˻se�?�����kkl��q���r`l���w����s�4Ij
���8"Ј�b����ML��,��x���P���E�Ip����e�s`�K�}}r�޺�ߧP?k�dB�*p� � (
�RB�ʒ[(�f��#��@a��bD)��С�w�˿eg����A��'�c)HD�|i��jf�����l

Kئ]Qڟɴ�@�0�9(�T%*������e�&�C?s�A�u������6ǀ`"��c�G�`�������_t�K�逆�w��e��t�����A��;3 ����DC�)A���Z���0������FG�u"m�Z�T������o� �M�2��Zf20ߪ&r`*=�t��̬��<6ʯV_�G@+T��)��2#q�篳���f���64�uc�&^�ڄo �y
޾�'&}����xS�r⾖��O=J�������$����� "?���כ�$��u��oW�O��
ŗqƀ�t���,q�2i�����y(���,@��.#�GS�0m�p6t�`r� �S���,��#Ƣc�t?�IY6?��59
��k� ���fB/xI��m�A]�8��W����G%q�1��d��C|ǉ��|s�c�}N�ճt���2����Fe|sh�L#YcS�ք�����5�*Ā_a_�,�I����c|�_���G���^N�A%�����_D~3��"$�[>P����JQTW,����8��i��s�����\m�:~�蜺��Ge��Φ�6}#�r�U�=&�A��4��&�9l /��F4����ȃ�TW>�����A)�({�D!���-QUe=��y��p��B���ʳ����o-/B��Jc��g� D�L��tO����Gv���f`�.����+n`�J�F�!�*a_�
d�����7gē�2%/Aw��j���n�B�ׂ���&V�2�n��䉐V�y�Ud�����j�Ũ�n� �}�T��r�q+��n���?��I�G�f�j�� ������7"h6Qx)�#��eD�W��Q��免z̄�	J5�E�l7�YJ'� �Q�]S�pU�!�H!��V��󜉹��g������v��@47	�+��:��r��N>sg�T^��bN'Nr4�(�a�k�J�p�yFQ�bВ`������ �z�Z:�9j�)��LnЁI�.�Z2���u��o��U��X�����w	Xq��'��d�V�����,�Uxx��i�Jj��~�۬Ř���C���x'��w�7�(e�B
�v<D4�g&e^������O��T��]��m��1����"H�F��0���x����ޚYY'i��<��9NF�^2ڲ�����GZ�^Bu l+Lu�^s��v� ߼ìP�����ZB��uf���Y�%���2R6H��� �w_Y��a�[�4o��EF�k���:)ܰ4�>F,&���!��my���UWRL���yȕ�0x�J� mi�plg��Jd� r��w�<���E�M���0��O�2V�]��J�^+>��.l����(�o��&z��d+6�'٘i���ݑ���q�b?{�dG�>�.��D���H�޼���M�w�Α���YS$uk1|���9K{Ns�b���r.1��M��҆�߀L������\�K�3��Ý7�Ԣ9�0�&�mS��~��3S��Ө]^�Q��,�cT�H��������(\��LtH�/T����X�;�r�Е�F�͂T(�?j@�?�G�NZ�����oy,�͈����Ź&$��Q��d��p���j:�'��;\�Q�q8b��}�U4����!,Ù�E?}+�?/�3��Q��[���m��6^x�%��Y
J�?�2�ж����	~�kv��A�S������V/| ��Y�<���G@0�d[5��Oٓ/i��n*u�w���d/D]S.?an[�3�m��up�P~�y��ۻ	v�$X�L�=�Bu�)���[�T#`Q�c��V�̴6�*y:�фu��d��$�%��!�i^����kb��B�Vp�G�8�N�á�1$}髺�6��\�%��[��ϸ��Q���~ـ��E�s��� I/&���pԑlg�M r����#�/o��H.Rw4�z��������'4�*��j� �N>�Q[���.Y�0����2�9@\�D�U�>+9U&�C�K�@�ߐc[J���9:^Om���,�W��3CRsW|�eצ^N�- o����]Z���-��<�dDQ̗n＊���Jq��<�Q�ڌ�MY7|G�L~�u��㠪2ԕC� D�ʻ�DХ�x�s�>��XGx검��5+�!� ��#��(�� � �.���"�Ҡ�0�@���ZOg�]�������#�y=˶��u�G����]`�;J\lF!���/�׌�[h^e*[��$����^IO��M@K�Գ!�~�Ah��uG�d��;�\��k�dǩ�YpGr���G���[E `M�qOp�]6��W������G�e�F��q�=���S�z�`�����b��T�C��o�~[w�nn�-�����%m�8v$��{O��$X,��� ���Vu~��N6I�����4����sW�&������y��Jix��M�Z�y�36�fc�io�P���ܿm^R>�:F��pu�Zd��scYNRR�M����9�`4�˛r7�\��#1�f�Cc�\�ߕXo�w[@��+S�F&Yr��뚐hCTj-�,(3���3Y�Q��3�J��Jɷb�q��+�qT��ѱ�
b��`奻+XWHZc���i���	:Ӝ�8c���r��?���D������Gv����mpuB�f�j�.��(S8�~���A"�1Z��b����d��\c�ˊ����� ����x�,�B 6Wp-=`!u�0qe~�п�
H��1㶮da�R~[��� LşF�zgk�f9-f�{� En@��8��)	��-֙lQ-KrI�vE�E#U�ׄ`��''x�DH�����Oʦ8�&]-�q�˨�j�����J�7�Ѡ[*��s+@8���o"�-!D��Ug�> �t��_Ϥ7����9�����[�1���|�&����,6�z�ฌqUK�h�'��ԏ��B'|�ߞ� �����}
�D��=.�?���4���S��ke�U��X���&iDV�˓�H�i>�����_��) �y�)�@K����U�&���+&c���Y;+���7�O/�� �Ƌ?W�4zT�~1�C�M�J�֖朗�ޕ�Ѕ�e��$ⵦ%J!�H��2��,����4;� �H_8�Q�
��G�	ʹ?�Ŗ��f��`0����n<��K�\�%��X^fv���
F�'��t����P�lU��a7?��
�d����뮊,Hk ��(V�mT�jp��W��5��-��1n�;�JVe�B2c�ъ���6���&*���S�Ȱ�c����O��P�%w�a��Hp�Ǎ�c"w��y�q_I~���$`y梻��[��x8�w[�K��J�3��PW�L�b~���1_qvzW���ԟ'
DI��v�E�,: ���8��<���J\u �r�z�"������Y�[�;��{��wo��7��|��XQ3�����FN_��q������?�Z�}��P�1��ϝ�R)ؗ Zt�.❶�b Q��29T{���q��������ㆨ�$_d�ۧ���wiQ������A��ضUp�Csm%����с0�<_��6I�N:Y�<q�Ӗ@���_/�Y@@�)�!I�S݀�f����Vs�j��2���� C�fN�9L���� �\��LZ!�a���<!�CdI)�����+�%��?D�|���f�ᦵ[N�c�/�����{ yv�E� ��P���b�~� hq��_���H�"=�r�4__��}���و:?Kޚ���,)m�̨q���W�g���~r�_m\��-���L.����h��R�Fs�� ���M
�:��}�}r�<F8�����Ay.��vmYz��v�*1�A�
AF�gV,��1��C=��5��F�>{�E�i�&a7散�8H�w <g�P4 ��-�s����+���Y]sV�D�&2n�P[yF�����ԃJ�U��5o�u�Ġcg�N����o��v���Ă��=�X;3,���A��pϕ|B�����x�"�o��/���:�v��'I������&3�ff�I)�A�v��⹎�sv��鷝t�4<������Tm[P�Q�$�Gk�s1�:�t��y�#Qf-�a�7�H�Ӎ���NV2^��W�'�Ҵ?µ/�,�6�X|F��o�zS�(���A����J�ޜ�����E��K�mT0v��c
�X9F�
������|�����$b�_R�;U���Lj�В> �M<4��5	W]<(����>c��Ɉ�Ry�%�I]z����b�$V�t,���3� `���b#�
�
b}>}��^�O�v랡a�*�5��{����%3�2���?�6��z��h1�~/�H��R�>���6l(���~�I;}�|	G�j ����/��l��v�M���&��l��twj�1m8���[Y��r���f2��0�1f.]�R톕r_�]h����eG���q�Z��>ֽ�)V�&g������$r�_k�����rJ�S ZW\Z���&�4T��!���A�ND������8��#���T��1�E��PsEo��S5�:����Ē���se7�ٖ��ߎs!K|���"�[ƍ������\��:3.^F��u�5A�&��3�ܥI��P~��2� �jJUt�o߿��iY��1��v�U�4�IRmfa���(�,^�2	�񙄱�8��e����$�a�n#$ޮ��"�Zi��z� �x�ʫ�������3��N>W6Re�n�����Ý���߄� �x�5ڥQ˅㥏J�n��-�~����E��K�J��33����q��gchjB����5&�n�Iu��~��)8��T�.��X�bad'L1�<q�����eQ2�46BgO�����T�Ш^{���>�L�O��:���Y{�ޭ��0P���@�7m�O�E��oe2��#V�\�Ӧ��^!�'ی�X%ԧ˸� w�B3��.R��K=4�$,|����7��g��ik�ۚ�\�Ϗ+���<�7��Dkq�+��[����x:i�a玢�������D�I����y�?ˣf=Ju���h���L�7չ��kz�aJ?o�D�M�w3�t�>�_e.�<�� qZ^T�,Y��M!�e ��f�>�*$R�+�h�X:��B�Cr�<|xvuI?o�ɑ�*{��2=�!�	�o�n�lH�@���j�4u��
0ێ����E��z�1lݯ�@��0�4��^����K�������Ǩ�PCYz�F5,Zd��:��^�h�c�k�IƸ����m��kc"�-"1�=i��=ʙ�
J���?� -d%�W<J���O����n�s��"�S�nf5��dp!8���@!-��o��\姉�����}�rڨݥ/r���#"C���` X}B�4��۽ׁq�g��k�'���tRG&�L4��A�1��>l�5<Ʃ������JlG��R>z�J���>����9�.��O�Ի�G :�Go�	���7�9 t�1�� mg����90dsL��Ӕ�<�Q�+�tI�7id���j��7X'x����2,#���"�
;V�I��� ����D	F�D�R���8���>���w-�KJU��� ��� �ڲtÉ���_��w'&^$<�l4���(��1!�/�Sg2RM�t�o�ш��v��Hl��M��8�\���ɽ��
�V~$�
��'���ǝ��ͼ���R%�ܡpQ0�TjE���@l�:�x\d�I�8��G�������P�0����>�����Y��J9("|,k]��b�������5�~� =��e�Cٱ	o��U��Mh��ފM�n��[���c%���́w�p�����:��/+�J�����5��V셊F�~������Ǆ��'/��]֭a���)�p8���D�L��(�åT�馩7S�%!�0]C�{����<? ����8vI"�� 	�׷�^�i��4B+�t��J�;����_4���{�i��ɷ�t��ٴ��[��)�[�=�����d5��`�zj�r��-�?�ќ^�f�u���fɧ��_X�/֜0�Ք��0��dՙuڞ$�v:_����^KO���y��X�H1쭲�T�Tmk5��7��v�^t=4��F,��,�GڇbaE+W�	��^�N��'n3�s0w��pI�?��3�FV&'���1yh��"?�V&k��rMĦ���#�����諸M��:���:B���s���N�=tX��-�h)�d�6�?�����{�6D�zꐘ^Yp�t(�����(�h���0���3Y�e:S���9�}��1_C)�׻����@�� ����ն	g�O��@ͦD�ϢC�pTB!f�u��v�]�����WsU]�KI�Sr��_r���j�����/��/�;x��.<��HȑB��6��M�G�5��C���/�Fd詴�c�������!��vH��XW����1T�B���g���d���LJ��+���h��̻fL�&펼���h��Y�M�6�'�B�Ht(D�ONK����5<�L���2�ߧ�J�,Lnq���5�c%�7����w����ۧ �����\�"��@�h�����s�y�K/�ӽ��!���,�m�f�[���o��t�g���\��޸��"c�0ۑ������dՓ0�������W�Qj��ҿ�j�Gg���܉����v�0�f~���:@���N��@Jo;�����.�{,��l�Pc�`�M7m02BH�]�c��?N��VK�)E9#���*���@���\W����"�CJ��:*�Vұ�r���W�lm2��:�рt�EL�"Mn����l�k�KSA�DIؼ��Y�:�6W0��g\͏0����q���l�PV�$��i0����;s2� �����a�f��<��?�G ��4AށK�U��lG�]�e߿.�*i�p�Y'}A =^���R��аV�d_N�<���h<)�����U�8�(*bU������K3�'[�V�kF۝.�=!_�B�(�б0Ճ4���*����a���O53����U��iN�iS�*�e��e���~5E���������bn�C��!��)��4�T]�>�;km���(#��Zs�ExøZ��3DqÔ,7�A"�9�������ۓhe196�J�2�,8�)���$e���P���>ʸ����[M?�E%�/y����=�����d�3(��.Ӳ�!K(!H$C� ��|ޕ0f!UgTF�5�|FRU��gD�O��u�/�Yڼ��ť���'i��r�#���=n�,M	I��k���m#���?d�-�Ό)�o��đ+-���f��}��M��*��c�<6r�o�{�6�	R�	M��u����o�DE�ˤ<`p0SP�H��{����S�q3X@1g�pQK_��_�?x,�#_����k(5�e�O)��h��z�ϴ 6���16���ʛQm��7r&e�K����>fe/G�6r,R'���c��*ѺnĄ�t�Q�1.K�A��\V�b3`+����74��K�T���Z
g����<va"�~X%���������%�QOqs[��x<�gc�������� ��q]�ջ0��|6K�w�������

�hm ��;�v��P*jk�������Yg7ځ������K�p<�E�)�bJ=j�CF��5�(�é�Տ�6�M�1^����I��Q�@a�P���G���b�-�_r=Z5l����~��Kd̡���{G�o2tBŝ���A ̉�� ��]&�Z��j�C��&��:h�6 �����OW��lf��%V���rȓ��n"�hՅ �uj_���}����iPl��t�(��I�I A�7$�j��Ӧq`0
�x�ho�{�����o�_��L%/Z$h�=k�^�)�=Y�ｳYX�Pز޴lf�zFÔ�
�XV;R�s<ȡٱ���JIx�w쑘��h��V*cVv]�8����a��x�y:��W�G%[��O�=�p��ME9睸����O8R�Ѫ����jL�)��A�tO�D�V�nf��&�{��y�1��Xť7��%����Ҳ����PW�t)G�l-�·������M=�I�'�g�+^N��$�lP9�������LfS�8� ��.u���e��׃��	�ͅ�<Ln� gg̊{����:N9s��s+���QT���ҁQ�Q5=s����1nT�B |2��7�F�;L*�_�����c��B��ƀП�a��ZkX������KV..�x�KD�9S{IW[��W|r{4`C��^q������)<�ũV_�I�c)��h#bM�Ԣ5+�-#ɵ
��+&>�Ă�xv��H<.�"��L�i��ؾxWd}1	�A�J��16ֹR)Z������IO�%(0����]���"�B����Or�@ubSQBt��[�~�ћ��H��1rV���0Ou���55L�+_i�������~�o�OdX<��s[�n���ʗޢ���]�4�P��`��#����o�PN�g�na}\wp�E{�]��,Dl�FK�gq&p58��.1�VM3�)��3��x��|�Q����A[5B������>	x����!�8�K���t����8�7Ѱ
=��)�~8k���b�^���!:������b#�٥9'�"��uLSУ��z����[� ��}�[��u��4��%C�1QJ����?�S�\�����:����ǼnwPF�����{���G�;ɧ����:���5��2�k��U�Z�t �0�-�A��v�A��t�������0�5Η�ļ�+���4�t�xOE"���P�S+��
�^y�+,�����_ܳ���P���^YmoU�_����e��i����׋e�~�NGҝ�V�k`E�2�D�m
Ù��3�[6g���%��Sx��[��fz�Op��-�z���3��M����B��� �4��-�I�� �����&�g�n�-U|�*���AV�h��Uy�X�A���wo��rC�~H�4��K�7��ȧ���v�z1��PZ���c����1<®K�-0pSF��1���f[��4D�&���-xE�.��&���.c�1@�$v :"V�Nj�ç��/�y�Mm�,���ۀEk���ш�p��E�Y����,vB��}6Ҕ|�7����\КNw����x����� �o�?$(󟺵��,u*��B�8�5b፬�\���H��P�-#C���a�
?��x�	a�P!�mMK"��+W"Fs���n�Ļ�����ǚ�0.n���D��D.����/,���F���ns�0D?�kc�&�iO\��VA�	�3�7פډ��g������M���k�����&t[��}_���.�cH�Kd�o���-�q������#�m��F��{|�e�tYV�5��TF��Z ��Z���x�*֐Xw�ƞ�R���3�5��)ט�h?�)�0ԯ���75ӊ ƚ��a?�I0O���A���[;�ԛ�ki��㎗�|�Ŧ~�2��j�V͝d�`�U�pa�!��QbM�����q�,�ZQja�����d���2겖�sF��bl̆c��Vee�/^U��)�b��1�q:��u�h�5$,*�8���ӺE��2��sY�G��ѣƠ^pH<A�� >ۊi>�Mɨ��loE5�mU�hJT�V�y���czF��(`y�m6���z9�3#�#/��(��*NXڌ�t=���ƶӯ�g�0HH GqC�LV�{�Zp%#�:x!Vy�?�����R���QY�jrf&Ŵ=���"�\b7'�?B�7���ľ� �Y���{��\Yk,��D;���@h�����xo�`04��Vz �_+Ov-��j�LQ�L`�#U<�E-^
�3���?}&��Ҫw�����X:�]���g��F�拵��%!S��A#�Uf�w5V��B�> �z���� F�,z�dS��Y���#O��O�x*T�6@0��#m���x��)��q�E�iB��Xp���9z�t�t9�&D���x>T�L!��8	]�?8��Y�a�4�Z�Dqe%���4�Ѧ�%��M*�}ڼ২����Y���if�h��_Hu��z��謓UB�e��I42���/��P� #/m���,,s�'꼧�x��c-ѯ�i��t�܉��d�m̶Pg+��9�����ts`��y5�����ѝ�;^�����u� ��#��g2��
F��<#��s�p(gmi1��^U(����Q��h��-���P��<C�6$�i�ڡ0KS�V�{��~�1�<�d�8cb$�?�Oy�9g�%HR�b��ںM�ޥ�����o��X�k�8�S�bڎ�*9�b+���ّ�{;1<|/����_�9�2�|ʈ�w|g��`X<�6u���@����P��w��?�H�.x�ѩ�T����h�ő����5�|6G2zFr�p�ld�E�&�xY�-���}�MC�k>=f���ѣk:�}ҕ1ٌ�����7;���PY�L����ط�H�	�0qʤ�S���HD�|����d�nC@�Cy@�m1U����<w�*IUv�$RI�<��m'��q�O-<ڞM��S����� �JX��{�D�_��Q�2Y]�{Xk��]���.���B��e��h��>��m�Ю���ع�.�+,0>u�=�{1�ѓ�_�-��6���G���0��%�'wQ�e�Ƨ)z�������(u������,A��ж��E����E�'���W����B��&�ĳ�]� -_�Bg�
�x֪��qÌ��_��E�i�w�й�*
I�+����%����|��1�w�Q�`O�$���/5��X&�v\ɞ]5�,g?7�g(��]N�����ٲǳ}Jp�]?)Q�ױY0�s[��ަY��B|[y�@j�~M���"؁
A2��D�>��?c�s	q .�P�B.;嚆����ͅ�����x ��/ ٨RZ�J-z7�C3z'��C��K�F�
!o0�*��:��R�մ�>|�W
��w�A�S�ß������$9�`� ��P���7|P�k)h(�2Ⱥy׽�̊C��-�bc�B�Ա߈�Qf֬uS���*
H��s�B���I�Vd�����\iŨ�E{)��mf����QU~�s�܀�Qw*�F�Q����̮��Im���g��c-7�3D��|�1{���j��I^ES��1)�Z�$%f+�%(��]pH�s�`�x
��NCl�ǜ�"�vT�/�ᑠ�_ێ�C�ŚIW��&�W�?�f9�,�@�6�M��U��ׂ�b������
�,�����϶4�ͽ~�r�.N��������4�g#gVITH>�~��^%c;!�CU�h=���%�&@��w�'�*�Eݳ���Ȱy/-�^��X0wd�%e�,=_���>x5��ң��DJ�3�M54hS�h���QF��w6SI$bG������D3�!Hȁy�br�~��n3���<g��R2�?&��v	�_��K�_��r����$���e�Yr%� !��z���s//,�E}��ʮ�e$�d즈��Wԃ\��B%fJ!�GpF�݈6��Ƃ��O�!��x~��H�2W��%�{����,�%�F�� ��)��s���^�C\��}�TQ��`3O��/G)|��d	O��Y�^ȔDsa86"� Lɖ
X���G��0���PE�z�Ћ\�C-]k�g����u�N���E��R���Ι	�G�$�_`k����MƝ��Z��,��!�L�2/|
l�}���G����ԬH���:+��ƃ�>�-�'��: h�N��x�4k#?��ٲ��~*UKz�W.jN�H��/���pnh_,�b��wɽ��l��)��n�TwL��2,Z�ջ�
	��0J菁(�Ƅ�E
�����*�'�3�%I �n�1d.?�N�� >��������:!�W�Z�����C�M�.�{)� 6]:	���0���(�2�s{�f��l)<��i�*̇������5u5/��~�=O
�΃��6���{\8ܲ�8�9<j{��8���J�2dYC$K:�0��C!a����mt��d�*��.���^�t3�ސ�{�KC�P�Q�.���!�5#fk��S�&D`��OƃV�p����Oy���<�|k�,�IEU��J�����^RH� �Jq)���t#��+�������T��'VM&����-�i�̴2������S��.���1lf�0�hR6�Fv���.f�#u�72�&o�!z���&��e�s�'����y�4?�}y� ��vu3�	�`f�Y�R:(ޜ�U^�NS�D�p�^�rl� j�����~��u�W��	���}�iA���0��ǳ�4T��([�O��������+P��(���X�(��w��n�G���N%��*����]����[f��֜^hW���
2�p�� �/����%���m=l��*�W����R��*�|��:Ȥ'ldNf����˦jot �.�ךѯ&z�x���f�
t��߽��B3�!dK^<(���e0xJT;DE����{m�+C9�wC�����	q��D0qaw2���_����3����R�`�`��U�����r:�Y��O�^*�+c^��J���_e�l0������"��{l�/�:2�� ��!@�?��Z�\�,25NK��A���dj���Q����ר�w����S�Ɓ=���=���	#5L�r�a��l��*�Qy@,��|��y<S�D�S�Qy�'��m�DOi!�zK3�حVCðd���"_�m��d��� �5���x�19��B�즷X�%�A"ET�1`a#�}��-���$D��wH���/���,jBq�c�{��_|���̰�#�ת^v��H\��,�H�P3d*���/.I����^��
�W͵���/�$���F"�q:`n�6�&��홏m���v���L�&D��un͒�$-8�T���(�Ƞj�G��#{����$r���Dj,��9z��������5?���e�.v�^#W�WN��]iaj����^gr���{�M_k*�����I��E�t�t�K��DOw����4Ŏ#a���_ֻ�T��i��"��m��o��܌��R�����I�R\m��R�=]b�()�`п��e�&F*Ѿs�S<5vH��&��S�����ٞ�u�F���R(H�U�!5��Da���&�6�e�V�Nd�II�Q55�'�@�c����~�Ъ| I���Z��pU��wfs��l�o�|s�-�r�U(Ʊ�U�ܞ�uGZY��m��Ώ��b��t$F(�7�,P��S�3c��������Q��	�`�E�tv%����N�q��r�8�sү�9+ͯN
Z9�v�T��C��m�ׄ��Sʯ�z��/� @�JBN�UX5C�V.��slz�;!S~+�)J�����Z�Z�Y:�]�I��!�Wz�:�&e<G1��*=|��\Kb�r�k�4D�9�w�ײں��xi��]�炧Gʺ���"����`\��2�IҖǊ$&asL%�}���a>;p ���e��P�r=`�-��=�l�Uvk�H��b2,c*�����?d|���CTJ�hED�#�/�WK�<��ܚ4#Y�B#EU8l��r~��<s��ku�p�V^�8D�+ �����s���)�,]q�Y�z����pżA��j�f��hB*A�a1E�e��β��`�o�qĐ�羡�i7�=ц�[��6O�)��I� 'F�w�Έ�ɯ���d�"*^�k��#��r��50�".�V�֭���s\��fSt f����8���Y�AƃK����_���s%7c� `z�nup<#�����y�����Hձ��&=]��-��.��	����j�,mZ0�^�8��,�"�eC�u�NG��]�8��T1b"Q|�ZD��SL�=fz튶�~~�ĭL�%~PA뿀���<�p/����_�-�����$�G=~�|�*'������rz���%Q7_�T���^Gj�7Z��ɩL�QG��n	���	�tҩ˛R�^�+��D�M0�J̨ܳI6���� ��̵�����؈
S1�*����a���e��1(����.�9�"�Sf���b����
�rd��'FUOտ�Ԉ\���� pT�<�wk@��n?�^�D��EưU�ھK��5Y��}[˒�D��2W��=�8�
A�8
�Q��Ε7c��\����졼ׁ7�;��}x�B�y\{�a�ڛ.���pS f��xrY �q�w�;iX,۬7�;V0�4p?R�@?�fNGG�b}�^1b::e�1*��0��6��ݕH2S
���#���29���g#��TP�qb�ȯ단'����s�S�ho9��[S��l�/�/8��񭆖`���A���f��m�$~�|�:��S�1�s�Nx��~@���3�ڞ1H�#��Cr��xU��/n�#���@Ԩ���	7q�uv)<K�٘��K�'��{���G+�{���g�*h�j���;1\�Xr���UD4΄M�`�{�v�t_�v�S����k+q��`��H�Xa@ѢR�u��)�Mr���[��5��9p�L��J>�i�����%�4|z�Z���C8�F�� �E*�����7���j���������v�*���`Ыvn+8��/��@$��M@���ni�r|�=�B�)�O�W��6����(.�ɐ�T�"�~���� ��LRdx%�T����gV�}��+!������N�f\��R�U}y����c~��,k,pcߚl=�O�%%jq��f���"&�����������D��v}�y<��Kgg��~�/�Hq�	�NQ�����D�������nԒJ���&�ݧ1�6���ɛ��D���ߵ��]Q??�5��@��G�}_�»���rոP�?��
�&�"Dl_��o<ʒ�:�,#����X�a���c�wK���k�|kyً�/g�������ں�pY��S&=x�3+��3�O�A������BMO�A�1����)`C:zb_M����Dd�%�9�`�e��[	�q+�6�t��z ���&��f��(�ԏ|��^_�Vҗ��* l��*^�jha��i����Q�p�f��_�%��v ���XN��W�� !ѧ�u�Q�Ȟb0~~P ��B��3(���|q۷}bI�j��;lώ?�%2/��z�*%9��G�bއ�5�_�����Y���^�����(܏x����v#����J�z��.��x�hm�Ac��;�X*i�;���z�ʱ�څ��=h�9������.A��V3���)�G(�� ������rŨi�i��pW{�3���*|$i�9#�mº( ��\U�c$��pA�`j�A��?Z��v����$�1����*�����pPc�x�� T�Mp@��)��=]c鈓,�����E?���X2I�;#P�6��V�D��3HV��kB��A(����Ƒ��+$�f�1��������®=q6�<�a�D�ӫ��
b�M�7��4P�zٲbA;~Gn0�����^��*S�P5��M�����#5����6h#�*5�m�=�����&�Ʋ����Q��~ږ���E�o ��~LH[�sL,y�G7>�vΐ���&ҕ��L�������Q��!� .>h�A�7���(��pX�m�@2��y��KO~+�u-*˗kF7̺J_+�&��(SC!ٰ��V��fx�҇����A��,%���/P�VB|OJҴ�r��u�?�u�zHBwj�a��t��1j�hkPd���%�me^/2��Q���2�3	F�Ԍqd,���q�N�� ��5�M�L��G����@��K�p���jW&�?=�?j8H�滯��0�8�����s ��T�͓��j�ȍ�'	2��{䮧��^bm�KWl"w:�+o
�+d�`E^�Ž��Z"҆�M����)�cn��&ɡ�n��hu�TL��x�V�ԾF��^j�c�9��&!/h2]��g����)��G��jd��JT����NK�9#���L� ��5�Ώ�iZ��R`���7���юoa���>S�����S�_��_&�j^����󼁪 Đ+��u;ks���\����^6cݬ9U�����+Q#�7%S����g�e�3�n�r;%���@�5*�O�8 ��\[��#q]J�9���Z��0��9_D=!�8��EO�����;�ƀ�0��b�`�2h
錐�L쨑b&�Z���UW����`2��Yn�z1������~��}&V����ENlH7���N�ˤ������kLxq��\0� �L�;/X���'f`?(�ߟ,R��΃�K�c<k�e���uNު4v1Q��"#~��u��-@��X��;7�yS@ m��0�01&�����8��m�n<eN-��uX�`��A �9�4g1�=ˋ�9 Ά�~^��]�Yp����E�&㊠��6��ɼ������9���e�Ȥ}��?��;�f�$����ѰK	��qt0� �\�*�O	T��=f:Z��,��(D.r�b�u{��=��}��ɖ�s�G�:��-�/R�E��RQ�5�#L�v{r���I��Nd��h� ����4��p$���T�xj\[�ךZ���پ-cu�mOԭ�R�w�,�cE�6.K��\�*o�o�gO`c�	��DO,"�$+8��@�5�ýj2`�����z~M��'�%��O�#�Pi@���aa~�ؖ��*�-S�_XY����U�Je���ŗ��n]�=m�yl�6?�k�N
�����`�;E��Hx���?�{ ~��q�RY�����RP�F$1��]�/h�jf�ͧj��!�ҫ�E�E���G/�r��$��k�eK� ^,%���fW�,ì�����&h��&g�7�ψs'Z*�<�.�MHf�y�{��|�ᘈ�31{��SmwY~�';��yP�ڝ��zA�S���;�;%ܬ��|�,jP{�{# �M���nGȣ�E��)g$4��ݠI�%5%��Ȅ��޸��_[�(��}\���C��D��%�T�Y����s ���=P�|-�U���1��4 �{%oyZ�6I����3���htn�g8{���9h��S:͵�;F_ͻ���+Ϯ�<�����v0K��J��+��Jʺd�L]����2Z�����~2�o��=���D�0��V.�E�Z9�C%�E�������Q�Nчy����Xã����0֌�V��ȼ��:X�Z�QL�U�, 5�*"'D���$B[q=�d���c,���Z:�h1P|Ѧ���c�(0ք���͌�̖{ Zδ#��t-�!�q��Y+�)M�C��xv���}]���$�F�r;���������8g�����z
��tD�3gӢ���D�>��h�v}�N��3Z�<}W>02���)9��k�_˜�̢|>��Щ%7wz�����Dn�(1�%��,���@{��&v�U��FQxE-�l�4?�|.[+a'��^����q��-�|�Jɩ@�Q�N�HR+�Ց��U�y��%a{Z��|A����C�gZ�F�̻��a���z��ٿ�]M�$���7ѐ�����^�b��V�.�Ʌ�o���O�PJ����>����n~.m��-�V5���ub�n���F�.�`@}{Q)�u�p���Eܠds|C���8V�a�
�]z��t�w�c`��ߐ�:�"��^gC�=��q.pxӎ+6y��ʒ�(I�S3�r	txa�(&{$ÓƸ�;Y�����!��QF$�
U���gM��6n/�}Y2p�W���n�4�ӫ`sL���%���a��zR �B�я�j�da{���.���Q6�����_��Y�u4\S OFܭ��RE�TE�Ą��$�"8��sE'J�}�$0G��ݭ�n4R�9�{�f'T��^P-�|���_ �%�!Am�p���W~.�\�B��d��ɺ!�����ߞe.��zèJp*aD0�<5ߛ��ŘU��6x�=�2K!�X��xw���/�l��&g����6-�m���cYE)b�.6͞V�)�@DA��� �,e��>f��F��:��Lg�[�Ħ���D��k���h����,${ٻ�Y�ſ 2zd��{6�4��=�V���f�I�J3��zkyO��\�ޡt����k���Muڤ���_�p�~��Q�v��T���~H�InRYg�@^䙋:ʈ���C��}�6g�tʀo����N��UlV�m!Kĉ���.]�w>����d��ø�Md�axZ$�E9#��Co�K��z�[_��'�y��'�7fh��Ѻ��k���i_�u�ʿ
G<����R�|���+y\��k��|ǡ<��G���i��N���R�u�<)󱏃�2(bN��C�N"�B��[��K4(����V1r������U	Ҹ��V����Y}K I�/�6��av)�D�Yp	4�,�u ;u-�����P�o��:)����S�t�F�;"�K��
�A�����'2#"
D�(���[F���y��,`�/���E��1�u�e��T˱Z�à�"���D��L4��3 4�Ho&E����(L+�sO����e��"��� p�r���I�S��_)Lo���S$�R����Vσ_����X�$(x�������-U���'mL/��y��)�I���-�F�P��z'W�G�}H^���Ϛ�-đ���O�D�-�\��
�b��JRd�d��~k��m3�}`oI]0�kv-�`1.�kR�DX��z��+�W�� 'k��;��������j��ē	x��S��<sy�(���ĉ��.��Y�P&��EMC��1���G����!�fh_'�R��$l�|夼�׋24����
i��S�{81��N�V�D%�΄G['W.�m��XIV�z*皐�V#�$�=��Q_t�`��y��4׬+�J4㖧+����7�@$&쎀�k�9<n�S-�K�@�W;�X��|�C�/#��~��>����5
- <)�J�����7;j�͙�Bt�d��9I���!B�z�,i��ҳr�x���ebD�njS�T�T����Y`x2LD��lv6��~��_��|S/I�ƥ '�ꋧ�/H+v]�[M�jv���=|d;	��ǉc��k`0�ќ�N�M�����ly�D�V���2�t��Y�cmK�I0���z���X.����"���e��mu��]e��..ݻ�`�A��ˎ8F
Ns�ԯ~34w��a��\U�oL��ќw�Z�)��� ���uN���:�о����!�tdQ#����<d�gzOl�܃�l��'�15�����[J�ݡN�=��L�1򘢓y�Խ�ý�wĎ��(�+"�乱�T��D,�eP׶uf�
4vǳ��/D�Ϙ"ɾ��I?�8(�WV�kਪ�K�9� ��k`����L�n1#���eJlO:&�����^g,<r�� ++���
�pڀ��!y��t�<k����V���69�F>�����M����U�0$j��C���ef��@�<Q�l3��(�ƽ',�z���f�2\�3�����;K�W�G�4"WGX����b��D�cK���>X���-��
��iK���'�LiC����w�a���5җ}��Sr�C���K�~��*�s734�d�SMg�E�1TtIy�O�%!|�P�+1f��V����%T�O�7D�86����;&wg12M�M�����'+�����,�Bpȿt*�L5k�1e{	�n}����S�Z�Kӧ|;�{�ͣ�9j���\�t�W�Ji�1I9u��-��l"IkN����ȿ|��U���������:v�F/���G������B"�i� #}G� �,�������鏹�1���BU�b;҇�j��Qj�Jڿ��L@{�aX>�����\*)&f��	��9�r���Ǟ#wFOE%�Ky�� �Hy5�5`�
+�����A�H�jԮ�����K͝_JP�t�M�e�\Y~阈��'�,���=�M���9��KHA���?B�l�ڳ�%���֗��C�Fq|03p�2]��Rpلr�����	v!��5Ї�~EK~[���\þ΄Wʖ]�[�]��7�,��ᚊ�d�&��GX���ĕd�<�g�}���n�q2�$.�N��F��]��	8h�v>ΤL(��`F)d���qY��b�C�g����*�H��v�0�`8�@�(ef��|��7��}��*��X���,k9�h�9!�\���;Q]�2�+�1T������T������b�F$��Ӗ������|}rn��N�V����c���L�Fe�O�J{�����[���PP�ʟ��zX���~T�H�&��gd�|���SR
�d�����h�� ����]����&���eSnI\�#��S��N8�Bw�z~Q�QnNf��ɱ�O*���X�Z�u&��� �F�:#
�B��/?�sa'���1<bYk.��<5$���ѽ�Ϳ��]$��E�?��A�u�HR���5�K6B��`ٸ�B:nb���~7+Q��m]�X�*�����Uk�*@��)��i~���,'���$��b�Y�7��`�w��;� {1Li}���9	���������
]��zW=�������Q���럥�L�c^}����ܟ�%�[��9Ju��V�z)���P�2�A~ۋ�8���GO��
{�䈼>�=c:B�MU��;ÚxN2R6����@l0�����{-;��@Ҵ�G;/� �����u��;��f{	]x�5�/�&�P9'@��g��O���逭Aq$�*	��T��A�ur�X�^#K����V�/�)�w����}�UO���\���ɯGbb>��4�c2d�ӊ<\0�Wq&>�՚������a�v�-p�Y"�ѳ n�#�C��O+�]��[n���vSY<D�A������d�V�4�-s��D��8*�q��{��n�w��?���+d��n��c�DC�#N��&���v�M[���:�nٙ7��OJ�T�����o�PQ����ΰB�H`	Y����T�Ýe�I�&(�>9�[Qw�u�t�6�7YK�i@��9�B�efwφ�D�mѩ��?���;b�G'� �6��p���Y��(��|.����A���%�f��@�x��L��a�x �n~5گ|�o�3���e�oy ��.W`�7N)�������oRq��q>$�,�kx�J�K��>4R��2a��^Ŧ��7~�y�������������N
@cP��J���Qm��s���q�aڳ[��m�j�PF� �ƻ 	ہ��q��b7ri6�%�[/� ��3�Y|!1��x�����%��һf��r�qGQ.��tO�@�Q�mG��M1��{ta�v���}��&����x�Bb���	 �~P����U* `�̔�S��j#�ө��Q��%�P��v�s�%��Qg)!r/��OJ�
�F�T�ߗ�X�<�RxfE�+M�t�ד%��v��d$��&Z1A�t��N�����Y��֮[�B�s�oi���ah��{�sm(0�,ti[�ec�J�uP��e�&4�iN���d��KY�v�+G���L��{��J�+(�[а� �J$[T��6���F��+*:~���BB��? ]d�V�[w�.�Lbi� �-6#��_!����xB�ޜo~a���A����IR�C��W�Өԇ .ĵ=�A��Ȓ	�N�2k�>�.�`��`#;L�G�����d$T5LUx�����3�נ5�g�}%Ktz�a;� �����?��)�t�����v21�oO�ex��6��}.���bxAf����B�}���ϖ�A���N/����赌[�Z/�f`H) ���i��I���5a�Ӏ�b�F���?q�����u>%��@���݆�ZE���iL����� �#5�-�9�Q��*f�ub��Nt���@�@�Id �p��	���E��@�r�W���dǧ�K5��*0�ik݅��u��j�E�z"�q�]-wSD��+ܾ5N��������$>	X�
r����x�`�V�j��ʁ�M�݋ Sc#@\h7�<�2��l|�d�Ӑ؀�{2�JY�����,������������6�Z��n��^��e�U2'� ��!��0�ܲ>\x!��8����";��i�#!���sՃt2=����f|/�u,��-a(~�(+R�{������ /�􉂢) �d/���	5Vr��;Yͧh��b�ID�/��&���@m����r3��p,(�`{���F�z�����a��n�{����w�O��z�-�1'}+f^ ���T��[3������_��(��z�����,m�T�qܣa��7&��)mBJ� �'��W=�ζ�/W�;}!�m���_IBʬփ/��
yq|#]��0;�
|Z��v�5Z��{��lt���AIWv�=U�p�	�g&EȨ�����O-D3a��a$�Y�c8�;�?��LPyԓ��Z������qf�}��m,��3U���N��3�'AT�nƤ� ��'��� s풭����p;0\a�����׿f��(�W��&mQ�i9P�G�Co�\��-�ĽF|�m�{z��E���uu>1�]�YIb����u7��{�1�:2_"��e���<��m��U�T��V�$��R���t,�Sc�>ƶ�+�"��g���|^4O6�kA�V���4���o}!�}Aᕍؽ�C]v@Ջ0����#��s{)7�����U ���K��Z����I�s���Ծ��4��+�&ۼXz8��� q,>��Zo љ�œZ��6�O&��OsO���\?FB����"0M�0�b����n�N+X&Pq
�kf�.�Ʈ �\�Ά��u4]�<���a�7V�wľ�&
jP�$/�����#��}���گ7�ğ�d��U�<����,o�х�mHo�Oy *09CU�3d�rq�\{G�3�Q`%8Rq]��E¸�z�;�WO��4��-zv*�dJ��:�g~�vɟ� [�ʲ�z��OKI�Cˮ��P�&9�����ؠ��}Z�����I|*P�ς�������d���"}�@SsM^s`��*��h�+�������:�q�J�BG� ��Q\#M�0��?��ܱ�t�)b�@�N$��e���j���wr��4͑Q�� ���&i#  m�ӽj>�k��y�ԅ���o3|�iPM������Ƽ9�����u{4I��W�
z���tKꬵKg�5/��1�
Iq��M7�=!��"�$�f�I�1�pl|&�V)��>k1س�I׭ ��` �\��v�O�������(�֕#5Y\��Ơ�\����2j��Q�>�q�l��>������Y�(r�[0����70c��͈�~Ƅ�H'f#T��:��g���p���i���
�J�mO��31�fҷ��b�*V�/�����#>ט�׌�]-� K2m��]u-h�.
>r7��-�I�7ǔ���?��y;&�=u��n����CC�ĝԲ����[GJT�M�g�9�
�W��V�5a�k.QA��FŸ���O��ff7%�y{�҄iT�x�{
�`e�snnr�������?`%���5��rA��5��J_y`����S�NzW�)7+�^���B�fP�(�W��l�[�x��$�H]3�����r��u#gw�<������:��Y���[��M�ǂ�En�k� /Qث���y8�m�h�w���yt��Qj����\�1�H�]�D��c��@F=�*+j�4��U��v��SL5� x���k�0��:;W0���3�.��Ki+�צ��~����'"hU)���.Cуj�za�n�?]�6�2��X�v I�Ì��[�/;M�6F�ӄ��C��ǠD��L���F�%��\?�jt^j�`���(Y���;n�p������讗6'\ln�#�N�3�|Dk�GJ�=�uҡ��*�ʍ6=���=��tnxaɚ��uY�!��{���R*et �O��C/\��L�S��2+��0z�r��#ܣ��EVf��0�.��G�L��9����|r�)�6<�|G&�H0X�8����s�*H��a�%֙��g�E2ӌ ��KԢ���������<	��z�s6����_�s>�&On7�a!H�S[_td~��ye��1��5�E��ƴA�� ͣ�uW����ۻ>᜚L!�*�j��j�9޸�¼)�xAܑ���.�d��/&0q����Q�P���t�h)tgDg#�ݸ�����&{@I�01�G���up�p���pO�R��⍿Y4D+3I�y\����2W�^n|�xַ��(ڿGLV�t?��xm�/%�Ey���SW5��������/� ?�4=CMk��k�.F�Ї�<��l.	���R�k1Nͬ.�(X��d[զ��3f4<��0����(&�����e���b��7<TpI�Z#/}���@)�މ�O-��n��ː�K�v��o��!�P	^�r�Q%�����q��:'b���,�L��{q!g��{����W6��NL]�Z�E�e2��I��ܴ.y/�������κh
Z��kn��,���Vz���H@Ba*��a��'wu�scs�X6��l{ ��9���t���~=7"���H�±�GT?ι�ҫ����^��+Z��4?w
��R��e�!8�,f���]W ڡ1�3iDΓ�>~�1����^�Ӥ�i�����v��3���,$|����z��4'���l��(�@�z�	1�7�B�5���3����t�=W��V��|&/7[��N?�6�(��M�J�U��U1 j�&�OR��}����dJ2K��of�!���S��Ҡ:'+�(XҶ��,����s� �sv����AZ��ڄ"�&:؃Nڬ���������-8� �%מH��!������o��(�oIr�2d9��M��f���g�匀��Ofr���sY�v�����30��@�v����qgR�J��\�{�]rL�q����cF��BD�P�t��C�۸9���9Ƚ���ʮ��h��\R5����0���W�Lfj�]60�=6�R�P���z&�e���V���(��S��6�.y�]��qB�ve&��\&*�k��[�#C��QwXo�xLϢ ���s�hG ás��%�1z�d�"2�^��1�;�\���!�X3gx��V�x�{`�c~�r<��V�͹���4�ZT�?i�♭Ŗ������S����5�K���Z��R,�A�i����Β�X���	�.��W9�\I>
�o2��~�-Z�^�l��\2������v܂xK�K��=L�+K�=M�h�K�������R5�Q�dzE��f�&��d�պU��4tH��+<���f2���۽��ƈou"����:q�)��	���)*�u��X��kM44�����ϗp��Ųr�p����Ef��c�}EP"�A
}eI���K�
[�9鹙����i�TF��C�*C}�B���_�P�Pq;=��-���Ӻ<�)`��wky�l�Q�;�>��2@L净���!Od�#��������L��嗵vv[O�mLU���^�/�H�6���txȿ�������)A�y��{h��L�ɇ}@
G�� Ӓ,��T����ʩt�c)R�(6��%���E�!خ%��6A ��;�Cd�%3��y��چWյ��h_ �*E�z���{<��9�@t���\Aٴ~���G�\r4�ԫ�}���~��S�B6�Aʳ �m�,$r1��@�C���0��<�	�i�W�n�J8�B�uK)x���M���Y��P��⅑j����g��b>Ґqԏ�#+���j�qW{y2�*��2�>��, 	~��jx3xT���e�˪`�=�#<��[�nb�NqUSÑV�3�p-�|��R�5:IC�j!I���@��ϖf�q_�e㯙��mc)�罋n���*{���-��2o��{q�O���pQ�UV������!�s}^���'����z�!K���������*#l�)�w&��ߞ������r�[}y_���iee��4i��N@&��%*eUp @�]PWs���Oo鯮�>4���o��p����q����͡`!L3E8�k�T������VK�l�g�C2�ʔP�"��O�L���k;^��S�a�k㯵���B�0�E�h�zoL���ȧD%7P|)k�bm�d��a�.����#�l@��m�K�!7Ǌ��o[�d�Gf�S�y����f���s����2h_j�5����4V����jcZ��h�,У�pK1A�X�����y�~	��]L��Ĵ��r�L����4��PfT�+F�p��n�о�����y?��'L��<��.�0e��QN��HW�%�b���@
��}�	5��f[�ѷr�i �c��C����J�F��n'}[�D��ꤦ)ʺjc��u�*��NaҴ�� ��r�������9*����B���,��.���^�l'�X�Tc��Z$GC6�<T�_��bӳ[^"��%���5Ǧ��S����My��g��@B��ִ+��ŮK]jRl�u��ӈa�q�"UГai��Z�v�����e�l�Z�Q,���5u��b��F�j^:;�:��&: �M4��ͿM�2U��	�ѱe�lY�OaVi]��de0�!Mט\�
���M��,�d����a ����J1$4"���{B��y��v�xB
f�4�%�0U���I��.�l�U�'t��������P�W�/�
]��A�xa%��,�h�th�@dzxҿ#��:����?��ڎ��,���!�:��DO�+w�J�<9(+�i�U��P�7�mr<�S�e6���;]��N�f�ȉ�v����P�� cCR�^P�B���M������XK����/
�J\=�i<g��O�� ��7z�z�]""�k��x
��oVĮ?F]�>�[��L٬������~r�"�O�n�����f�r���'d�>�hwR�:�W�'��) o��(��Oݓ�*H�a$�..�����I>��D�2�-o��x��qM�]��L,���(Hݢ�2�w�;��e�FP~���	��H�S:H�3�����*����1��ZW#G�9'��;����E.rz�&��v�@��24r�& �����t��Gbr��6n,Z�g���h��7	��p��o,u���*���Rf��C����Q�n�$���`a6-����.ؑ��6q��A�6�T���LH�:�9����O)_)��D��_������>�N�d$	�1c���C9����	e�t���2$Y�~�Y���T=p��\}ݟ+<���j:hH���#��r]�xj;�x� ,¡O��q8�l! Cɷ]l�^y���������GC�l)R�O:�1�+�$��s��M����~sO�7ߵ��:�,_�2=D˥]~�[�G������?��4ꄋ^�I���@cc�Ja�|בH�N���iGB�>Z��6؍'�*РY"��-W�4Y����������7��-��_�7_�S�]ؐ&�w�=�ҝO��d��Nhҝ�Y��F3Qh		�������G
tu��s�h8&C	qvU��K*!��jb�Z���u`L�m��������R�y��M��@��Vߓ�/�H�)�y�Pk���	[�FE�����(jj$���uq��Ҷ7*��0,�L��bJUl���V���pԳ7cF��QjrR�v #7� ÷r}�+7����ߝ�Q�v�6�m��:ob'���4ɜ���[���qX�!;�(5FW�0���M�~�.
G8;����f��� i�@f����A0�ٍ4Ѧ���	Yw`�_F���g%I&0m��Y�u}�%+��j�/�7l+�;���R�Po��-�
������/S���?����he���H(��״��/��s6U	d� }����tv�����o��W��󒿭ɚ� ��
\K�&N�B���*�+�`�U���\�w+x���/��Y�'�+V�*�)���/�u��*�Ɛ�����p�F����_\Z��<����1v�+^�V	����/.��o�U��h`��/c���^yo�sh��������kH�qޡR���M〘u3�`���ί��ʃ��j�<.��ʬ7T�F�I��T�Q��D��Q����!�[clt�|N�/΢e�49IW���)��.��׏Vt�Cu�]@�AhJ�"�D�7�"�-�����'�>�F�]���h��c�ex�,�!�{���d���KH�k����/��qh�����>]���!�oP0�!Y(X=(���
�n6J�V]=.(��"��\1���mzV��̜N<I��H��T,��,V�����+!bdӭh�dw� ��y�d���FNp"a����tUZM��D���CrP�ǰ��*}J�4�9�̭�0|���<"�{̢��0n˒f�p�b�5�iυp�*��0���cEW ��ߜ�h��>!��+��R�0(����`%lߞ<�%�3+
�5b!�JvV�Ȏ�<Wv�p^e�L_����>ْ���m��7�:г�h:P��J�y�P�nAu��`z����Ĵٌ%�@k����s�iu��2�Z�����ϩ�D_&kx����mS��<����vG*�Y�/�-�%k���r9V3����=�Ke�TA�Q�=P������	 �,V6��q����!��iH�T;�vJ-*t�-�Y��D8��Sۊ�9V�͕�*�U�Z!18L��Psw���K~��1T���a�%̩��w�ɐl�Ut��ǩS��M}cc�>�m!,�%�ʊ��'j��,3c[dmQ���<\H�V|�}���,r��R�3Ci����ٗ%I�m�iB���}��"遬g^��\6~�������:9+`C��G�KO�eғ���C1�'��X{�~�����27��� �^Ş搥M���ޖZ�c�ŕI�W/�
S� �{ ��[{��}Ô�껞35M��DC�(��ҧR��<栅&)n_}�0�yE�A廐ۘḊ����*/�c3E��K �n̟^�}h�u��BrP���������C�f3(�j[�?Q%[��=YY@�-��g�{!/&����C	0�R��G��p̞��n� �&�`�-�>������X5��_W���t�<L�s�|�@��LE|f'����Gr�+!nӘk�$��5 �w�60���m[�����6f���L��w0t�'�k=c��W�{J���5�|IwVJWM���P������8��/�m��)������ۉ�4�_m�U���|�S�AM�9�'>8s�n�m���%׊cʳ��] �乂ZB���ྔn�N흏��@��x���3��˝�U3GVD�W+�����8������(�~n��7컜�����=�.�a0[m��s{�j�~�j���1M�:��nW�]z��o��WP��7J��tꮵC�9\d�'r6ֻׯQAR��G��~W��
-rh��D5�1��������`l���<mØa��7��j(�G+�9f���CIkr�]��[D�P��4�T�4���=�K����ŷ�6�%�m)�I훻�{�{��4��d� ��@��| ��\�d�<8��JصK�}�U&L�U���.o��_]n?��Śۇ�fS��Y #9Z;�������BD�t������Z�ĂM��!�Kr��g�y��6����d�C(sQ+ $��ٔz��ּf��wA�[��۽�G%���(�K�$�������b�k�r�}���Rq3��i;LT
+^��Fi�lب�I`�&Ԑ�����+�J�'H�N�ؘ��p��p�U�t!L�~�K^�ÚD�eU�B�td�X���ǚS�1?�ju���|�⋘���ч8��4�%�7xC(�q2u�n�Ltó/�j���y�3	D�~�{>�xBY�t�Lq#�#I��`�.�q��y ��gXz����EeQ�r	�'|"�!e(�z�.
�-�F��p]�Sp b�G��4��p�����Q3)<N;�H���&��+.�SGU\�\˔����	��� �p������Q�c�r#L�'P��=�+b��t��耷�+"���$ķ͆�v������钻rvYDHL5nW���a��CY0���b#�^�DxN��J��y5\�d����~6���L�WZ�V����y_�B�<<C0J���@Ī	��C��!���n9�N۞n�Z� �zl�  ����SߌQ�c-?�Z���P�N��>�9��OL��R�
͢��2�0Z����l��~3m����v�������T���I��t�Y}����m΄�W�k+
��+��=�Rǎ�#b,�҂%9&�:���.#A{�]���!����ٰ��B���z�&�}��).�P�1e۟I���X�ҵ�@�z#6}s]&:���gR�7�_��4�8q{ �_Ai.�^)Pb%h�z���j���H@6e��
����?��痘XA�=�)�[�?�|�"'K����U �^�mϽ�Vy<�e̯����K������㦗�]<S�|1�ʳ�_{�������|����,�]�8����r��Q/�p�t�j�.�U��0�UW���)�86۫�pJ�7�$�5Q�a'�!��'`�LjJײ ���B��R�f%����)�ۻ����ʊ����d@��`�Z|���l��R�B�@^i�$�w�������/���}���������bԒ��H�%��gs.��l��?�+J�Z���o{W���j^�R��hsJ��01#�!0�\��5e���Tc�Ue"lɯ��62���=&(,�5b�IJ�-���bz����8��Ϙ���{�ŝ�e�<�&��/L.��k�ׁ�H]0��I��b�|�*ws�
J�n��]�T���R��'�4���0������Ij�-%1I�3h� �̚`/_DP�V�jH�'If���Nʁ5���瞐�|5*˧/�m�6�ږH]�Ŗ\9F�ࡠt�H�GZ8�	?^L�-�/����4H�HG!9Y��Ƃط����B����,�lG�Sa4�U���$B��?��*UO}������T�[���)��QAS��N�hm�6�Z0�""U�ǫ�+�(O�M����LȖ4��|@������HP�%羛���C�k��Dɛ�f����1X'W����t��;�J�����ʖ�u�˘/6���99EP��[� a{(V3k,�a�X�di��mt}�?Z�X3���<ի� �D�d��r:�L��+��ߍ-Uӹ~Z�D����̞�X&dh��n����r�`N��4�m��!�})�C����)�����}ʋ��htl���#یJ�Y�ݞ�9�p1T�&�UK�d����t�M|1?�}�,����p�6ng�|/��t�u��ڦ��^.��"�N��8�2�[!�4�jL�[�?��3�	��$�>���:�,A�A�$��XOk�ڿ�5��I~�����A�=a��;T�P��'�7�~�&p���0*����~�2Gp!���TҼ�����e�ws�<�ƒA	��h�U�b��n�ӎr��_�]���7�[b-�;���i�MVzl���(l˾�M*	a��q;ِY���Q��H����u����Ė��򠑆�%o:�36�����%�6
��ֽL�����ݛ�����vd��"��G�������A@��́�6$l��Rar����X@1���\�W�jO@��T��i�`W�o����=��IOpJ	��#G�rV�IQoV��Q8	�~P�}�h<��t��C6��$���<o��-b�`����%r�/�;[Ӆ!,��۟4�6�P/wKF�\�-N;��A�P6�5�y9B�$r�YÃ&
�q)]G�V)&k��X��{\�_���Q�f�FH!o��$�y ��?�E�:%�&!���y�&5���eG篊�w�Eo�3w����@F�" � ?���C�ew�O�7��z��KFv�G	��M;�ع+Î`�SR���n'�>aX�BJ��|�juT�W&���0X>KO��X�G��E��"��$��������q/��ZZ3C8��OmV�W�k"�(k���^"z:�Ǣ7��B��:����{Eҏ�vŅ�6�x�B����ྖ�i
�V���M���p�N�Vn���/����?.D�{���rLB ��ۗ2�Sge/M�DL�D[)�����H=��M�oKٙ���_l��݂�%��h��T��_j�/N��Ys��ES�q)(6>�Si4vPHΎ�f��%p����"�.2�;ԙ7�4�>�TaX��aV5�M�i'��@;�a��2?%���d��7���]��qO�q�ߺ�!��EA��oX5߂��e)��`�C��|3Y2�)��
�k@�t^qr~F��-�7���;�g,�k~���M�eh�	�>��A��SX�*���%*J^��ب�(3���`p�k�
uu��Z`LGzrP��K�6��B'�T���psp`�Z@v��:aU��BB�p���Ǆb���jJ��[��(�g��&!B�:v��?�2��?���FB��ߢ���q��e�	oY��V�;Qw�@�^Q�tGH'���*�I><���\�����;�q7I�ﵭ39���Y{x��<E3;{N�:A3�ՒSS��g�q<#S��n��&�k	E1ؠ�)-���j'��| ���VR���
S��H8�O�̐��F��j��f��3[���ܿ�zﮏʗZ���M��,S'�]h���c='H�>wET�Q��xY���.�?����� ?*<�y��A�t��=���t�*N$?y8cDx_X�c]h4^�R3@)���x0�e����Y}�[��$L�ѐ�<q��O�{"8�� �03���{�?�&T�U��C�/<]?p4�eM��4���.���hb����������4f�2������!����U�?l�v�x_�v����� 匝b�sPf0bI?�V�v���j���]`�^�l��BHԀ�����'%И��r_qa��3˸��)ыꥻ����0�3B�eMŅ!1x:��qk3�u���j�1�
��$���\?/��-1!F�9^z�`�u�����S0UV�+�����?.,�d��?1���A0�-�Lύ6-�"BR���NDO��'��yTݒ|��yx�xL�u%]��hHF�%��Хky���P6����O4�����߯����h�$�$]��$�ti����$��P��DN7�iߕB�a�.��<<8F���b�ի���xv"��y|gi�C�=�0�4��% ������]�3�Tb�J���\��7�UZG���qiAc�:ap�mp��Ͻ���{>�:���Մ�5�j�&w���e �o"��u��y�^����{��p���P ��r�od��ffb��/��k��lǥQ�%����|�5	��ʀ+I,��I�1�` c[^q�[�Oq�%:���kU�O�*T�����1<`�͸�uJ���@+� �Χ ��d�����R����7�	Ӎ�_P�:�6��B�Whk"�v��7R�<_ů�TR@�\�an�0�oΦ@�.*aR������Ϙi8b�5�����f�i���@m{�Z0.˪�M�>���˧�4����X��6)��������v6�("�̜�u�����Du5�9��C�p��$w�1N� ��ywl	\X+1#�N�6���qe57ȣP�X�W�#î;J��|�ٴ���'eܴL��zm�aF_b/$r�+��$p����Q�ϴ��G)�1$F�u_� ɹj9sn�^��5�V�^��E��s "}�����ڑ����A�z_���ىh)M�S��$a��`I�z�dM��m ����^�}2߆�$��r��Z~� ܊axt�+�1���8�"FA����|��|8M|����������տ���+w�#�]-O��s�`l���;��^0��v3V��~�A�s�R���xl�Ep��ry�����'I�_20
ƍ ��%%���GB�(� �<_�rLb�l[b&Ř0��A�;)K�L?���+`ݹ<�Y��J��h~��E�7�R�[��+ ��%:m{O6�
eYt�Å�<��q��+�/ǃ �&<j޷��y��w��W=oqL:���"�$�c���������"�e��u�~V�D�g��slU�|$�_��c��I/VBNY��I�&�u�&C�|4�9E����=����D`~;a3��w�z*��X��K_m���E��Iܪ�1�_C�7l�?�>���S?�(�k�ys�1��)��l�d�N��«dQ�����C�>���=��a��T뺀�&����BM��8�bܿ����������N���p>9�eQ�w6C/�w��21��Wp}������9�?x��]/�a�ׇb��������Y����D��W	���F}��{l&"�yr�̥i��<,�� ���#�̦��_�Ѯ�� �4�q=pp�l���p�(zrYG>R������S��LM�=�(�x�`<�`o4Η��d7#�,xBo<�ȯ��R��Fp����7ўs�AA�2�DTr}=	���W�`2B�Y�$q������'�t=N`_H��O=sk�`��`�7N�X߬���ӥ��K4C*�]��U�p�[�fd1��&��}@��������\�I�%�@6�g�\�WK���Y�o"ǀ�F`S�b�3D��T��,�}kOπ![��n��k���.g��������zS�r)+A��"�6ᆳ^��/�t�n7����t��` �H�Hn�g���m��h=^7�����/�S���8�N�.��/^�$o��O%�2�F�8¦������pEc\�%z���<7=a%��
m#��?�Lie�Rh��*rcy2���g*ť�w������[�ᗈuI��E(�%��ۖ��Kd��2R�^Q�ޭ����1���F,B�~:y��+{�7��E��v�m�.�B���dR�O^u�C�����
�k�Yz�@�Q9���=���8g�[�̠K�%Rp]o�}E{�tT䨕dB�=��v��$�W]�˴<*6�ք��K����L%�ţ�BX_��
�"
gX�yw*�dR9}d�bp��${��.�����K
6���RD�g�'�F}�d��ì�/$$�h3��7�%���qV�+{d�����v���o�~SW*�k�|{~jvMi�<,��z3�75ʼiڐ$���ż���y�-@��^�x��!]��0��Ri@xZ�'I�!��	+�Hw#�~}�2�6l1)a�U%��Q��|VY̲���
�I�#�\�<@'�o�va�9��ǘ�i��^�ZA�=at�W�mBm(S���/[�����P��,���@Y<��<�&�L�����@��D[R����A#���m(,Zd�{3�����5W�89����Y��"?4�<W�y��}q��Xg��7M����+ ~�[�	�/yR���C���3:x��\�j�-X���	}+?�Dg6�;�]��.qPlӄٕq�8W�!��0_�z������5#��h!9M#뜫F��î�!@���)C�Ⱓ�@b�;�֊R��+��]j r��M?[�Ns����ƫ��C�܉��;��s�Mn�͌S݋�ǆbM���mq���n�$uIkk�$؏
Mxi��d�d�h����Nfs�����g�w���HN쁺��@����S�J��:On�n�·��a
�����SnM��}]t%$��=�C;��Ƨg%8BQ���7�,,s�yo'�0T�d( r�5����&\[l�����O��F��T6���&z�؊�$���̍f��bj�]Q�B+Gc�g�_M3��.])��؜�j&f����V���v	n^>�I�����v�]|MJ�^�����4 ����'�%�z��k���EL�
�f�򌴙:��D�*dˇ�s&f��VVG\�֝�I��������a[q�h(��9c���*�l��;[�mr~�?� W EϽ����S8h��7�)��)�
M��}�^"w%sPuvlѦ	\�|�.����Kβ�r�{����Ք�T�k\�*vó%7���+E�4��c�G	�f���_��~6Jl��u��K�����ˀ�����un �/|�S�L]����x�y�����m)X�5��o8(��=�_��z����S�C���(Dh���`X%�	�!,�m�x�j׾����p����>%��/���q<h�s�G�"���1ҍ�F	9���ĸ�2O#/l�i���u���0��Ġ���j�+����W�vV�,���p��D�X�7\3�D4����G���l���ŝAœU�U�M���0���J�9�(ʱ�\�$�i���Hq�I���u�6�j-*���Ie�o�X���:��E�po�O�xWh+���g���&���@��/��@R1�=,%�S������ڦ��[���K��95�I�j/.�� �"�3�×�i����d��.��Q���N��#����%ƈu�L��[pp�=�g����.�5��#��5�	���s�%����*��I��B�sW/��V)ԑ+����X������ڮ*�dm9i��"��m�"����.�!�綪�|9Tr^aX~W�.wx������8Ӕ�5[�����V����8�\�6�6|��'�h*�<>zfD܄̧�G*L��b��_&��G
7��L�DCMT`wH��ɵ0�an4�z�Ɂc���sr��V�IG�#���x��oNo(��J����jAc#��f�P�+LJ�ml���v�ɴ?�xo�R6s��M�%�r&X!f�|�b����f�/�͍>Z|V���7�DG�4!B���0�}j�!9�j!����C�n?�*ѓ�gzu�(����п�D�N�[�'������$/�$�3@`��d/㖺&*Q�|�<J�yxgc/�4�K2�	-�8�|�?]8@��b�By��Ǵ\�V��)�+��"�HEgvѓ$�0d��n�уcU�xCX��4	���o��M�UY���C4(�G�R5 �;���L�������Y� ���B���	���I-��[VAN���������?[��lx�84y`�F1<�4)����*�`�¾��'1߽�m��?��Y�W���V6.u�޴M��O4�q�����Cק�I�%��Do4����@`=s��e�N
�m�L�Z��믪����yފ���r~(��e9��"�}ō��
�Y�֐훽Az;�ק��ZvDv$�$y�5��E��q+��_:ES�T�fw��[Z����`�+����3m��%P��y(CD2�e���{YRGB�a�ݔ�I�0���+�����:ˋd���__�x�ʒ�4��
�
y� ��(�6�U��{�p�s<��z��w��~��9&{OӦA���	�޶T��c`W$����y��th��U$����������^AH{�7Q� 7a�Y�y������5�M�r!�Dw�F�k�J�p��z�3��(�D���q�~"r� 9+iH�#��~k{'u�EU�b���Mj�8�
�]؋ȴ�NUhE}��OB?��BT;���(�l�-Dü ��{�vs(B�p ��h��ӽHc�{?\�ꟺ'h4�u�闱���v�Thi��R2Ꝙ���q�ga��Fm��嚽���G1���O���u<ƂrɁ��ۗ�
V�Jk������:X�ƙ�C뚿Qe=�)���*4oM��t���m,�j�#���v����@�sD.h#����ʍ��H�4 �.-����uu��K Gd�u�.�CW�a�pe K�Ѽ`^[��ܳ�M�х#g���;lbɮF���UW�t��a�¥���pVs�#1��rb���)	:����-A���E���O#m���c�Uޫs���������_�W��1��g&f�Ւ"z��W`f�1�	��s���(�{��d-�=*�,fl
9n�
X�^l�v*`�P%�����k퀏�k%�&)�~�M�U��s&���T��L�<
�Cl�e$JSI�74��"�򝏗�j�pb��߅)��i�&7���XH\a(�K�Zļ��h!���$.6B-$._��7���1.��N�#���)S��7�n^G@o�(0�Y"(@Pc�D�ױ�@�Ƽo���Z�>�lj��L%9���#��y|����֋�o��Gh�OmJxP���w<���/L�2�Јyş`É�bY��ِD
����oɂ�F�RJbZ�� �؟�"&9|��pL-I�۾�0�g���-�G�N11�%�j4HMǣ�!&R�g�IR#�Wh♉�VU�P�<J����~���z�Y`��c�h�o�n�cbB���S.�}�������������0> �5�Cq1F�:%��fνS�U���I\�S��Pւ�>7>�y�	�]q���6�#B�p:9 ��$ie;uo_(��SQv2����|`��Y�5�G�S%�_��J��Z�ו�%fO�x+��P�XWb�����R��S�����G�xP}��!Mqv��X|{����Q��?���ʾ��V����ː4����ܲȓ]孧�L��#R�qE�Gg�O�@t-T�I��=����R.*�r7�d��j 8}�u�z�CK�m�z�5'^`%c:�e��5��`�0a|�8V�D!��p�Y�dK�(��K�3��������1#���`Ҥ;ol�X����l/)�@�܎��{x=�y� �� 'φ�2�a�����@)}�0pKf���;MI���M�"_*�*�O;���,���2����&���s.q�x+<��/k�i�O���lPC�6���Ը1�gP�(��2 c��>t��ZO�RG'�NiD7�｛����A�
��I�fDN9ƪ9���&d{��A�DY�Ҍ�+����.C�S!K*�mj� �>��Dy��غ�}Io��� �I������-����C�QB yEz���8��p�S�z�ϭ�k�0y�z  qH��խx�3��G�c�[�케�X��,�莎� 7�J�(�"K:��>�q�������,zmkk�m��p���}������A�t!N�,�~�L)��ؿð9�}��`�$���x=����H���X�N�\�o�YWp��gSo��6��dI�h/�QXs��}�V׺�p��ro��>�B{�����Ո�Fb> KRf����H'�u����-1��)!`�C��dׂ�?*���� �ܥ��x�S��A��!8`W�K\�ê)�%Σ=u*��.{s@kAvQ�+G�g�	%�K�I2>���'���k�Ec�
�r�u��$���}����/�s�+��*W���.M�j��bZc
���g��>��C�tL��,Q�#O�dY��As�����ķ?G�"/nH�8[1��Ycs.�N�T4jE�u�us�XZ�� |�����}%ݣZD�N��~3!�(L�|H5	",�Y����Z>%��)v��v^
s�&�P���i�n�A�!�h���:38�he46�DJ^�1[�[#q��f}#wK�W7�tfC,�nA��M�h�u���B�;(b����n�3x�����������z�
����~�t�m���
	ã��#��࿙\w��s0���5l;j#<���a���F��Q �NN��Y�1�ˣ��m�!����$=�g���ƞ��@�T���rK�:lv#��S:�����G(lV���+,ۅ�A O�i��64���#U��Һ֔v�g����>k'</xY�Y~N.m�n���E�J}����q8μ�\|	�T��G���@��H�y��h8X�Mv�4���klB�F@4]M�-A�
��6y6�kx�s,�zR�v����6���f!u.�bGuts��F��-���4Y��k��Xky/�>�Ƨ�����U�L3����B�5�{���0�A2f'��ûya�	�P�%���1C���W�+
 M!c��2[���uL�M_}+�������j�Ec�K;Xo�|��P5� �/[�2�luI����j&�C��a9[2�}_E�����V�r.�(�Mz�IL��k�LM���r�h^ћZ�K��
��V-R��<J$�ܙrr:���4m�gh���צc�����S��ĳ�H�ޜ������t�a&���=٧t�M�|3t)�B����muihN;؅��){���"�,S��Y�p}���6*}��J2��7����(�Z',�����?�l�9���g�ٮNm����F��qҎ��̅P5� }[aVB2���r2|��}��_	�~����)օoY���EQ���&����}�±Q�0ebo6/�峼�1�&�m[���Ô�&�x'K&
��������F��N����єza��k�HO`�=}����I��3�}�uG+������i}��8@Ž��N@f�T�id!�[JnْwYDI~������mйe�g�'�>Wg�,�4bD@�y(�L_ͥ��WX�.��9nH_�(Fe�3�h��ζW;e�)Ml��l����{q���K ?W���o��NY���[�!Q��j�&�}_���a�"'� �*�{ř�a�M�1l�z�q1}�����_�@hJہ���{��py���3"zÈ��c�΀Ɋ#��581�Āj$��8�h8�%��.-8��^�ߥ��������j�Y���>��漤6��z�9�Bd�Q�y!�ʥzZ�e�:
��-�胿���}����J����ҷBe�~����/;�R�0h��=�	��hj�V����\���bI�*Yy�j/#�*��t=-z��@�P:���6s�j�3��]����(��:�`Q�q��z�=q�Wu�dH
��9�rkxu-�m��Y.���!a�	@������eO��uQR�E��A�S�W�ɝ�3~�P�h��!��M'p6���7V`�P�������9��85���?1��f��bGn�8��	K�;���4y~�k�(;X�ʗ����,�T7����M�K���$H�*��Aa�kYu;�H�Sr�lL<LUd���|:Ek⇶��Ov��'��BF��d�UH��2�wwP
������'�c�"4_#�8��ed��� �ACy�����![��E�����t�O�.��r���Y7	/8�YaM��*��%����pKx�k�{s{�ꈉ��i�g�ſ �m�cB�,���O��ik�F�a�.e2�	������
AF$�e��/5�r
c~���5��*���_�t�$���`vp�M�����&�2��a���\�WlA��� ��}��՚lui��\�&����Ђ(�w��X<�I��a7�J꼶�i���킀�L��,�0�a�4���ߍ���Dr��חw�m�e�eNz��/B��l�ӓ: ���ױ
��2�Z�<�i��nY��,���$5U�uV��Ύih	X/X��p�@)d'�4�&��T�;�L�wÑ:۪��n%��0���p����^�\��$;]�Ǎ�������	ٮO�'o���7�Z���fG�yi����2���g)�7�Lv�gw�}�O丌��=.h�a�Ȟ������{k��vߊ?�G�$G���H��F�bj����v@��)`��������ʻ"
"ܓx����3�Y�*�L��0��S���xRlE��ˣ����.����n��}f�nM���{-�5���Y���dtu��I&cԭP�H�1� =�R��Q��H%�T��R��R�o���ճe*��p��7B�x�=9��TnA
L�D2З?o��:�����L���K�9D�p�/h�C/-$�1�JK4�2�؆4��k���]��V��jd9!9�>��ci���`G]�x��Nd�;o��p��T�ro&Yǎ�Ai����ڼ�H��j-^<�K
��������`1��e�qkU���\�m�4����շ�%����{Y=�-:�t�>���p��蘺3(�	���k;"g�y?��9	�juh|����6��-�x�������q�UZ��J�Lr�/�ؖ�UB� %ᕷ�����Շ#��o]M��Q��d�i����"�k]��z�B�L�ɸT^6zJ��S��|��c��~[�s��Z�˶�ܺW��O�
��p�З�9�W�˅��nsPAMc�N�hV�~��絅;�M�p�dk��\$�G;�}�;�^]?��NcG�����+�}E�����VR�-�rf��g��`b�PR]f	��(?9�J@.��%�
p�[��{�rjC��V�d�Yh7�� �O
H�4.��x����`����%"ָ6TMs�^t~����ǭ�uO�����[�W۫{�NHC�A(O�\����2�NM~��r:���3����A��8U;��'�r�_q�{LK��g����J��+~�TlU|���m�)8��8�);�=�	�� G���fpZ����zTY��W�h��8��xM���[���,c��+��?qG"�3m9#���uM�J-��`�2��Le��}��r��GA5a,��J-���R�Pt� ��+�;M�vZ1�����dtܬ��c�k��U,��潗�Siߢ ��lk��D]�!�H��������ϭ�H�Nbƅ�O�n|�B���>=Z��38���`��������~z,�RCޏ7¡u\��ܻߝn�Mŵ"C�����ϋ���l��M�Cd�[2�6��0�`�d%���� �-�0l��:ba��|U��֩��\98��Sv��i`� r���e�
�=f1�G�u�}���^%���6ԃ�s��x��nO�*0��d��J/M��n=�AL�<�"�(茍�w��8���$*�m U�;�+�����������
��H� �������*��ZwC#�w�pT�_��/��T�m@6��u�F�����e�;U���������;��]�����	��N�V��j�\q��� g�7k�N�a��1�5�4mʲ�|����*���bt�=�'>@*�8���? \'�%��F���l"]Gy�1�Q�_�g0k��L���nC�SS�����Z�.�>�(����)���Y�~0��:��q�6��6}Q\�YK���1���(���B�Â��\W͙U�������Ӹ�`I.�n�s����Q9������B�=W��/#��V1��x9٪�9T�K��ל?5��{���e��4y�)؂�,[�<h�F����D���s􋦶����f���+6'���(�Ǯ��`�56�ZL�L�\��1�d8ȶV[�8�#�h}�._5���  �oLy?z�������NA�}G��ʹp��B���|E	���S�!�H� uWӵb�����p����L^�D�����%8�ww0����'4�)]A��M}Y�U��6���^hx�o��3>9�m����VcW?T�I�Z	�%�u7s��&�`����!�P_35���ٝ��)��Rc�K�Q��4��qv���!dag wâ���d��%X�}h�ˈ��TM�H:��h������5�$6JF=����WtZ�l"��%ӫ��n�e	~!�4v\��`4�~�n���m �?�vn%f��b|m�*����HX"H�zk�r�/���P��T
���U#�)ύ�*�^�{5��+i�n����&��"��S��r�^} ���i�7/�H����	�ZK�K'��ć<ƀ���x� ���3�}�t��d�K^��/쇪���T6�XݚЧ�[�eK�H-��6v�Q�⡩?%���
h�W�i;��hX%d�	-�'���ir ;��?�2��&M2���a$)�g�6M�,�$���iΰ��	��k��L�M�>bηu��=�MHWCfQ&����!ہ#k:���d0��J����W%>P�Ɠ/Z� �W9�t�(�9A@yK:AN��� �k�;B�U8�J�~���z�y��sK2=�Ė��c���ZmB�幌��g׉��Э�}%E[�z+k����ӹ���z����J�2�#7��П�\Nb"�ٔ\���9\��#Z����e.��H�b*�$H|Ɔ�Ȭ/t��~l������D1b#��v���N��8�2���dT��;O���Ï��w�.꫏��9�Y��1��J���!q(9*@���; zW���e��Db�*ҩOʌ�Q�e *v�DZbz�"�Z�q��^�VD�z��Q�ԡ�d�Tj~w��Z���v�=��PZӘ,����ї�`m�YY�)�t��}F/�N�Vݺ�66�YI� ��T�2��?M#g���@;��O��W�
 -��q��9B?�+��;G1����y�a�sս��0Lcb�|���7��/|pْ��͂N-�y_L��4\,��.������t����
b�`�Ovϭ����7���P�N��F�&��}c�����A�� ��]�ŋ����-#��J�������9�Ƙ�a��]�F���+V��-��V�k �G���+��r���vÏ�^��E&��yp����N���e<��µ���gw�J����KT`<�sOK���2nI����<U�9M�^|��%d�jP4Ӻ�J���5����<傿
,�#��I��|� _=ĥE�Ίm��K�dQ�y#����mQM;�C���n�1���a�U.R��
�]�HO" L�?C�?޲ש��鹣9�0���*��p?��O+s+@+��I��Lt,C�KI�$M|k�h:2Ud�~��9����[�7�%L*��_;��֨u�$�q-6���-�IP���v����ߦ:�2�����~�ϩ������PW�n��[`�J�/D
H���\����)�8����z��'y�u�5]3�(~�x�	r{J�I�}}��ܑ�����%JS辀2A���_&����������:��F���M(6��3���l>�p/�x�_�<������R���l���t��x!t1���㓍)?���A(�G��`I����7����+������H߾��v��u�5U��+#x�<2�۔E�#�jG�O�pr<@�VvMF�\NIH�#{�`�ۯ����ln<4�	�03�W��Kb����!PY5Vy-=ࣩ���@��$:��z+hx.�����!�[2X���쪓����[�Nd �J=[�EIA]D�sG�x��L������/�[[=�8�ݰ��L�U�R�m�����է[�3=d̳��Z�{׵�����#T�4xo��
���ҳ@�-����o����>^��8�ꏝmFGlß	�\���V����^N�nW���������s����O
�[:���]˹1������Xw�ن@W�m݁H�R�k^W-m��O�U�T��Vp:�w3�3rN����m�*U3���=*�n��{�R�Cyq
#�|Ȟ���ˑ��d1gEFd�2B+NA��s��oO
^�ͣ��m� �vGaM�4�F]A!6,vmuƚ�07�+�LT�F�Fٞ:e.W �v��Ā����3�� �P�,�	G8��Mp�~־��uD���K��FuI��{��z�^dR�0W m'�_�Քx�����C#h_��ҡ���t$�6X"�w+t�|p�S���f���oP=��*�ε��h�%��O�Dd�'���8�G����u`������8P���ty���}��^�L\����o�&G��P)�i�DY�<������U�D�^��Fz�:!/#�1�w��:�T���?8�6�F�a���羛�+�l�Z�e�N�}�����&��>)K��G�VEE��f�`G��~�8�ܴ�T-�G�G�{eU#"DPaϺ�<E2x���ǐ)�8���L�K���ظ�G��n��R������	��N�����8�wУ��nA$qF<;'�����24w�"a|�e�	{��y���h�Wu*�\?��	���{hbx��6�X&�h�awM�i�kl�%*���ts[����#�m��N��������k(��#P(��
�����Q~B��A�i;bb�񔑼<�~��(j��`��I?XG(�>7Ze�%f�\��r?%������1 \>�2#ɚ�HpIy�|�x�P{@��iq�íf(AM]/3�҂���Ӷzg+X��*� Ɛ j5���y��)K�kMf��Q�����U�[C�@ ʲU�7���F�7w͵v�O6�=����ny���>��,ӽ����,��!U����`d���*��.,�����zI�C&q'Y�ø�҅�0�o{Bx�q�0S摜�|�T��qa�Cu`���WT5����c�����$���S����4=�z�'�?ca���s-A����M��`~~>�6Ç�f�c�{J_��YM�=Ƅ70pe*f��x�ʧ����L�Ez���0�k55J��Iڲ�m���ݰl�)��5���ejc��1�,N88��͉j���l��Vȉ�"�� 1���P��$!�`��XG�F��计�<�9��w�����z�g����Ѽ��+A<F�R_�9�\�&}�Ac{��>�3Z\n�����;�cW_��e��J�#�)VО�%�`�W<齫�o��>�^�4d}[��%p���8K�O��THքY'������NQ�/^��͸�(0�6ܔ���N��l�Y�2ݐ��j�h��$+��5��&Ki�U
��0�ϣ��@o�K��T�M.{27�eOG/�(��;G`���o@8�$gߪ��R
LD�9�t><�?���Cy�xc���	Z(����>����|QT����Q;��2�0�
:TJ(�&��7�Oȝ~�u��3zeĩhB�:��s���ཎ�ύsq�&�{_;�1.�(���� ɡm ���!�"�5����;��aط^b�����0)�F#I"��+� ���=�r���<,-#COߪS��q-�;����q��k3z�#P��)x�(�cy]4��K����iʒ����϶��X�����g�zq�V�:�(Q&�N,hҰ����,M�V?��5��]�v�w�R�u-�	N�"����t7'>�t��q�9��n�i�|�+��Ώ��N"p���짖��G��m����D�)e#Υ}2$va�0&�F�R�]��x0��M /�F؛�T {b��ޟ�Ʀ�Ij�W��saa�7i�U�g� C��8@�����-�~�%��4��%�Y7S��H]";�:<��Е����Q�`#�O	:�B�M���{��}�օP�g��^��k��Ύ�=���t���k�럠KϘ�t'>���~�4�e�mv�V��cw�d��3��Y��x��R���qQ�B׻�$�GԀ�WN��k�\;�	#|x�\1mxe��aU5�ڭ`�.�;P���AE �	���a\k�ޅ�B��џ<x�Ζ1r��)ڄ7��\�'��5!u��x�]�Ab����Ĥ��a�lP�ƻ^��^�-S�Y:�zu��M�os��/�u��c:���crEeZ<�Ǡ3��LE�T�g�Y�����}2�Cz�)t%C�w��q�w�jLϪ#t[g�Ms霭�ގӒ�����>�Np�M��]�P^��.j��#���j��� �(7�������' 9�g���i%Rp�(�{�y��XWBPq���qj[>���٢l���$)�#ި����/�V�6�'�*���_�{� �O:6rgf��`�*'������E���� ��{t[`��S/�
H"@��a���>!Q�1�ݳ�0N�WΒ��[�d�D3C8!#��$�:=}$��
}�f)ܱx>^����_�2e�D��=�m���kN�%[q.�J1���:Z��5.��t"6W�ϹmG�T�Zjb�s[֎��X��ҪN,�EI�(I�D�zy�n`#�-]*&)��uh�r�,i[�h����N�4FT�ĝ+��<�ｩ�|��V-�#'�ά=�&>�%'nEEsp�2��D�aemWI��7���l<�Z,?O�t���a���V�<�a�J�Y����jw�s�J|"p�����[ٔF�AD��6�'%��f%fʥ����ts�ә,���,�k�:(2��ɑb�';HZ������X%������a�b4߽�X��E'�=�Ƴtq(m��}���qؙ�gR$�����u��y�{�]#�O(�G< n����Vnͯ3*���bb�E�h�����@t� �o����p� ��Қ���E	lVP,�;�xU��z�ոsĩ�N@�,a�/v��pd���v<��N�e��&-��?�%?C[�=�U}4�	�DOl�2eM�x�R�
�S����S�7Ld��L�6\�B#c�P�#�
�b9\�2����[�̆��&̏"��*(Я���OK�=�NEN�����s�³<a��W9��F����GWG��j���0z��Nd��^��n7~���Fۗ�~`�'̍����fUt󾶊X�7��s)��k���ض��EN(�Y �]���>q0�1���_d!w)zS��<hWD=Ю��~��-!���ݳO��	�mӞ��M��M�jȅ�B����gG@Î�\����~����ߚCt���©Z��P�&q�B��ǳ	[*���R�)�G�SWX"���*�����A"��&�x���oӄk#��H&n�phDY������Ε�"$�g���N�*j:0%9v}���e�0���D�%����������!Oǰ+���Gq�������?~�X����0�Ex�J�է,RÏ.��b�,�x��[!
f�w�	e�ӄx�7�n���qB?���Y������9ӕ�t2IM�0����\��X)�5�(��zd���&RL�ćf���sw�a
EFv���k�3�r�m{!^�Ɲ@���s`\��=�[.`�����E�ǥ����j̻���\>Duل� ���(|��؇��*��d��._{��\ �|�I���;��a�~v�����x�=�x�'����v�(_�P�g1�� B�m��Ѹ`'V��]��\| Q�m��uȻjQ*�Ϯ�\2Mf�\�44��D��C�AH(�Z;ih�[�¼���iSQ���}�`\V�I��qu�3�b������3���+o�a$��!��n�F:��ɔ,~�䖘w�`\��0L�*�(��,�Ϸ4J�R������9rmcrA���瓘���ʡ���V�w�'���:#><C�E0���=���/���C��V�]D��Э@�x�rrW�B��(�kQ�Po�@��*Q(�`�������u���V�EY 8iW��.\�����U�̜Z#e�Q]X5����_�s`2#|��|B���%wb�~o��N�b���\w;Z���0�%ъ������3� �Y�&�#��]�v�݇S�T��
NL�x��!Ŗ���Չr��0��C�>���5�� �����p�5�l{��i?��mҰ�����D�� ��*;��e3*�L2=6�<�v�CP��hD��G�9�T��G)� l�J�<�p#�S��9� uh��;��R��!*��^��$7F�-t�\�a\C�]F�泷}ARbP�6�mO��HȾ��q��Q���Hg�+eE~�L�+��pӁ;�<���9�;f~�RE�c]�SWo�s���4�����_��.ܓ��R�����%�l`J����ָ̝ח�T���i�F�Һ�t.����焤��Kߺ�QFN�ԡ;d����K��J�tQ�۷ו=�,�`��$m�{���S*����e)�XP�Rƨ1��Ӎ�On���u�~ۉ��i�bW��l�S�9q��DN���"��e���x�w�Z/r|�	+�+8'N)W�lkl�1�8a��Е��Cc{����l���Q}ʔ���B�EC㜳�:;,���*�-H+V�fw�4#}z�U��<�A>�A��	�7«]r�Nj�>���
�[h�i^�\O:}�ضI� �u��#S�ĸJn����DӵՏ���OVtu�e5=N��`.��龕�]i��xz=i�y��x��7�`%�l1�^0�9���OM����p{$��I
��>�H�`�?�r�}]yn��G�(hMުq��ɯ`�z>�<�}wpL�,�0���b��j��?����op�wˀ�Tt��%j��������h>2�X"�ٔ������r�z���[�1u��Xj@5��}�՝e(([Onia	k8��u�49q}K�N�p�a����T�����0B���p�!N�`J�y���z�9:/��%8��h*"!�Mb1���y�_�=^���AȬ��:��Ãqw�}�beB?	�t���Ԋ<f�����E�&F����E�A�J%��:�5�´hM�-j��G�X��|O��&X�E�HN�a��/�:1��Z�9V�F�*@�n�I� ���N=�v�ƍ���y#�s�A����O�������'ߘ��d��aa���B8���8~>�w��u��O�$N�v6�[����Q����\���@����#��A��SkQxss�1泏F��V6+�U��-��/yte>-D@ƃ�PG��w@�y�=�4a�F0��T`8)1��+V�;ő��0$�c��:;�5'��BK�������o'��A鯫��#��+�*��J�t��H�JLѻG�?"���ظ'��sua����[��5�*��r�(L�Iɯ>�W�x��L�k)X�V2!,�j������|67�p�,�7jʄ�vJ�G���z\���gA?����{%�d�b�����!��5w]��>#	י��M��z�/�kӭ��Ԡic�C�$HCJ��+��
���d������ȃ�W����h�C�p0 ��2�_i���|�K�=�g]�օ	�+:sz��?m����轣�[��-EI�t����qr��X�	�����WG�9���U�� ���t�|pTc��4�+2�RB[g
��l<����)��A#ĩC��N:ws٣�c�0t�|�!C��#>_q�o��L���9uS=5=J��ګ[ߊ�n3�צּI��G-�@n���Y�å|�|
}�ȼ��cᠯk�uBz���盘H5��X��	j�i;1m)��vS���%���HT�G�I���)Ez��!����e�P�������(7�®�ƴk0�&����d]Þ�;�)aQ+\�����X�}��-ż�iW��}��)��N^�n�!;&����cs7�.%��
�P\�H�=�� �Կ�����L ^(P�6
��샖+�2�w��/3�Ko����9lO��~��"ֿ��j��#�J�����uy�&���=>�$�������Z�%�X���Zi��;u!&��4�;�4#��j*D~?�Hy���FE���v���|.��Ge�,�7�h���*��k�g���O@�˵���
�Zo��a [��~*�6�pulP��.w쿳���@��yy����a���i8+D�xO�|��MH��'�80 �&)�z��T�c���,(\x�*�ӞX\��c��Q��ӪB������t���}�Z��Y@Z�-t�%��������'�I�F6���"`WqǔT�*�ָ�Z4g�5�C2�W�
��,���*l����o�r�Ҝ�˾��Q$95��1L��)�CJD�*�뤚?9!S�s��P}	��*�|#�U���&S�̝<8`����j����N��#��S�Fȴ�mg��R,8��'�os`
Ik(��"^<S?<�i|'-�>%W]j��>�)z,Յе� ~`��WF^�Ȕy{��@P��`*�+!0���@=�xB���-�Ȥe����mb�Jie�]�ƽ?�6�e"�z��
�p�a�X�[Y±�|c�Uo��eb�*ܛ�	m��F��0@�G�0t4��=�ơ%��h]�g1�oF���#!=#P���8L���1D9�AmsC}XF;���1�d�P��沎����t'q�ݒ����DW��>uud���;�rX@��}����
B��}�uZSӝs�КfȺ(|�Eej��}I��u"c����ܔ�vį�\ϗE�ּ�[��4��ѫA�sΙD,��ȍT>�o�����%[þ)\��j��7�3���4诩��KX�)^;�V���K�����B�R���;�0�{ElH��#ׁ����~�>�����22l�G��g��{���q��O�¼�F޺ ��Ѵ^9~3o�~��P�FT��� �>m��A\��Bԕ�fp)��T��y"�Wk�M /�(ϣ��5����j�!x`�B�6_����}���%TZ4�rC�����1��q���]=�ۑ��a�/GUTJ�.K���<��:�O���Ic����u��P �Q�} ��	ɦ�����
"<��B�'���Й<��WOp��! [#�}�l9)��ˉ��O�g����e��h���q������D�m
���H:=Jtv��5�A�8�`�Ц.�U&���<�L��Պ[����S>������O�����k;U�,Y����׫����w!p�����c��y��M�`��^1�c��1�!7Rp	2g�2l�z�M�	�uN�v2r�ģx)����W.��ޒ�`tso���DbRDf1=�WY��`��UKR�q�v�� �m�H�xp	�@`��ph4�%0�T��GO�{ ��BSfCF*��ϼWm{롯���Q�) q���V;/%�߬��<��8�FK��\��q����DjLVf_��{�Ǳ��`��G4�W,�	O�*�FKC:�+/�u���--;���2�UR���.�C9>u���b�W���``3��-�
Z!%����6ڔQϻ�����n�����8�q�#�` �����}����P��%���)�$���|�?+����S�ŵ��X]n�3����@;DQT��pu��H�E��)<��ۚf�k'�ɱc��E�{K�A���0!���~�6#�0d�X�@��&�S0DKs�Φ21`w�̥y X�~����[�<��ƍ;�P2�K�Z�AlI	��%�#w����J�c�UAN
�f@y�����9P,�e�]�2yh[Z��4ц���)�����l�%�{��"K��+�,�ё���G���Lk�K��1�n[����Y_�N�ه�l���!_/	L�g]Y��xe�
��mq0��pT(G�a�<B���Xg�wpaP!KP*Y�.,�כ��JY�`�v��Gs(�� t�I�<��T�D�4RNG�k�O�D����^p��x������y�o��T�:�F�A�y�7|�T�H�ݼ/n�e)��j�0�U�#}٢�-�4�[(ƻޛյCoR����s�~W���ȜWc?��i�����S�����M�7C�/:C��6�+���i"�=H$Z��y��ICrg��?1RcM�a�X�_P�� �ȏ�8�gv�&!I�D�Ո`uv.9,���RuB~��c�X "��M`m��j��2�qJӥw��lY�K�q�p��16����y�>��W_UH*)Śss�C�i`�:���
�z�4���Z��[���5��I�\H����2��q'�
y_%��A��nYD�E�f�暗�pt���[6	��,���?)�)	̕�����ai�9l{�\(�i������MJ)�f�z[ Qw? �)�K<E�n)���e� J��n�%���\�,���Ġ�$��B�����a��p�U�̵(��������X*����e�$�� ���Ν�p��7�n���+��Ns��B�r����1�a����:/�f��H�Jz!\�<�t�['[�%���#�l�<f91��vWþw��}kTN��� �"�ò���_!v�6Ba�q���J�P��lyi0
_��5��(2�m&1��<�I�h�
��C�R�2��5���?]��i��3��'��Mi�)-'���xz���}k����=�Z"�)c��5e�#�_��$��XS�"��3K���V�	��w)vBy�?8����^;^1��-�ΖN6��<��t�C����.�T5��Z����KXD���ђ�o4S��2{1�`�N��y�g�D�D9���J��G�(�(ϫ_"��w�B_��bÇ�PtO�.D#룫�� @>9�тr��l͌ئ�#	�^ŘTJ	اN�Q��W�\;B���Cl�uѯ0Ke8E��d@����/�6N���J�O�ao�,7���ˍ;,f�nHf;�e	���9�oi�I�����ҧ3��m	��v�~aox��j���{CI��{��d���Y1G�C�cfT�az���p"�e����I�InL��T��v�K<A�A��<��O��Ř�$JGG�����,���$��9%C�9��(V8M4/3� ���y�~����
��M抄�-�ܴ��4�
3bR��$N��1�Ea��׫`c>�߭sg�yA���J~����J0��48�H�`']ôc<�v���N��H[K��
(���1��):�o��G��S��ԗ�.�<xLZ�U��\di���L�I��V�}��ʒ��OX~N%�U%��T/���`���S����L����s�d�LY�=��F���F����]�Ա�Z�fs���)P���wǪ=F]̏�D>x*��1�o�pɎ�ݝh�6�(�;�)Ο����/"	�̑_ǁ��$ј�-&%��1�0�J�
�\���Kp���yh�?=�Ř��'�KB��P�M�O�d"H7)s}x͒&�?-�L�2���^�K-��#7��W������V�=S�?952��3N]�Z����L��t^�z7p�[���|��QD�wd*)�ReZ���a�-��q�ٱ����?T�!�u���L�`�$����hg�'t��vWbA_�$^�fʚH��Ԏ�E�#@���0O�W���G-mR��W?
N���lxLt�+NٳʙTpF\P�EW�Xg`�O�:���|�M��k�e�!$��,u�<����BHU{0�������c}L�K�`��׾d��Saa] �H`	x﷝֙i���^�ǝ���d��D�X���Z���we *���k9���|��F�of��:�UߤLRP��W�Wm$�R�x�q;�
}�g�%^7+/@���D�/�����m�IFB5*�>�V���6��}^�G�y҈%�uү:?��j����`��8�HPr$"��Ŭ#�j��9�5M�s�1B���[��MMc��gZ���!�������g���q�2��n&�"b[�]� s!4���^�q�=Sw��:��~����E�4u3��`���8�Q�i�%��b/��n��1<��,�����q�>�I[����Q�v �	@�Ҧ(��kv�M�1�D��?<���cH����WvuX�C�)�M	�-�er��p�uI�j��g�Q�$�X <@<#�5����C����W�޻y����sv	�4j��'��,Iz�V�$i&�^]����:I���5�;�}����.���� ��ʀ5������V�:�\`Tg���y��s�þB蠥�Y����<=wL���8��zp�7�ϖEr�ۙw)O	t��b���o;�$b�#@����C�z{��:U���u��@bM�+n���,���Hu�i���t��-�>������eHĸ��F��rm[��\�7S�^e{��L]�:��e�h[�*Ԧ����v^��y�ֽ��3���K'��0�ᯭ��1��wl�ҷv�)���`�ʈ�jAь�4�~l#E�Uݬ(~��B�M��N��:5:R��;{.f�;c��d�0i���U��>v�����h �i�τIy.e$0ک�сV�߄�AMD�/�ߘ�c�s���ӌ�eՄ�����.x��Tg.G��K�K˟
IBbU��ɍx�r�gÌ4��moZ��z·�"�Z)��q�K��+�PlA��Pwä44'л�N �����^&5��� '22���9ZcST\W�KQ��uCMAc��{b�ѯ}�̈��Z��	\)~(�Al���ғ��c����ꜿ�甜�Wp��#���M��Q|g7��=����>0Ш��dW��iŝ��x�i�����,��*�XE޸���K��2051@鷰.	�=Q	���ji�{�
O���T�G[LrO����J*|d��S��"yd�J��	��iJ�u����9޷ҜCxs�pP�%R�I*��ݴ�F�C_��LK�ԴH�k\�<����L�J
��s��XP.���Z�u���E�3�.�ׇT>M�Mw��az��.G������ہ����|�b�D��]�W��x����F7za^ߋ��%l*�E�ĺq,rq�~/����>`� _��?���@^���8�]mޗ6��Q&��&�؍h3gw�M�M����o�%�d~-ڢa�T4^�,B��<[�M���U5����)�0fy1�e�ů���߿ے%��.����dҭ�2����j�z��.�_��?L�����4��q�ǿ'=�?0F�8�{���(2\��c����Mp`zi}��,������"�"P�SVN�{��ۗ�Dg'�pa���:�f����:..�����u#��8�V�"�]%�(��U�;,o0����c��(�_ǎ2��������6+��m��\i�6B�j�rr3�w��+�z`�Fa�YYa�������(�o�v+��^����O�Z�wg<���"��c���Å��o�N6x�����o��r ���R����^��y+n�nl�Ot��d�����@�%r&�A���	w.3뙎ƘnL��H�0�iX[��+ݗ��m�W����W�N���t� ������#���2����*��N�W�PF 1�Vn��n�K?��,��O�t]u��B vAM�t륀2
�E*���n�$��Y��v��W��y4�Ϩ����QZݨW�+[����8�~$󋺏~p�Α�~)�yx(L�Q��o��b��̷�S�d�[�79��k���We�jn4��@^����6�o�g��&:�������Pz_�K��<`��J�>ү���B���̱��Sm�]�`"D(Ŵx�-&$���3�`��k����Y��R `����bj�0�V9utt�1Q�u�A��?�4�5P���܉=>��)sEj�p�V)��l^3$޲��w!XU'@㋜o����b�D�$�/���.X�vG��bפ��^�Ka�{�o	�O?�S$��em@���[���`�t�����O�P���i�(�}K	��^z����&�K��;�uJV�b�x�/@I��T��V��!
�FP��K�_��h9�t���+u��a��-��}ܛ�)��Hr^���k;�JO�xW�~���t��|ezW�L�5����O.kkB�t&E��d��� A~T!�B��2�2O��E,��^�L�_$�G��?��='_`|i>��C&� �\��$!2H/l"��HJ!I�����NyZ���Ut?B효�H�t�ϟiԖ�p�r�ֵ��¤�ݢvѿ��2�>�4>�2V��SpW�]����`̵B�ƃ��n=Y��?��h`���K��un�m��*��k���M>�T�v8ݖ<d�$|���-�x�S��4����^��A�L���3
��n�8�p�b �/e���&�bz���
��}q		_�8$�
��97������Y�ܠ)N�)��ѿ��b�:���n��$���\����m�Ñ��Ik�-#����ld�Rm!xF�F&�טO�||w֬�̔-nm��2�z�H�DA��+k/�0�O����\c����Y�5�t�XWk��s�H�{�(FYS�Iv�.P:;U�O�;�:"UZ<�ӘA�&���94CAq�ƃ�Y��H<��z}�֦B�
�Q�ɨw���8���!��P�tuv��K��
.J�@r�X��Ҡ樏�?��+gB��f�KN�Թ�#�0�,��]�no�B��<�1xs�^���\u��d�uu09h���{��V���*3v>V�Y �,�	�a*/k7����!�*+��yGO#�c�u��� qvĪ����QheU
�a藾Ԧn�'��4=5�����@���!#|�i/Z-�V	�'ʟ��p�����8u��C+g����vMg����m�f�2E�QI/��m����;���)��@�Xi�5(2ڃ|#JQ�}���+�G�R�	�+��j鶵��LZv씺a��?>��»��D��U�e��x�^	� ���x�7E����u�E����bM�^a�\�z�o&F�g��������
z;�C��~��n�F���wA�(��L��`��4�th_�'YM�_���3�Q Û"�LR��M�p}m,ʥ���� ��̽l�
�Y�hW��z+?NPx�����F�l�2�������q#�ˑ�(��Mw�� �_:���\M&��r�	|#cF'Z�}�D7�)2RG��*<��x}e_�{]�|- �!u��W�S�$t�$�Lf��iA�<X�@��[�\
d����2�9MHi�T �����Lҳ�Fu���_�	��_ՙ������mS҆0w��O\m�;%k$��S�૧1u-�Q[rgz��*��b-F 8.� 1~�����)��V1�J�����Ҋ�bFa�B�H
k��~kn��*R,+\~��2�H���ꖩ���X���]���$��/*	dиS��)AJ�Wd��0`D�z�C��³��G_���eN��!t�o֬e�~�s� ��J�_��vَ����n���'�7�4�`����n@��X�.-t�H��`Ճa§��`8��s{�4��
�'����y^߬�m��.��Ժ�i=j|=���=�I��2��~(�+neVc䠫�4?���bV��k�D��uB�'�u�4I�~���=��p���40�ѕ� ue��'��lb��We6m�_��������=Q�-���lh^�s�.�8�&���x���P�M�q�m��V4F�(E��C��F�x�����[�
cz�$���f��%b���J������F[��-��1��$�)���i��8Ѐ.�e0ފ��#�3���'<w�X-�g�Q�P����>^	�-�����aT���}�����U�� 'G�|O��}�O8�\��B�R�=�J��zނ��p������1�`�ŗƢ
-���)��TN#T��b9��?��b�ţ����~�Q�F��V��"�J �`� ��(�q������'q\�_c	�#�H���r5����:�3��e�C�~{�9,�ѩ�DQoJ�G��k����`Oe�2�d�ް.�.�F�3�~q�	k��MZ!��ؾ<2 jg����#aX�хD�nq�!�]Mx�6��{G��b��Q��+DQnxT\�li�C�[���v4�{�L�'pGYf6�|��t�l�g,$iʁ:Q7�ȁ	�ނ���g�M��^�Vh�E,�l�}����j~����)�	vf�-ː����O���#]�_z�ܾ��d'|�h�Ʀ�$��%�g^�1���^�s?�Y� �u8�o��_��	�%����4���nk �U�U��S�EI?F���ǔ�7�
9�]惵f��5���%��H"�y4K^jgKv�NCb_�K�I���3�&*K�?L�8��B��*���n8{'s��(q�����zvu��ߧ�Mf�b#Amâ��i���`}79@��Ba��1�����~fv�nDl��D�h��[�)u��+Pl�iY�l^�q�7@1gK�{U�5eAK���>��QZ
��R�Cl3$�L\��ՙ)�=��F&������
�>Օ�V����k�"!����1k�3#H�K-ҟ�خ�N�gjx���'U}��$��-A�_��@��=H,�=ZH�Ϝ���m�ү�-�~�f�!!G1�x�-@�V�kZ���aMD0�� �!���
�ҹ6�x�#���>�x�D�N]7Ў�g�k�q����L�4�I��	���^+���������Ȥ�OվL]~OH������Y�)Ř�A�֓5��ə2��+[Wx�Qf�PYdN��_�
X��1]:-Y�p�.�;g,���Nu|cv<<h
���-�4DB`�I#Ϭ�a�x��~�ݜ���q�c�WJ��	�W�Njl�X��
�Aj��v���7<���5_CՂ��� �90����LŚis��w����d�3�V(2�"��3w�>�_@G�k>_S��2��q/�q�էd�Y�È���_NT�s�HӼڠ�M[�b2"��|s��)��ke���,Rƻq��������M^�k��:<�1��y 2�e�@$j�/� ������h���"+�D�����H���[�-S�ij��t
9?�6D���N�4lX2���+�L9c���N��yT��D���m����ɤ�k����d�F��pt�C4,,71׭��~�'V�pv�̣|�����~ �b��>~z>����t؟����̵���3�v�����e#`6�m��Pr_uX��ʻz,̘��Ge0�ל���͖� ���<vgS,|e�{M���Ԟ�'�;�b����J�#k~J7t�5��4����1���@���ў�C79:�D��A��)��MI�KpW�J�"Q�����:\0�U���!�" f�gɠ�s���nV�k���݀�դ�.�� EZ�Qs�J�P*���� ��TW�%2r�.�I-��kev��Q�ٴ>xy�V؎�u�z�N툷�@(��p3�ĎT�s����	�8��_�	�u�t�Wi"��)u���z_;2��4� 56�eF_5��+a"��<{��8��R ��'��S~���L����������86p���ivW�AS	��@�gXR,~,3�e�xɏ��㛖@F#���+�V�����ʍH��xs�N�χs@�?'�����M���ÁIfXs���z�j����n�r �ٛ�$Nq#m��m۸���`=���x��&{P!��0o8�0��|���J�ڐA�E	��l����`
Uc��0�Qz�m7��Y�<(e�Ç9��5c獶ї�	�m���G�S��=�����h��U�0��9(ʯ�d�R!?���j1�����#�J��b�Ն�������F�Ŕ�ō7��,	�H�>]��/Co�5���,Q�{�I�,�+v��(C�kJ�^󚔚p3̞����o�d��T�XG^�f��F�~8���^"`��{�#��$��ڎmX^���0{ ���3f�)���k���7�uV?�C�ݬt��ug��������L��Q��ٯ��\L��D��މ�/M�]����l�[�����pQ.\��/1����n���Q�_[���s��p4�I��P��>��mр������Z\˿1�7]kT1eZN���B���KT�@�
�P���_)�L5I�缁�''�4Z4�$���9|��973�x��~����3��x���*�0� ,��?�|���^�՛#f�Y.�da�s |vU�4�f�I����~���6�z��xڇ#+��[&QDj��}iJ��@ZV��yCKJr6_��a�r��������F"�� ��$_�S^�me(��ՋҒ�#�gu�)(��cK��I��[�F� 5X���6�7�Lk��4}�O�{��h�8�P¢H���.�A~�ڟk�{Ƭ(U��[�D'�e��p�qX�yr��v3�t>>y�IF�OW;l�3TXQ�g�&��̧��������JmL:4Y�u�<�������x����On�8�J��l+p���l�̅Ie8{[�Ⱦ��TThhyc�a\aspY9�2pt2���Ohе��;��fS�NP� ¬�e����л�ԯ0Ҩ�&r��yn!�b�&/s8�(���\
�U4q0V�\9T��o �Z��P A�)2_Np�c�����:�n�L�yj���$-#�tо�7[��C�^|D��cpkMA6dR�J@����:_��3xEv��Lq��:��!K�Vg7��PwWU+�4eU�D?�;�%����t՝F���}���O��7&��X>��	o|,��j��=�0��@�T�,��zH��j�~����Ћ���p�4��_yՔ~�v�D�1�c��'U�s��M�B-���`3� �r��p�s���`���9P��Dզ&_Fz�x�.Y��V��ȣ�DNkP���]rZ{�����Io���	9���J�N����>*���д�� 3��WD^tCS��ڴٔg�^e�@4m�8�xx� Q8�L>.��~���v|�D�{祭*Ap�&��53�}_�c�D!�"��x�D�r^�9c����#i��byZƀF¾�|������V�V�;�/)ā��)�ie�m�f4�����C۶�5ND{9���,}us�M6yr�Y�5����ݑ���#��u��K�4��ʿP0R�Z7'��rS%W$�3BO��6���Q@3+�>"�F�F�L��5�?�fmo�M����	��[k:ԫ����*J�g�{7y�AL&�)�޴���&K[�!]��Ӥ��0�L�x'u6�4d��gp
{f�����z�8o���xW-Wȟhn�r^���]O#��jt��w��Z8�үYA�▮�u�6ع��8HK܁z��2@�x%�Ad�X���x8�^t�\63"�9z��>?������c%���a5�O��L�H���Y�"E������q)��4dZ+���&G��2�*X39����@qU:dA������el�?�S~ʴH�ࡥ����<�J ��l=w��eD8�z�>��ԕ
U�;��E�i�އ>�͢�DZYR�v��`8�b[��ZjUqf�#P��A��xλ����F�x�<�Z���W�E�>�B���zW.�t1=�֚5�Y�9y�z�~&��b+C��L~A��-�ɖ`�����wW����F�Ӈ7������\����)O�r[4^��<BN�sgU�mɮz\�|gC����6|Q���W�KJy���@����#!x�k^S�r�������ͮ2{}2eP��sx�Ѳ_��#�ۛI~B
`�w�W"D^n�.��2���YV�2�)�c���X>�1}��Ԗf
Ks�*1�'��r~����!���,������ ��<c��vh��H?q7-��IǮ_i5C��꿒x�W`&ީ��ɯ
�F�i�2�x����Bg�V�_�q��T��(H��<R#:��-��_�)��vIM{�D�v���S���V4��8d��"uׇ� ��vWt�q
q�j��5N��#O�
8����Ię%��Я���u(������
���ڽ���e冱��@�&�p�a�	H;̗A=9�-������P�1��Bhް�w�vk�a*�5ß_��G����8)����?ɑ=��q��/H'�d�j�L�'	��5��V��,������f�ɤ��*D�y�����M�7� qǶ�FG��\��*��D�2���������\��P)��,i��WF`>�U����\m�5I��F}�hJ�����D�;+����ÊU��ޓ�����xBE8���:D#_�4�l��N�s=7�I����o���4R-�|e:�����vA��>
ȑ�Dr�3��oؐܭI�l��RTᴧz�*{�ݜsk�a�ϭ�%SA�&�ߍ/�D?d���N��ûo�}eR�7�S����
����Q]�#wW�e|t���:�V�W;\&��sF1�"pcç���(�7oz׳�g[)-��ŕ��3G���Ԥ��᷇K�sc&��R�P�8����M�>����ۉ~a��L�rޞb�8ͪ좌T��2�v����g�vՏ�c��u(��6��Ʒ��o�O�BU��o�<	L�w8��Ԡw 2�LHI7���z��-�ǐ?S�S� L�%��ag�7ܗ1����j�2͘b||��U�iM�D,�V+Ǔ�m��tl3�ŒK �����qLx�c�6u(�Eby��Z�>j�2�B�tT���.�9�z�g60���XF��.+S1��`hftR�}��;��/�fաi7�������n�-:p���g�0�!U�����v/�Y�E������10�
A��ɔ���n%����J���~Ax�.]��1�T�	�Mf���G�P�0g����`�]	'�C���KM�t=W%�@z;�Ьu=�84da�תQݤ�}��Tw�	X-Z�PQMq@<\u��,ݤd+���`Q"Â�$�%�5q�
�CEZ]��O�.E&�	Ҋg���JJ��K4k��U��A�� vh�1r�.he��w��Y~s�c!�R6p��L�j��ibk�m�˺n���A����?!o�B
�!��Ӕ��RO��?�M\��07��a-d˅<�}�P�k����h��W?�5������EX�����6j���&�00�)b�84֗���ۓ�ؔ%��#�x��u�J�Jى�f�sN(e�
0k���y�3P�x�H`�?�aka��`�	I������*�$
�9���?ρan"&��Jƀ��~*
*n�~�T�zM��6�[zH������n��2)X�P�n�UH���S��ԃ0U�_��g�� OU!� mq��1J��Ae+�h�l���n�NB�xC]�W�g�*X�9��0��V�$�S"���L)���s@��ӣ;ѓ�Z1v��0���_�W�g`p5��{�	x���=j���&����d�s��ZfJ��1x�VA���g��"׹ψUU���c��g�h�&"����S�7+��8�JW��c~�PE��eH������8A��tֳ��.|�C�fɰ���L��C*ᑖ�S��!������Q�OĪH��ܐ����eH��-����Tǥ�-��0��x7-�\��5���4k3�r
���/��wsمN Xp&��q�>7G�ۄ��Q_��Ɣ0�X<Q��j��R�[l��}�"C���σ9�wE�nj�O^��b�ϟ�th�	�H4I����Yg�q�Ԑ�f2U�#dz"�<k컌Z�p���Q�A��p#D��A y~���r	���m�]_m�9�b[��=�d\q��R.�ؓ�o[�Qbf���񦧱Ո_Q� ��v�K6��w6WQ�y�P(� ��v�rzsbpPFCށ�\�m���\�`��@	��2r9@��]O�ʰ�X�]�
���U8K��'$�"�˼�ľϢ"ϐl�h|�W��%r�G/T�m��1S$���?{������i򂛬7�1��E'�Wrn5��&����x��9����G�}�@ZBh���o	��Q�5�i'=FFq��u�=�'4��k�b�s�h8�G�R��&�AĞ?e/3;��J�!�b�Bl=M睫\4����	��t�6P��01s�[�KφċZ.��N�c�0��wb� ��g
����ai��)1EP��f�s�?��M��M����E�#@:��TIc���J$9���F�7m�tx��x��GU�GH�3:|�ӿ��n\���{�J����-[Q!�g%���ն����~7֫��v��h�P9ð����6mOݕ��t�����$!]ێa�_��ޮ �+�*�
?,�#͘�v�(�,|.�2a��T�e��Lv2`ש����Wf��	%ߊ)q�d�{���3|-�u3��Q�a'��+���mN_�]^�����L�~&�K�|�:J ӣ��;�5���s'z!�[xB6��.u���b��f�EU��s��P;�ۢ.��6}�Y;��:��=��.)"<e.���'�Ľ���WVyR���_1� `�U1ߚ�^����T���t�,2�d�U�?��Zi7�ǘ�7μ���dVX3�������@os�pF� �YܯEVBN M�;���aj 
����j%����Q����G3Q�h�^����iot��yʑ����ಓ�i����HE��-sAEؽ@�R���Q��6�ڼ�E��&A���V�[W����o镖���l(���+D�xV5�N�0�秦߶����yf�YB|��8���5�z�.�"N�5�ٌ�&˙�\��wW�����ВX4��?_b�X��Ҟ)�
��ޤ5��e�pZ9�A�N<\��S�
}�5�������SS����.�\�	�.'��"�v��`��L_�/*�3�di�ӎ8*зaڬ�ݘ�$!�'��j��zsw���D�������1Q�Y�&:ߙ�!V� ����p�"$�G�ƙ>�z�s�ރ]8���}d��e�ݨL��yn�c�4���^��1����T�)|�[f�r�lL��p䷏R����
$q��|f8qɯgFDSqD������1�j�by/����h�� g�w*��;����T9�4RT��Nb᳊3ϠCe1����[�Xq�aHA� 2@�H�u�V�'����rĩ�j#N��R��K6���P�f5�x��䋓�B��������*�6��C��9��js��`X*!k���	ɬHs�2W��#��Ĭ�$��z�e8d10X��+)��Q�E�5���1h��{����� --,S_�XLAL�xƈ5I���J���?a���煖5�#��e��.A�;.ּ����J�p$��^�=��� p�_��k}m/���VRl�_��v���< �9@��ȋu����-�}Kz<�V�lL���[Es=0�1�Q=ٗe�,��'��+�^����!���[��tBi�OG��81����l�n��޺�aAT�J�Ι-">\\�yš��V�E��3=񴑒@�)2�-s���|��AE~�5R�:�h�<�z��MDV�Q��Yp�Og��L�jӠ�(,������<=�8�����)8� �UE���өu�I]wJ�6���O��.���.�Hj�;�ss�@�z|&u|dq�В���-�gº�S���;����ʊq*�m5�:3��,.	9��L��ꪔ-ʠ �k��uRS~���<ߐY��-�,9�������dИ
�Ԯ��w�iZ\SC(�6��I4V#�nf#o��	o�0��ugs����?�ri��`�?9���h���6	;M3*š��Q���Ϧ-���m�B6U�({k�������[����7�YZZ���(��C�z~�@y����蔺H'��~41��`h�p�!�֞�l�h���	���(Q�մ*O.^Mx��P��R�w5J��@ʖ���kI[Q�P��m�f
%2�ا��SB�3��g���m�/�H��3^���R�n���Nd��o"�.J��!�XP�\���hGy(��9��.*��Y��.��� he��z~C��w153¿<ΰK�O������q��,�d� ���B�����V�{���I���[�*���"AzS7M�[���9�+��iq{��U�T��� }P�8��WTIQdO|���Vα��x��^^��H>�	��=�u��EϮ��\^�"]�4�pJ%{R�
����C˻�m�Hw�}�Y}��.�����\p�<X��&�P'�G�{�����X?�y1@��b���'�����"�I�s߄}��%'�<S��fGaN�1}H���g��?~	�3��-X�f���H�<�'���1k�t>1E�"u-��MbWt���ă��)J��S{�߿2,ZN��uf9~)됚���͝l��v���� f�a�u��(��_g졎pТ��9U���_k�EF6�X�)`��x^�q>R�BI�.!(\f	��R�2)e8
G&�_���&�o]�F�6W�	o<r��_:��ɳ��p�m�� S���P���w���d:�*t|�s�;6��=�lU:�4?��I$��/�vhލ)2�a#_]Ƭ_wi��|z1���D?z���Y�,�䯄���ˈ?z��,������g������)���W�.�D�����H�&��A�M,�;0�Rb<���&~�6�+��{\<�a�)s�P@��X ��bP��R���uSKa��b#98k 8���C�)�K�ZYܙ��zc����9�N��6j����^���ߏM
$�����`�7xq��Y����;ʲ��ُN{�Ҽn�.�cs�̤�V�s�z�{�A����;���Z�\<Q�"�{e����S�]ܶ���e�;�!xD<�b
ߍ������B���Ai���L�>�3��z;�7�c*�p���	�0�:��Ɗ�����|��')$X.����Xr�7�ہlq�=��$��9z-#x`Ϫ�O��N���
7p@Ā��jS���{�)ήg�=Lݩ�mi�$ ��G��`���h{�P��v8�c��D��ζ�\�_g V+�z\cH8�������Nh�+h��&31e��(�D_N9VW�=��G~�͔n��N���)����򏻄�^�:�� d�J�������f����EP��g��3EM:������U{Wc��ԗUE�y�(�A�䫰U���O�ˣ�Z��r� Ք�QBsu^/�6*̙�M�4����ŀy�byw�%��Ԝ����-��;al(QLA�i�|�YK�=��͝r��C�ZB�i����`)+�y~���_�]�I�Қ^���>��L��ؔ6�^S�Q'Ji3y��g� 6�}��X>|�l���Yx��b���5�@�0Z,ʉ�F5�lM�*�`(�<a�M#K#�o<4q�)L2P�K������w��O��(�I���'�6�r��*d���X���d|L���YH��)���}��׋��c����YZX#��e��)�$���@��X2l?ȘZ��v�=v���n~ݒ�'S�W��㐎��ו|�s��[*��4CE`&��>4u�:��+F��[�M��E�6�u ��S�_�?�-'D�)1�$̚x�$��"Dg�,�X���NZ��D�a���zǎ}���d��a�.ke3�h���ol���Eji�����]�KH�T�ߵ-�����֯�V
�ʇS�y��x�����-S{��T��	���L@�ly��hce�ک��H�yk�'�(���w�8���� F�j���9]q�f�����ի�k�^n7%�q�ݛd���⻚m	Pjp�;���O^���.�������G�Z��. ��t��J���Xuq��lw��X�D����W���c�hB��`���pY�b���B��Fkk��'x6�Saf������.���5�&9�7
�
��H�}h�ʙH�_m[O(7*�0|��XhHy�;ga롇'��_�?�J�����\�[#C֞@�|��iv�'u�l��3J�������/����^�璟��>�X�����=�O����ķL���f���W�m���a�|�"�ۇp����u~5i�@b��y�*T�E�����]�O���ǎ��t�]M���t>�/}3{<�� �5D8��j}�ؾO�ʽx L#�O��2p >V�:.�6C�
��|�c��>�Y�E7v&����N��e**�A�;�~�m���Cݑ���A	�ǃ��HM	'D��8�s�Ϋ4������,:z��_鉘���O�c_,�:���f�g�zX�Fl�6�b	�|����f���f����8r�s��Ϸ�F���Z)���#�C�Cf4^z��f1�@�/��yN�8�P!���. @x����/��"�e�q���X��ܫ���p�Lc"�=�HB�t���|6~G�|���i�����4y�^m�C�&�mi�S*;���;P�=���{�eY�Wtypp�
�.���~)�6�4���t����q��a����% ��ZX������I��^|i��(ٳI֛�!V��߽�iebҜ���/)���4�Ki���!�L�g%$E�f��h�Q���!�0���x˘�xd�9�k�yq�	I����W)������2���؀�-.˂��X�����P�-hT�o�튿�D�9��衼����K���(qZ�L*������/�ʌAj���3�D��>��q��w�C����CO���1c%N�w�U! ���R���0��Y�!3�-W��o|�s|�7g}['�ehLڱ���0�:�R��ɼ{SZR�3�a���;����|�N��{* �`RG��
�9����Q���N�B-0 ����D��p땡�k]�b51r�3ǜ����0P�p(�T5� :�p���΢��%�vC���(A]���V�����z��)�:���g�����,��Q�A�l�nC�M����+<�=���.�-��U�")�/Y�(,�XvK��;�%2e����]�Jh���;����"�P���x$Y�r)�]+��|nh<��L?-L�<�Tf|+�\���qZ!8�Qz�F���� �%_�B��,�	NN�S��1�٦�[�k�ƭv#ي����A� ���:nvr��	���7k"��t�"-�3u�#�Et�M6<��d7��a��g�T׏��w��_����HBt��ߠ8�b��.i��@�q@�Z�t�i}��� W��P~��Wa��z0ו��IU03��s�U��ݘ�_����G	zEı ���G��lh�!�n�w��:�#�H;$��b~K,?���K���S~2��ƣb��𥳐5_C�x+X
:.��?2l����\��~��u�Rϛ@�<&�=�>D!�>3wK��97�w�wˀ	�$���ߟ�@�0~26��VU�T�+��8�|��ezN�W���ڜ�yg��! ծ*v@��O>��00������\j�� W�Q��]n �����l�Bf��x�l����-�9G��4��r�+9����I8���Ғ?N*�MP;��#�$�����P��zk�ǌ��t���1��>�kJ
�$;W4��p3O�db�BG��||V��:h�&���;HZ��qp�`���$J����$CLS�DG��.�a�sn�%$�v����m�����+��e�������6�L`�C	c�Ipe��ݣzϒ���iq��/˲`>|��i�/݈.%��ٳ�_g��J��.�1p���{����l	��AH6H�6��E�>#�h��~�r-h��"h��!'&X�(��m`���$��F���P��`�0^�JD_k;�� z�hks��9IƐ�lz�ё�ڙ��҉ZG��{1`�-q�@��2�_�e�g�?�dT�AkX"[��D��|"�`��>�x���C���ڇC�ʈ�-��eέ����p�P3�jO�NV���� ����]yOZ+x~�6APN��,Tr��V��k.�|�	��.�`uz"ra�׏�o���ք�����0y!ej3�=_�[����.Z��+��˦k�6ը�ƴ2;�]����To'��o����ܦ�z��9�m�����Gy4�O%pm����h��I��Fl|⫲�'͑�5�φ~N��q���b�1a|W\���#^�MoǨWl1.��U�(&\���/r�>����zK�1�a���������l���.s���^��[H����=[���^�@�#�t�l�
tC�%�\*  3��^r�v�x� �JTC6b�ț�e�}�t�=d,C�ULT4UfyŊ!��OӚ��ϱ�s�0��:״9(H��kA
kFI����j��&l�-�ݿ�VV��O����t>��6���B��2C��Y���΢�uD܀Z���{ş����ߍC��)����Es�!�Z D��4��N°�F�N�VD��k�U���+��Վ.�k�|K@M�]	՜�F�f2��u0ެ�_�D�,Y~�?-�!�:U'j�k�y�)j�'&0M�=�{��ս��a�+�XH��Ԃ���Wj�_��uטg��?��j��\���9��+�1�]=�3Inۧ�Ks����&0I|]�eۨY��=</�����|�`ꪟb�f�^0xn��[���s�I����f蓤����@T��J�R���� -�H�HQ��2q�b�wMT)��%�mOu(��3�1C��t^��_:����,C�^��{&J��J��Y�'	
���P\�
x��_ڸ��Vߏ��?��9j�a��35�f�o,��D0�D+HW:H	O�|���u0Ӳ�T�E+|x5.cqC�0<��ʝf��O�&��ӡSn����j�w�B�VWN3�͡:���T���ئ؞y�;V�DM��ןS�8^KS�� ���KM����/v����mpS��~Z|X��x�:��]�p����60u=��YgvC��|�\C���$���8��-R*�"��H��X�;nV��}{�U�ݵJ��$9���E/��]���rG�;�מ��gQ@Ugg�8����]�cӛ
��HX�˟�j�J-��Z1����8�_��_�߇�=!��<Y�pF��?S�o�cν`��u���Z�1�(��xƎ���`�v�r�����s9񧹢�{��6ט�g8_X�J^��(MF��/a�"��G|��!�q=���IK�F:<JRNG��ԕ�{q EVԪ�s��W�<5Έ��6�8�$�X&��M�n�m�d��p<��unM"��M�����8,
P��r���Ō�V����v1��rw�I%���@ET���Ը���+��b�r}m�״_ة"�Hty�m�)�v�C�cr��~��%=�C��DV~�/4��\d+�9}sSr�H@W���g�*��G���@�6����h`�-����b�I^�JR����,�U��[�Oδ9lW�`bU�@>(lL��*@�;�R<v�f|�f����XbƜ$N+�w�{(�ٴܘ^�3ۮ��4���M���M��Ы.�\r�~0�� M��(u�Q�n8O��\�8���b���M���hlB�KB4�dZ	���u��/=���/h��<�Op}��P�t�#ګkL
�D�T���6=睷�������}2���Dtd#�p��h<����:Nt�CZ}�.����sCP���*�Q㈶ѷ:��,�!�u�Zl�H�%���b�.:���L�!J�V_��{���y�DAuP����9�����S�B9f���|�b#�q(G��= ������z~������� �(�as�Y�RN��i-�nh�p��4Y��S;�Q�#J�.#��3�[/�j�Yd���l
~ ��v@`O�XQw���o����
���}�Sd4Q�� ����R��.��lc�vĂ��]$�!��j�h}��C~0I�rFeᓥ���Z���~�9��7	�c�	U�Ylm��D�=@�Jw��~�h�V~e�l<ڇba�x�,�~���nՃ���9)�ʂ����5�ٓ$���'��u8j�h��*^��ј�b>�# �����C��D��d��uc����sgB*�Sbݬvq�,ĹD{���'Z�TG]Z���
@ޢa��-�~&>�5D���b���F�._���[a�5��q����Cgo��Z?@����Al�CR��BLR@��Ũ�{9�>�w7E\ߙX@��Or^�>���}��E���cw:m&6n�����PFĦ��KF���y���ȴj�U{3o�Q�ly���Mw��K�U��5���;�di\���$ !A�y ������'W�hg��5���9�K�0�7�kߨ���(J��T��nr���CBl'��nE4
���d���J�6
�[��U�*,��%w�8�Dk�ּ6��}�Ȁ�-�=�s��~��	��X�Ǒ�o9h}�F�5�^��&o�Zq,�����Y����5ӑ(*�N��~��_`K��"Ô����u�|��e.Θ�(z��a$q���o�#�b��m>�p��U��m��h��BO��́�"�h+��ab�C*���h�	����a�sQ9(�N "�i|�6�W�h�O�/�u�gh��`�{�8j�c��QK8�7D��7?����h�P} 9��W��s�=x���v��q�g���l]��sG����z�1�o �������f� �H�bZڻ�miB�yס�r.�1��|v������T����c-�Df?�j�;�c��͸��$��m�2���M}r��cx���q�a�D@�p����2�R�ެ�c@��4P{� ��d�v�u�I�`�S9��tF�Ѱ+>����Ǵ�P�6�P�a��G�)-�?)��g�6[z��u_�X+�^ye�ꆊ%�k�V�b"N��v�.�+߻u�h	{�Wp8~�*�fd�G׃�ho�������,&-WJj����A8?o�!��L�g��bLV0���y�C�;��u"����C���̱��Ά��X��tգ^?��l ���}��g��K��L��f��ijŤv�KC��T5Z�5�9�0��k���Jr���b�+v1�����RHy�v�ql\"E�`�0xuf�*M㥾7]��YG��UM1I�]����x�W
;	m�,�nc��Q� �-/��a�2*�P�ɼ�Df#n.܆%b7P>��@�s	�~�2��i{$���L_��8KǕSɃ��a��ݚ*�-��ͯ������Rg1j#�Ӝ{�!�A��"P��kr] ��8%��tt��V �,��` '�SA�[�:�>��xێ�ǌVvC�1
#�N;���w� ��m�W��z�]aA��M���)�m���:��|.�\Fߑl��h��	�Ն����-�9<8
��Q�,]�5a���?�"�R�@�Ɣ���fn�ĕ���g�r�5��'��!6m�S ��H�+�1d{x�bE�qn	AЭVZ��\X�Z�z��N�եdݬ�����$G}�@Uc���z�[A��  �Xf�V��?ѻ� Y)�nW��i�M����eo�W躜{���ވ�8J����s�],8ʛ���E.���s�m������������Ld���b�����Ե�̀l��d�L�F�lW:��K�V�~�ׂ��WyA���ܑ0�=y�ɩTU��7}��z���6�g���P�}Cf�	s���I�k�z�\oҬI�+W'�����Y�O���%�,,���(�?/�:KF��x�a�Ēn�$��FR�#�Pn��*|����^�9�{�}~�@���7��G����Xa�"?.Nbo��v�p��2�^*H�%y�w~�S�6��g�4��)]Ѐ����y.[�����ŖB,3𢡄V:?+��*P����N�i���#E���$�:=H��>��Pzi5�92���6"�m�ToŐ�J�j�;SQ��9��-�]�@�$;�yu��],=PwD'�Di��7��O<���BM��� ��T2k
.=HO\���C��6A�,�$��?2*η�9]��C��t�0@'vq�"jg���jgXF؍��L��%��(�2Sֻ֖�	���G�@�p�$��N�Ů����;��V��^�84��t�^}w�S�X.�&���
��~(�b

cO;�Z;n街�C��$F��R��l
ޱ���lfV�^�X(����jes7Ozƺt6ru�tE�� ��"��c�	^�3���cwI��W��n��ǫ�W���9+����R𳸑%� �x��aE{r�Ɯ%�̨	��5�q4b�x��_�%�(S���65�~��E#Ӄ�<	dt�#��������iNK��״���E�\�\x���@�������X����?��$}��DF�@��`��V��$���΋���nȑ�D������S�0.8Bt������Q��+�_�g����y�MV�eȠ�\z����O��F����QR̕N!�q�Z�Ñ�yeV�mmu^6�@��'(�������YLv�7;e�Z��PvܿN���=�rz������C%�g�C��vwk=:\R��>|}�`m*�u�]���R���lc�т8�A'���9�.�p|���^��+��X���|��;4y��
.��?����#�[{�"�/3u�6��	�+x��~����y�qlYe:Nr?�7���l_nS���\��Ϩڀ �������l���=��N��4L��|9���x�ڝ�\
\��o9q�S]h����q:x��5���)	t��f�@�O�����Z����6�?��C�i:T��5y�D#���� ι�S#�f�4����u�E�j5�g~���ͽ�!��)M�Q�����ܗ��Fv��2���`!ٔJ0M޻M7u��v(�Z�wT�<���i�Y
�}D�t�Ծ]�@s.��!��њ�-A�Z!Tg+ȹĤuwF�ϟy�k�&�T��~�?<$FSE�\֒��0��7=�e��Ԥ�"^"8e�~��6�ޖ��.o�r�!R�7��t6�u�����c�v�%���e`6E��]���	뢁��?�9��Ҟ�[*➑�Ű[�|E�⫚Nus�<�o*�έ�B��R�D�bG��')2�׾߆k�^�*���}wɈ�;p
��:.��sƎ<',�:r��*����sw���DD
�K�L���nC�uRNe ��T�TsnR_ԍ�XB��~:ӷ3��	)�̩s9���ʚ�r>R�.�ϐձy��a�������M�J*彧��T�~BZc<c�����ǍGS�zb�򃟚89�D�v����[=rU�ۤ(_>�q���O��T�R�e���U:/�qͰd;��:�Їդ�S�!�KE���0�����8R�`�׸��$4H��|-�N��M�1
��.��� Z�'�rr�Q;������>S����9�ޫ�9G�9&CQs4��sñ^<� ���ѫݳl��Q�&QKl�R�[�I�� �p%�ݒ�5[Qp���=X�d�]�Q���u�K'�=�8�4l�7l���x�C29\`�:z�/����5;�Ti��iW�Ū������P�@���Gƥr��]��򝿖
��4=&rnZ�����������Ow��	�a��u�RRK"����.1a� ���ʏu̥��5�Ю�U�6�*h(�M6+h�$�brD q�NP1����I(C�C�����l̀Z��0ݧ"�b��.�=��%��eKظ�^�g��V�;@z����ǥ���d���> ռA1�icՠ�v���s;b�'<�h4:p�I P�ĕNz���,��HҀ�-"���=m�i����E�U?e��A��;��`����إ(sX�섀�h���n�ywOӧ����h�vW��9{�W!�/�T��K_��Ic�d#���n.���| �� ����H��uR\��KJ`$�k��%Y��B,��)�h�!�F��b�<ݞě����^�y?�D4M�ZV�<��g����z�6ST	��䀭/���EJ�����5G �C�ۻt�xqEj�X��(R̠r.S
�v��]��G�vUw���Q�nXNWMv�m4io��v���#Q�7�Rn��v�Q�Hn�eJ�:���,C*$��	Ŋ��H��$� $��D���M�^��;c	���|}��2�yJ���l��N��%lKy��)�$�ՠ68X;�-��2yxgWl����v�C��Y��j���u������.���l���K�z�aPy�5����:��A��c0��������Q�2�-���U���eṄ0J�w��u�u鹻�W��Y|�J�	C3��߫r���U���4I��N�愪��"�i�"����m���aʐ��O�	i#�����I"�s�u	
.�3%�����{=�є�@�0�-�6�/u�)oaQU��V�~�^>$�[�њ���t��Q�3T���/l�<�HLI��&�y{c{�T֕�RT�?��Ye�J`�\F$�=�9
�g��j~����Qq3�:��:��ـUoe1���r7u�Kӭ��
�Ô�?�O՘NZ�D��Cq}�VJ��/��1�Z ��2�����z�\~�T�u�,Υ����'���F�~=��^��0�xPF���):��`6
�AP����O�XB'5� V�9l)������YG��������@�o�*�{0u�,Ċ��xj#/������%�G��R`����5�\����KM1ְ�i
Z�r.>�z�ך��*^S&��8�P���6��{�����K����gD�����76jI�����,���K�N4�<>�5�?({���]�̮%}��' �gO����P.BY��V/[�m� >������Q���q�&�[l1?�Z؉x�51?�3b[:��Vܭ�ch�R�~�u�C��>`����խG]/�hs#��ϯ�� j�����X�����kI� i8�EԂ,p5	�VU�NΚ���}e�e�9�7i�<�៹�5 |E�I���2Kfc�������3q��֗^(�ek3D�i__%�Qb.vSD����/ѿ{+V� ߶�6,��{!S�N�/|�j�ZrHN�'����c�-��+F
q$;�CP+�H5���;e�tU��pB����{C:s��s�����ֶmΑ!c�
v���q�gr���(���C̋�e��e�nM�'�qΤ��Ҟ�tG�~�A���DiDUGSE�?��ж���f�P�J������U4�q�Us1~4!�G���6d�Vvn|11	}�_~7��|�&�og̀᧯�$�7:}��|j������-*D�
P��#����r��?(����Ҟ�Ax�;��w��i�*R�� /F5Ѻ���T7�br�!a��n/l�LLa��3���`m9󟻌��'���cb�,jD���&y4i]{�K�����6L`�Kd�R���U#J�����Y�_/�1o��4JW�f��?��EϤ����h\r����+X�]G����:�0u�)p$�����>ۆ]��.1i��D�΀<$rPV��@�}n7M�ɾ?F��:?��oȮZ�W9���]�y���ƵR�Lʂ�E%��I��UDvx7٪ Q?m0�S��h�p
p
�!��K[�3<e��#�:�M�B��&��@2������Bh�;�f;\��n�±L����3��Dr�H�XGF��`[��s8Z	8�͕��󳤷h~I�w�|Ĵ#�x�����Z��{�yy���f�4���A��.����� �d���_w=�3Ǜ�l03�'�J -0�볂8��N/�G|�jj�!t�����	��#����G(�F["�8:m�s�	��4c���zl���7�i�W��!�V@w6b�� ß��鸛��b�~}�n���P�?q'���Ϗָ��|8����Ѻ˅E���K���dl�������s����j��wmj����k��;?�|����550���/J�.2E��q�Ӎ��"Qs�������,ƥ�N�m���sh���!�J;'�t�~.kĊ.?��˂�ېV���ɓ��wS�gd)I��M�î��R�^��;��pFRuy%�i�X9��0�cCy}
�M�����&C9�I�����x�w�'���6jO�b�1ֆ�gV����y�p�,�Bi]��B�7��~0�V��HEw�m]oa5�gX�v��r��+���g�����G ~�!�]G�sR�㻴��P�b�Ψ3'�>k�L3'K��@�ar�<�wPp�,��$�;�6�ZK>!f+m����b�Ni8f �<���Ԣ�)�3c?��-�ñ�N�G�X������T��X6m���������rN�����t<��I���b�q�-4���&����Z	�$w�S�,^��?�諮ISGF]w$f׈2/�6�SN�h���t)���!%�T�Yv�h�����;F��M4l��ʟ`(�Br�כ�����*�'9ڡ����6����������ob�����l���]P���T/��Y�<�!�GCF3�6�Y�mĩ5@���WZ^^?>k�����̬�tb.{I��������Z�+a<BǆC�O������^x|����Xr����P�m�}�{t�@��iM[r���'2������`�$�Vυ��R��*�g��^�z��'6��Kd���IHt{����%��D��M2u�Rt��SK��7���	"F���,�Û�S��^��O�XSDP�/��XL@�N?�b��ݵ��,�1+�RH��]2R�b�4�!���x�%�Zj��p��6ܫH�1(B�������K����0_�Xt�ꖲ�\�������ñ���9�ᚖs�p4C!(����|��Yp�q���<VCI��P\�)
HE	ǉQY
*�-.E�����Y�)�`O�W$��������,2���u��ux�R�AI�L]�Ie5�����fb|1:�I8 /�$��%��Ba 4�X�F@�������߫������谏PK�����#�* ��a��-(P�?���P���L���xɒ�).I�Z�*�n���)� ���aT)�B�ĘVϢ��(t�M�i�-�����.*�`��꓋�y��
Y�p`���E�}�]�Z�����t��ͣw&,bTw\�p��3�i�����a#��h��c�W��tQ�%]|�^?W�}��5c5����e�$)���uM��T�|xg;מ	�%Y�P+P6���(��7ze��/25$)<����m�{	�r�!7]���Y��f���J�i�X��9�л���&I�ƖT���\������n?���?�"��R�i�2f*۔+&Pj�t�@u��G��~��@ݨ-Z���a�W��4�̇�AWa����m��2��øV]\�+���e2⨔�q�ª޶ҡ(H��-c^�d�=1��2�����F�;~J�Tep\\M��bO2�8�^n�GQ�H�i��s����\h�n8���ι�Jxn�d��J�/��1���w�H�@��`��*�(q���z�U��}IT�h���&)�Qb��m3�*���ޙ�u���p?_x�kEA�!^� }�"�������ۜ���,�������	z+}�9��W��.3~S;J��Ү����hZ�:[��w�	��2�7k��7�1�<��rS%�4J�����Ui�..P��� �������a�8,�B4c��V���f���N� �I
��]s�Ʋ3mN �=#�*9G��F��!��2�z�� R�d�	<�]�S�{,P1SO���*�0 ��Y��,����2���lv�tj?�&��G�wH��%������?�\��uc�ٖa�s�$���e�t3���2z��\�(��o#/F��2��&b��<Ҏ�HQ����Tj7�B�K���u'��u�@c�+�{D��v �����-N�(�o��٪�[W�t�<3`��e��C+��@��9�����w=SC���T&�(���=7a ah����3�uk�=����L� ,��	#h+���2�tj��T�sg�Gۥ+�<Pإ���ԋC�D�"���uν��r��!K���At	�S�EH�x}�3�}���A�$d�*���ܾ]y���M�
ξ�BZ�	��zbqIb_��c����h��tk;��N��VK�~j;B���!N��Q~j�������ǈD
�˦�A�>z=�t��0m*�5�o˕�1����59u
hq�`]*}K�6OE?uJ�W��.���,3�05w7��97%^�EjL��69�mY0��@�uّ���s��.��������������6
A ��wWyޫ�P������bf��z�g�K�2g�
����D��F7b��_	��Z{�@1����fYJ����Ř)mjHs�QY�t9�dI��������&E���g�&�� ч�ĸkQ�G�CG
��w������"�}hO
2z$�{��M�3�M�n��
�=�<�A�|�QCe��l����_���晲����
���|Y�.A�&Lx�W�hTO�b���>O/'��F��p���Ԉ��7�C�'�x~��X�ߍ��,Z��c5��|�g��ܛ����*������� �X0:i"y�X���J�$2'��5(8?����.����G�Su^�p�Є��ӛ٫,�3���������%[s����eQ�_�F:)��Lʖ�A�ڂJR)C\��U�w��=3D��]Z��c�F?7����H4 KJ�r@���̄�lZ&gꉤ���.�:j���@��QdC�ۃ��5z$��Q?1d��y-�Z�Y?o#���6�M�oz�k��c��bK۷�zBү��4��7F�F�w�C� ӱ��:R�������1f�E���~#�ER��"\����/���Wi�-$R�̓�-���_aŌLD������[@[���X7b{0���Od��jo9Nt�=f�
��K�H5�C���U��Q�K#�#@���a�b�+����֒�R1�4UFqr�'�EU�T�|M�#6	����7����{�%6�+¯y�T�ף9�{Ć��~�̖m��^����`y��x�C��1{hLn��>j����WX6�M?�b3S����0�*�"��Q��9¥����ū��xKBYp����p,E��JRb�SGܸ>|ӝ˂@;Mv�~ ��^�p�@����8*�T5ӗW�\��W���9�K�qS�^�&�P�rB��͝��6���,����J%�W�-�?$����#��J���"�_O2`2[)�����f��V�K�7��S��r|f��C�7�]��T�����E6�UVi�xJ��'g�±)���p�z�/��]�x��h̦�bR�U߫3� ���AQ�ݿ���X�+�֟ܜ������v���tl�����~��9��P%+p�C����OTB� ��(�����4~Dv�����W_PQ�ܜ��dCߎxI�A"]��7��)9��k;�	h�v>�x"�uL���_�B6����&&� '�^��6���B
mƒ YJ����$n�)3���N��49x������ՋHcne�b��4�1�\;��k�/��ݻ�����J4����{W2�6�������C�e���$hJ�135��s�Ҩ4, �F�����sz�o�=�5�c�b��{rM���T�{×�rt�۱����D>�Ǜ�kXY�ɭ��]�$&�*m�S�-�y���h/�_M�O��:�߄�B0��7�M
ђ��M��]l���z���Uފ~C��S&R��!M��~I�P�f���C#�Ը ��`qhJ�p�����2��N���l\Õ� E����̩�gى���#�����uq�%��	u�&���r�)�%�Z<dʠA���e~���ǵ=��B���ҍ:he�7�/�����@�q����c6$ٻ�Q�S;�k !���B<�v�s�cwiY<�bN&�hi���5_-��S��s��ުn�S��W��klS�!�S���㋓��n����jYC�V����'d��W�ܷ���֔���f��[=�E�}go>�6����/���Z���4��2�aK��M��
�u�n�r��J���WIRC.�'b���t8~��~(�V�t�=���Ls�!���M�����=�gV�M`����XOK�	k�hI���8z�3��*}L�e%��['�HF���|��*��	tH4g��v�Nu�)(+�w֪�d	�����������N�z*�lp��j�[�� ����������C�;9eg�b<֚��J�G4� +��v����,XF��$�Po�[�ih���'�qX��9Bܼ�� _y,_x�%2!ʝ������pH9�r�D-7UD^���^W{?F��;W�dHR֏�� �1l�>3:�j�8�K�S(R�8�KW�=Ⴜ��B�d�9M���l�E�C�9�c���S�i��cv:��Z�?�M�vBC_�4��hB/H��k#v�d��ఒz��q s �Q,�-���e:�h֠���8Ĭϝ��xǦ�~9��0���)"��I��o��8hm#��%Xu�aBG�\}XS���XJ�ʿ��վ�v���	h!<.�ubfu���~�f�s�S1��RT�v�n��.A:]�:dt:�N��\O���$똆Hc+�<��2���-��~k�Dw�l6��1��v���ohFE�����c�y�RN1,��(�U;LN�{֘��4�j��ؗ$��AQPU��w�A�$4*�d�E}�o;N�L��HD�>��W���~��}��a0ZVk7"ug�ZZ�B��E���4I;ꔧ��O�����p���Ix����u�e[h;� H�C��\��ݦ�����~�j�Yx�]�Ƀ�#U�)��p���[���;��y5��ȟf`"_��2���偭d m �|@Sү%�;MO���)�U�=��܎ZW����fx.|�#j~�A���'S�x�C�_R��d��+�/4�pRzQ�!��H/�;��;��|7���ٿ��f%��z��P���4���=䇇f���}z6o���ȹ��cçQ�F��~)N*����|��ux�~�ӑ-k�	����u�h&! �
�{��>�g`���=�r�hl���W�N��,�ʣ�����7S�!���D،��c��LE�����m��
�	�{���jy�HlW�Y�����B�	q��8t���FK��l��4rf��g�)x��u-�o�&��O9�ƃ���q���L����;IIک��O����!dn'��.9����]������#�y}eĹK���"�t�E����F��#�ɏ�g���lJ��0r��9+��W�v��o���B�]�&�S'�2-%J�Y��������DbP9X����~Bf�a{��r�A���K�����8��K8 (ԤT�[��xbH����j�����LB��Ʒa�uշ�H
d�g����}Q�S�h�|�O��~���ӄ
m}���]*���K��#�lǅw�d	���y���zsㆭ���p|��%�D�������� ~���(z�_��d K�+�����h�<W�57�<�I�C�����
[�E�Y�j(յMg�|S�~78U�[��$u�Yl'^��E�Q+�R0�oG��T����H�J^s�4K{���
e1���'�ɔԾS���taն��C��� ᐈ7r�R⺤�䠽 VE��#⡒�
Xi���������DR��"�V�sM� ��W�ǁ��r��U/�T�9ُ�&���D�F|^l�T����A���y �.�=�c!��"�~��_�� �c߮^���ܑi�)�%� p�%S��؄��@7�Ğ~��a2��z���S5���§c�0d7}C֫A-LZ�h��T���9J�}a��נ}jq{�7����t\Sa ���g���r���`$��OOc�f��;���N�x������|��[K� �[��K���zӾ����k}�0��u=��p�FP�y3���7�����VD���L f�,[斴��M�����*<6�"�w{v&�"X!�bD ����u�ǈ@������>��ks�N9��:L_+KBz\���l���՘���)�W��	�7��~�A���/[A|�4r�nXI�\6������{��^~&ى��ó��`^�g~�ܿ�5��k�k�8t�%�.8� O�p�
<��&�b/m=5��C�"��z����Sxe�I�޻ub$�8�����޷d[?���#�� ���Z�%r:%��?�i�T^5���s�AM�¾�q>���� ��iE�'�qH}TX`�"ud��V��R�}�9\^�g�� ��9"\���&$� Jk�B��e"C��,�q9V��S}c��^:�=����Pr���)�������)"�-�,�rU�`�Ҽa�,�,���-�1��@=��B��?(�{f�V�8�T=�/W�6���\��@��zp�:�(���#J�����-Fa{t�I�GxR����Ê��P�G�h�������K�҉-
���-�W�@��-d�z��ě�R�@�7ꇍ�� "��^#�h���U����{�0[���-wF��C5VX1�h����j�y����@$6���r�aA̡CE'��7I�����X�:�g�j�u�����ǽRv�J�S��X8�E7d�.�J���G�zE[�����3��r����5���e��)��W>'H��F��"Rk��xO��	� ���[��/�9�3L�x��<�~�y���R�S<:����� ��L��=e`��(�GZ1Q���i/�+fV	_�'�:���8�,�������:�/.���n&�Z@O��#5��'��r9����;DƜ�v��=�����к8y^�3z��,"��oS����Y.����:�W�|Sw��ʶ��Ɔ��P>�0i��o:ю8ܺy�a�k�p�7�9@�!yq���u���O�b��!5�u�Tl�D�-��S�G�uA�ص�}�@��sV�[�ר6,���W"��ꠡSfu�����$ �Ƃ����U;ۏ#���[ly�$	��)�bf:�l�9ٕ�Ht�/�2��ǣǽ�6�� �R,ޭ�z�F.�GQ� 2EmK����頽�|�����FM�~w~����1�t�"�Y|�v�ςT!�E%�ui�Ƣ���
�AqB��'��!�TQ�jC���ckC��xvu�:�=L�J�`�{��>��6d��*�xכ�$��<�wD��ɡ��sL'G��sC-څZ����1��������>�1N*�C�c�ʨ*b%X5y�s��]7E�z���\`��~i�9��w#T-f� ԄK�Hg	v/��[1M��L��+�a2��k2���I"�-�������&7M���;�DK��i�%�MG)��"�g��6�*�{Z�A����Vަ`��w��~+�l������|ʼ{��'���Ŵu^ZAɆ��]ȯ���9��X�&ԟ�m��^�>�m�%!K��D��ăv�������6����9�yh������D��@� -����{A�v1õ�@��>�,(8�}��=[`;Wn������Ә>R��~�_Q�iJ���� ��dY� �|�����\�׀{N�D�D}g�06��~p�f@�*��K�������r�.��(2�@�<�1~w��֦�N�T��9�͚aqr���	6E,�<����~�)L>����Bƛo=���>�ЗM�%!�접BT|խadFdh�5�F�[�G�D:"����Dٿe�\����а�����YL|��Ot����0�Q�7JP�W��A�.Vո�[aþ�d�v?~�d�8(�O
%��6�S7Jk.�&�������["9�mӄn�bN��'4�����<L9�X�*1�u0�+OŐ��52��o[`�&�x�vE�������{T&���y�'�1֘Э>�\ �����;'9u�ǺU�|����?b���k��'X��.�� &p���8;�-�c�r��m� ��)�L�/׶0�C����*��n���h«!�Qe�B���P;���7�<nʗ��,]���C�,�:6�U!v$�e�+��n�)��@� ��N���ŷ#`R�ne3����6��ƪ�^n'>�p���j�Č���hg��L�}���Q�Qdέ!_���Pէ1���kS(ҎK�t�qx�Ѵ�L����^�S
CZH���.��8n��a�y-u��`Hv��q���"?vJe|
�m��'�#�5,_�a����L���W�b��C�ψ������6��iQ%�-� 1���i]�'�m�E������)�$ӝ|����w�,�c�yJ�r=�\=�p؄�C�MM��`p2�H&�]�qUs�d��\D�7��0����Ԋ���/d�C�t�t�f�W��Cs�Ź�	rn�]S=�Vn�)�"%�s@$S�L�ZJ���զ�k���4�Q�/�~1'���j��Q�󽓆˦�óCQ��!��f���a�Ve����X���M~�[/@'�Q�T)>*�U�_�-ģ�|=,���j�7�eҝ�wKO'��oυph�Q&�O;ҭ��(q=2��ϳ��W�����3���}�������pM����H�f��n RN~kt������2�B��<�q���`��yղg�ɗjq������q[�P#iӾ�Eg3���lŌ)�?�$l��V�04e�B��O� X�t�T-����}�F9-��߆��=?����H��@����� XpȀ̄G��=Z��xYFU�^��q$m��8&
J>r�L!2歡`�(����������G|\=���8��3u��I�P-�Ι�����@D_�s���v�(�Tn�da��,LQvr��BX�4���/O�5[���)�9{���c���1��e)a�&e<w�}2��A�-�y��1M}�Q��=Lh�SƉ�g��q�k�A$LoW��n���:/��1� 8Y�8y��-�x�.�Lv���Z�Ry�������mu��J��0Ҡ2�.�����љ谗ᡤS"bF���+�/���ݹW��2��,������P�t�m�mƻ툭������@��ʷv�h#��P���O�z1��ݚ�Ԭ@X_О ���Rj�S��A��FLR �6+��)K����b�C�����`p�愸q,����zpv�i&tѰ�K�[do��K���z�ڭ���r]{k15P���A�Ś�E ��q�O�*��
�f5�U�NvE0��B/���"E�d���� �P���1�/�#;$6҈t�_oèM>�&�e
$W��"�k.vU �������o�3��PZʅiQ>�>����$E�ֹ{爨˨�q�,��,�-�-M����c��h�*Fpi�P�������[�1�׉��y�<�9W�_����&1nXv��৥�7�*P�����
Z�K5ﱑ�yPi��O����}-	,:�^�<W3�sX����,�ej��n^�R�グ~������)
5��!ɓ�R ͝+P�t�kh}��%��탼�W�@�����U�^	������Jc�񸦘iJj�6��;��S�׹�W��B�̻��4mb��t����g�n�i�H�qLE>�jG��܈(��,<�z��I���'�L�<���}��5Q���HM�I�����A�ƔF�$J�����D]��p��k��H���_��:�J���'��I��Aq/�7��p~��_�4�پ|�gO<7E��zw��{�Ki����:��\�Dr�<�]�_�V��D�O��f��c��97��g=���~Q/&��竊�A&|�@�>Df�h+��[�@�1��L��l�0�W���2ЉL��U��1d��@���U�wF��}���U�v�:�n������ڤ��׷�5�	`(;�7�6V����V�ބ����j-=g}�@���2Z )X<�:�c�}�u2P{����aT񐊜7w�^֗G"�=p�TV���5Dȳ���1�nOnGK�U�V=��(���V���.�-�l��B~�85�_F��+q��Ì"L`?���IeN����m>��h=�;6Ж�9��o�7*��6�LĄ��ȴ�-���^d�m�+K�G����������i:	g�%4��З�2��{7s�j� C��0`�)cE�u��+$e�}cŀ5	���s��;�,��E�l70^���dAc@)�F|h���Z���%`��^xZ��H���艦q� �^�l�� 3���?����|`Bٻ������r��I��gT�����%���dc�(��T�+�ѧ�ܿ1c�tB
�8��B���"x�a��:3��_���62Ё�h���6�4f�-o+��/��`[�X�h�D�OU9���ژ6�3�t`��X��k���W	EH��ب��i��͠�� [{�{���Y���gi����ϐNޞ�^o$qp`.��w�V?b����0�c>X�t�&���S׉�l�*�$(Z�>�\�D�|�$�����%Ƈ x���$����Ǐ-��h�.g�P�E럆Ė�>Y7��鄷r\������8�.<�8-w�w��1[?=�0u�rf����_���I�ŰS6(8v\`�15��nܤ�΀oF��H;��P�[���l�>b��?�+go'���X�ݢ�l��<��-<?��+0J��V}p�^�kQ p�+��yIĸ�ţTI$>Z�|d���AǢ
/��� H~���.�,B9�Vo��B�����5ރ����H��Z��mc&JU[��?f<Ed�V�?|���#���aU�4��=�t���=7t�:��r���%jb�k 2�s�_Cwh�q7�ު�\l�e��93!ݗ8�1�cs����u	2@��ЉSI�ַ�>T<���ۿI~7�!�yP	�3��%�q3�{�)Y�Y���3�t5�|�~�T-3r�:M/���Q��nB�M�n�n
}��D�F�����	Θ}<�y&lV�����j�<���r�H��(�؋-}�$�t�`p�S��Ε���I-�[2:pZư��y�x�@�ޢ�(�{�mI��iōF�ުR�t�'�S��+�v���%�`8N)�;�iv-:{-���JO���}��ʋ������o�19R�t����j4i��^	!�C ������9WwA�_�@L�nWR�ɥ�3@j�D۸r�-���Ѐ�dS|���p���(
޶�[P/؁�u?E�,�>>��բ>��ǈ%+� �׼1�jzb䓥> 5���_'g�<SL�Q]���!��&�.��K�yZ��v0Y��zb9�����H�e\=��i�Y&�ryO�8	Ƚ���U���H��ShLvk��9��,joE"�[��I��<��. ���`]��cp�$@?�k0c��OJM�!��Hԭ�b��a�5)zF䀿�M
|Y����l���2)��r;�"�1�ۀ�	���1%�VY��p��7��$�C� �7����t5��yY�^t5��x��A�݂+����T�7 �=�2G�3�*�Z�QFˈ|>�e�gO�=�7HX���35����t��A�������U͏)�҉�̔!��u0/p�9��t.�)����Ht���s�XL�6�ux'׾P�U�_�9����Qˤ�PD�����n�-}MB �0wY��D<����Jf<��jT��w�JQӛ� �=F�B5�m�����L0�,�7i:B="d/�q�o|aժ,���&Ih�pІ��dv��,�ɞ�ԟ��љ�D�����E�|u�΢�Oi�*�6)(~��a]C�/��-�$�E��x�?��Ph=���kɱFJQ��r�}��*b�V�(1�Q���T]�~���Y��N5 Տ��n�sXk���Ck�3ߗ�r��Ub��%|��#D��ܚ������:Ge���*^0z��]���Ͽ�8��j�L�#u���RbvC���=(�
�%J�C\w��^q�?�������}��S"�[�e*Bz>���oq��w+S�W��EtC4���L�� �.��`������檰���:w��bv#��P�:]�p &^j8fȋL'�珵�a�3p������x5���s�~@l��R�N6��h�y�kL���2��AZY��gJƲ�Kd��|A��jl=6�`���|ot�N�GpDT3u)6��!�l�ZY��w�5�����0��\9���P�]D��<���qsS�W	�D�%�i� ��K���)ֽ}T�U�н~�i�O?+w�9zT�j�L�T�	r��[��4�3:Nz������ߗ��$��Fp�	��̀�ѧ
A���ݫ��~�3�/����Z:���M}@ә�Odܞ��<S&Z��=�u�&O0ӄ��c���k8��S�A�G���p�Wu�P���LD�}���vN�7Q�"��_�D&���D���������ePqI	H@��vsþ�5�i�T띕���	�;��w�B)�`A`�8e?�e��2׾<���h�qD��j��p�#f_ՎqyLLZ����ւ
7��VYq`q'2a	@(M"6�ʬ{K��%'�e-6-��W����^3��(Pأ�⿈�K����2�'i�;���3n�R�N���x�q&;I���}�)}�ꗡW�XlB4�i�F����,B֞�K���<��y.�����$�����3�F�?�F�=���q��~��E�^6[^��hy>;9cY�d���P�\�Eh5�����g�3=����X��J�B���Œq��oaCn'�H[e��A���`B��l��h��	��u|T�Pc:���_c{X�����1��[�d�t���E$���(gNE�]h+�Q<�V!$�֏z�	%�Y ��>�Cj���"�l?j&��p�a?TnV��u�6�e��~>A
r,`��N=�r�����P/��}�pNv0�;0�@@@�]��8����ڒKC�gkTE�b��3~�xV�u-/����a�a?�}�����{ff��](n\G�]��]�Hac���dߧ}ӌ���=;I��=��"v��"H,
ăo@*����N%)Gq��O$G\��U��3>/5�z��߻[���@���j�[���8M�T�I�s�qYGꝒ$��`Ș��h�z�b��%���nʐ)+jG$�Ϳ1��/��u4+�������LC��6ѿ�Vǝh?�_�5�Za�i�����s�?rlq�x�-T{�x��ొ�(/���U=�vb�B2:�$�;J��)E�[�+%B�4lv�[q�`&1��+9J�r"�N�.K�{{r]ͯ?*�=+�֐b��wώ�6��r,m��w6�9b�7�8p�G>(�B�3�bt�j%�
�RMξ���~4A{�5TT����]�.)�2��O���(���Ʋ�U���y�\X* ��2�Z�����I�-no�gؼyW1{��)��ܽUނf���Ƶ�H)R3�Y\Ǡk�B��hQM]j+};fw*k��D�/vo ���ci�](>�Y𰋐��sG崮��̞�[�y�:��4�pS<
�I�6c��;�(	�x�j��#Ig�Gdƍ9��n)i�!&��Ʃ�lu*�Q�R���h&��k����1P=����=wb�����}kb{��ɜ-j$��:3�0���$��P�-���E
]7����v<�+���TO�A��nZ乎E>�&c��>�� v����r��B�]���6��"��ݜJţ���Z �
����D9�����o��1
��U��S^s[ռ��5��L�M�YzI�6����]X^`��	
i���]ɖ���(�H"�2��}?�T�����<�S�U[k9����w�ZtE��Ӏ��{�`2Ey5 ���Q󹝫�1�l�Tq�D?Q%LV%+���~�(�6!��]���xl�����"ڇ7NJ�^,]�b#vx�ђ$�ۘ�w�?J%����������-4��A:N�������>!��b�y���_�W�/�����Բ��N�)���}vO/���
pr�ω�c̗E7��}AJ�#7¸�C��:���ވt�k��+u-�7f����9������<�`�\�N���8le4�T�M|���,\���s�q�ʴIE��b\�a����^X�z���7��{eO�뇘.�f%�50pܹ%�<���z��C���ߞ'<�G.ns`A�u+���(g�u���S!} Fw6��r8U�T�o�+[?�
��_6�� ��Ʈ�%ū�/n����};̀�E�{�lR�}���
{e��������t��|�L���qaB(�KOʻ?����}p�7�!��I�˶�s��!zLa��*�d��.����{�Lr��y㕉wr���v���Ho��L} ����SN�g��f���u���a�/���c�tGz��;���Y+����� �_�&c�E{���&�6�$�֦�I]��W��j�*"����=�~��
-��E��`LC��7)���ukgn �a�~)�!J(�drE��1�j�Q�+pם�:4� �_PU��&����)�,�{�j��p~1�M�k�<�e;l�ߊ��ot�}u�\�aTI�9nQ��`&k�3p�gw��x�nR7N�;%�&p�G�=M�16o���{�BҽA���A$ǫ�]��,ٜ�t���% �P,�G�Phx��籇Q�C�]�@������1�i�����Fn=��|�x����dH�/�6��N���x����9c[��� ������j�ș��R� ��S�,��y��-d̄ ��J9�]���:F�������}��^���W1�j�i�%�}jU6
�Ĕ�&F<�qƈ�l��	.P��G^�B�`kء=�)�xm[�8qC��[�7�v�����)=�,�a�@��^�b�y�����DN.�'����;8U�Sy��|�5Io��hy��>{�P���i蛫pң��t�A^u	]�8�������4�u8���e�x+ነ/4�<�
ڔ�@�|8�)Μ�����1q?���ƽup�]��e�������o�,�J�D=Dඓ��^��\�D8@�M�w0M�5��dT��(��s�d�)]�6��*a�)�Զ�'��w�&(�#=Z�?n��ı����MΞ��m�Fp�#yw�8�X��b��@���8�����xF����OQ�T}(�2�+���ԯAֽ~�F<��o��=�ŷK�L��y���,mn��	b����pЫvJg����0�������8D��.�����g�S� �I�o.�Q�2L)d0��/��W�f �f�-4n H
/'�[�_��j�'_yJ�Ϟ�}��\A���+IS��?+�Cݓm"�봮1P�8u������%�
�=xZ�@�d����o�vv(��q��T ��5�yS���8�]����Gr��@���߯�[G�w��mk�e�NŐ�oQ��] �9��������� !�u�	���(�����;�~��j��G#���IG[y�+���Oy�}�Υ�9���U'6�k�v.�������Ո\��J�gpP�hU�X8������,���Y�f�;|��͌d����说n��B|R �d��x��?���pi����G�w��Lf�0����غ�.ͷ{�B��`�:�BN��,LK]��ŷPV�~�'nGD����[�����Qe���_�r�n�jHh+^Fl#�4Kzh�
�܍�ix��� )&�=y�����>���O����U���s�E��n�8<JW���A
�H�;�S��V �r��ɡL��/K}�3Tr��C?3o�6=xm���eT���&���CIS)�v�z��dCWԣ�JU��Vǚ�YҰuH�e�S|+_gßa��0pY��xiް�t&2���g^�0Pb�t�\_��+������¹�FM�F�/��C,"���5}G�ԩ�� �B�k��܌��KYcHI&P|;|R�� ��np���_�������������*�$�%}s����q��~��32bD�F��3��l*�7R�����r�$Gx-!inR��l��_h�G�\{"N��+�������J��1�C�wJH3�_-k����t�� ��~� ���4�.���g�h��{��$�/j;|1dZ��6|&$�kr[q�*[4�?��8z�_6���Xc��2�| ҏ�vϩyt�^c��jP��3a�E�x��?��#�ً��s�sᶊ���/͛ˉ�Y߬��^�����j�pS�Ypx�A��AP�F��_�!����$�͒���'�b���7~ڞ2)�A�#d���s�_^2�d���O�J���w�)��)�D�0��N0��{���S��?�3�?M���wS#?|Y���_�Ҿ�TP��/KdjDƼ#ޫ�9)F�À6̝�] �;��*�\������^uW�IX�b���
Yɼ��m0-B̸���tC�:>Wb��cn�=*6�]E�n̔�q��)$�KHK\����\q������6z)1z�6d$6�y�,��vZ�-2�n��L�]��xt3q$�gO�{����9��jAYw�wHm&��
�CZ�m��K�N�t
2��2�)�#}� �F����cM�t��BY% ��3��P��:�L�$����&&2"4'�������z%�DH�a���b�-�'-��Z�԰�2[�EY}S(��7�<P�o���|U�&��[��ı�������V�ϕ���N]�
�HB�9Σ{pބU�1a;6p2TC�u���XW�� )W}�FM]ښg�*:�n�4}ԼD6]L�G
L�wI�˿}X�R���D�df���>�⠔[M��<%��9jQ��m8��Ɔn�� ��R�5(eǷos,�X&���eƤ�E�t=i+i��zD�����u��/���fd/BO�wr9�S������_���BE�x*�ph/��)���ԭ!���0nąM�ދ�[иX;3�Nh�����U{>{�H���h?�qtC�<NR����a�o�?՗�f-�:��d�㈻�T�=��P��~d��P6),V����A����r+�@���"�1�䘴P��l��
�R}������'��W����. �^��yj��A�F��I�	\(Ujm�����Œ@�ˤ#
]U!ٳ��]��DQ�'#�]1�-��J+��Zr_{�$eg��֧ϱ���s�{$_���H1���9&oڴ`�N�OC����;uoYC�lT������A�RYqJ���� �a/�A�L���G�D�H%)M:���?B}��w�
�c��_��e}D���y�O�h6���?��7&I��5�,�m�?X��I���}��aS���� �pz�Nn�#�`~��0�3��9!����.6^���5��f��$s$�DB_�}�I�N喧����\O�]�CE���H��I_�.���&?��;�Q�y�{q�
����#�c��mAU1>�.���VD�?w'�_6���.�T�$�^m��o}�-��[��ȸ}^u���`L}A�#�f;�;����
AD�n����3�%��}�e��]�C�XOD���W��̮����iJ7����C*oj��<aؑa�2a1pPh��ȧ\��*��@۬ ���pD[b�=�9�6�m�0��[�rP��fd
j�B�jmHn����5��R�;Ʈ�&�H�0s�{u��Ogh4��u�-8e$<x�]l� ��nY�� �(kq��	��F@U��j)0T.�8�H*�	��ohSYKS'�M�K�%��Vu�b}0/����	�ti��։N��E�G�n&@�EVd�6*�V��dU3���l���#H9bA�z��T�C���qWZ�?!�i�$jAc���m�&E�}�L�]�C�d� �e5k���C������k=jSf�@�
�PF]�%R�mf�C���y�y(#5d�3�o�'J�r���U\j�����Y����`��i�tr�E�"d�K������'A��/��f��K�S$�0���ݧ�u��8�z��ܿ������n�.ͤt	}�.|;Ed�/]���J	����c�^��ί�l��@��|V�<�ua�k����Ѝ�I��b�z,�݄WYѠț>^��pB�I�Њ5��Oh0	*�i1��/�����:Q����4���YoK`tO��B!8�V���&�F���P���N��;l�z1��}�:��b�+nyW+;��S�Ma	�us�l�n1҆ނ���/fv��%W��o5�r;s��e�
��mP��%��ؖ��s��S����d�JX��+�n��f�T��Ƈ[ �8�}����T�~FN�C�r�DW��ECo���|���8K��N{�J��� �k�u����$ |0�F�iƝ�h��?�ˀQ��^r���J��[n�Ȫq!�u0#�s��[3!n �"��B�;R7_�h>D�����'�����[���Bf'�vv=1�љU9��Y�S�쌊:�5θ��U�1p�u��_��� `��������A�Qw�]/RȥVa@�$�/�S�$%v%�O��ʛ}���b���k��t�HL�/cyW�O�l�"���2��&';�0u[S�߄Fۋn�O�`,{��~��ξ�/ "�	āoQ�j��C�+��}�d����{���4��@�dvF�X�����G,Y>�NЁ�E��*�Lw��"�3F!�l�x���]�����{+�I�"��'�T}�����[�d��W�����;�Պ�� S����\=������u���1�����7���n}�f����㟚�,�f-�}�U)�g壀C���m�K4�u��5f�DH[��~F@O1fM�'8����O��Қ�X{�uU};S72����Q�������7;�qm0�Q�썈��ĩlf�alF]�Ha��/�[#ކ�.��I�I�)���"�����/jMq톯�l	x�DS���o+a��{U/
l�mҎ��ć��W߷�&�.ҎC�V"U��WeC	^�Ӓ�"��u^�ю�8)3;w��џ[��cn5��ch�#s�����n�1�������gO�~���hy�4�Yn�As]3�l92�s�@�1�w��0�p�@D	��!ܥ�ر�3�����4<�+u���ߛUz�R�/�5�ٖ�h��U�{��]8GZ*�b5p�sNb��L� A�����|��u���Z4M	8+y,��Nj�.���j�'� ���p���ƿ���.i%_l{p�A�� ݢ�M��j�8PKC�Y�`�)��*�l���W4'>$��
�d��d�5���ut�T۱���<f��zߋ�ow���ڱt}�R��q~8��o2�Y+|k��hO�7�G��iD�	��b9��p�Д_ �;Vf���@�f�t�^Z�(�w��t�
��f�i��4�3���}[��JM�ք>��k;��	����z��*�isӅ�qT��͑���p�������@��r���^\��nz�`7�2�vÆ�	�0FI=d1���F�H����ˉPl����L�=0f�h�s�����X+? 1sC� �p����"�O�*�K�˱��<3���iH,�њ`��2���})D�7j��u9O�<d���qy�'�W�a��칐]A�N��j�M9����9�[��R�'�������E��B���rfͼ��:�[�I\�x�u���,UF�X�	�C ��;���2��sF�Mh�w͖�qN�0�T�=H��K�J�I���'���,;y�W�-A���&��ˏ����<(�(sMc��3���HM#��$����Uml?_�U���_�Wpl'=��$lb�oN����G��ib��UZ�%�ǮA����6�gt��v�w��^��"� "/n`�sR�
w��d3H!J�`G���l�]S��|[5I����`!�"pMv,D�R�8��?+���V�=Q#	)�ЌGnJ�K,<����z��y�?2֔E��!Ju��,��o%�^��m�'�5�<^�z�������|�U
���lyz4<���J_��hŷ���MC}mX���йp�B�x�֡xHN��'�c"��)� ��h���H-\n��z�k��{y����)7�=���f�:H��npz�-�,v��SQ~s�t{>h�i~��'��T�h��_&�?�� ��?��-ٔ�TǑ�������Bn�3���m�l5�K�A?O��?zd��r�IoM�|I�#����y��Z����.�o��mb��+�0(��":e��N?���ʺȾ�@�5�*�Tx��$z���\B�����M�Ɂ�g~&��� ֡Qp�u���$�hF,=w!�Mc��2[�[��|~�2s�b�W�����4X�'�$��<ar����q�ab�Ɉ��Ǡ&1��HdT�ƷՋ�����GG�xF��H�l\�+Č��-���K@��Y�,�P�S������2�k[|r#����	`i)���u���+kA+�����$�j���c�z���)�Ew9�P����G�hM�V,\5/3+Ҷ��U�o���{Y�"B)�6)R��*�$��]�}SP��@�h�%Ɂ�I����#)�t���Ҥ�1
(�!�ܳ�<��y%�M�P��>�s�͟Ip���XaB�r"��Q!gϹ�΃�������pA>^���V��DF�,��q��9��^�5�-X��4���I���px�/�'�:�!���,#��OӑM��}��aI����T�EKQ�=��zǖ9�#_�u��[	҄n���'T�-caM����H�u���5�^�����¬{?{g�PI�#�)�tk?��wS��L��GUs%ñ���Aj�-��Jch��:/�K�lI��C؃`B�I�7���lΗc� ����AY����4�Rj�$w�c�\��$�m�功��p���?�Q�D���򍭗�]#5����#vD^˰��R_j%��[6%ݻ�H>?;�Դ���ᝑW����@�6=JF��?�Oއx�[�2wg�ť]S���M����&�F�� �,H�BY�ĦuWV�*3d�ᵇ�OP�<#�@����#\M^��<9������Z�I�!3࣌yz�K��ߺ��Ep�7�In����Ottd���S��������RY�S��7p�YW�ō8����*MI��?��I'l3)�����Z��y6��U�v=�ujD���Aw�ũ'�ǳDl����'CcjJ���`ݗf�=#��$�f,��{W���T=g��^5�K�l ��xG`Q�y���'_W�b�?�Ruqn���3H�M�TTyu����n�O@����$�F'�X��0H��xȭh�Ƞw����V�y�7�y��qm���i|�{��`p������+|;�Ѭ�L�eg����kf5�K�#�X���+�.�{`��^���,�{�[XyQo/�ۋ#!��*{�Ҫv�de�r����I 8���w����sg����-��6������nف��i���8<�ny8vFB!Q ��h7�ѹ�L:��^���irF��rJ�������'����1v���tk`*T��(�u:U+x�tƚo�`�Y�;:�NP���t�] ���UW��*T�����e#@o��A�ȆT���V����]�/2V�����2�)�y��� ��ļ�nbl5J= 8�<mגEP��;e]�L�#��MN0�;����y��b�݋2�"iC�Dp��+�
��:��Լ\�B��YԊw,dH���<�b����@�9��$��4�@w���@,D��=ڇ�;��[�EF���p��V�d.�щ��p�C��^Ϯ�T=T���W�	�-���!�u��$x��!.�'��g����-'���"m/m9�V��EC�\�Kd�rn��V�L�T��D���$S'	'��*�%)�u��@�_���y ���� �k������(��̅5�k�1ZI��&4}��;�:��v�Z�l<�Y�;�%q��`����ͷQٵ_lb���� M�ǿ��8�D�_\&H�a0�:���������?%��l�&��tIM,���x�OU<�8ek���2��������9ĤK�D�t[F�|�������S��3}5ʓu���xA
�r�1hR��-|��/&o�����ʩ?�^�=�����ģ��F�B���a?48��r��^�̴;�j�`���� ����d�͠F":E�|pME��K�vӣU���W�*��uoW:�rF��`�1�zԄ�F��R�Q%�0��!�CT��	Gp.Zj���1%"?�^&툣�Y���VյA%}����Y���vW}1`�3
�{��o{�`U���	�������َ�?�t%��+#����Eoe� wS�rY���ėa�|��d�_8�<����:���On�$��yF���eZ��_��C�H��-w���Շ��iP��M�_Jo�k#8w#޺v}��$�k(�@F��(��O�І�Fw�S;�V��I+&VEd��"R��n?Ev�E�&�T1ؗ��^ؿ͹��G�|uMc�<lU�g�����:�����Ŵ�5닢���WrQ�re�z-�+?�n�#��p�VcYq�d��K��<�e�B~'����HX�6�%9|5����N����M��u���A�7�8S	l���)��0���~/'�di�ߌe䍙�������?���˫mn8IOC���(�A�$������*{ȆV�.��ٌҼ#��_�*Ba3��崦�,�b��B_�O�Uh�iשqD3�P���6�~����L�$��2���}��w�E��Aά�6#���J}]���>��H>��Ͳpm��ү��ބ���q���Fqj)�C*���v��Y4^��mZ��m��V�r�F�"cƄ�pUtz�G��^�X�VWjh^I~�x� ?��Z"XU2��2�0�!�u/�Iw�����_^���тAT��V������	������o�t���QJ�%�*|f���?"e�#;��&wo{i�$������K��$�� �1t������<~b�B�3L�h��!������)�ch�.���\�7�7Sj��T��qU"����[܆���7{I�I)4 ] ��aT%����(�gF9i�W�4�E�8�ZG�E<�T��k��W�L|��	ED���u�#��;n3ͤ�P�0�~��z7i�ħ>�"g���W�c�)
:�һv�.��ؤH���Z3�����̣|0wqG��h�����0���!.�ZRHt����3���/�s�#�a��<Lw���#pa
�} �dG�ۑ?�)�(
�'�?8M�kP�d�89R�w�nq@��yeR.���v���~����S8���k=i�A�`�:��M�\��f�/�!w� ��"����Ԕk[g��Y�^pm�v�SA�B@����0�i�#�����Ir*�)��U��LH�f�Z�o`�Ro��n� l}�!T�	����Z����%#ƊlL��m����Z��}JJT���z?�ޣx���Fcf�}�@5
Y�Z�&��M�ؾz�X�"�?mjR2����u	%u���#u"\���9/�b���i�''N=��&P�J"������_@͞��N�l3"�/N^݌VL�p����,Q����8�#�_��7��~((��V�(��S�9��! A�(�F�U��i-n��˽�(��j��V�t)���2 m1{��:y㣮�iSx���p6w,��/=��g2s��̹3��+��2L�6?� r2����B�-mGʎ��P�ZiuGYd�Z������2��pE�u��B�R1k���9�C+ׁ�����8�F�\]}�+������k��<��-���%�ϔ���d��D��t�BE�m�6�O-Z��k�v82/b�YP_����Щ.< k�����Rí�գL��漸�x^Pi�ͳCg
�8=!Y?�%��y`�&4@��'W�F
>mbʲ��a`>��@�θ��x۠b��9V�L��F��-�(��`���xp�!5�G�s4-`^����e����|�J�s4EGG�<f�l}��{��E�=�ݕQ��X������L�/de�x�	(�6q��
b����n�4[ЦLE���֮����k�<o_q��>Dj�l����d���^f�h�S��ِ�a��c���[��g�"�˞.��zW"7�����-�O���/xv/��}R9ѩ���Q/$(9���g�vӂ+��Wj�xh�����	�#�������5t��t�b���+�Fd�w���.W�20�nPU6���o�t�ܡ�FpS�*���s+
+,t8��񚆃D�%�F��(.K���X��b�$��y��ˊ��J8Ut�)�0�I�=i�6�+Z�1��ጽ$�(�Ͳ�:k�SiP�֍-����+^]��e����meŲ$�����uxƚP"Ւ�s{���r���aQԍ���m�**e��!l5ܚ��.�Czn�V���qa�����Lo�A|�DX��,��R�r2X_a������A�8X��C��|(��:x5?QHW2���T�A�3�-��R����(3�l�k��Ψ�/1�S�ڞ���SQ�-KH���:�p-��(b���E؃����:|�݋�k��ܦ�?�l�U�H�/W+4q5t�x�8�%��#ĵ�n,�w5]*���L0g��q��w�0Vq7�>!�Z���OǈĦr�R{��X8"$4����b��~���uͅ�he*�!�D��fAv�-��hC0ٹ��`��M�*J(8���D/�V�s-֟��/����2d���`ܝy�ψ�E#-fRB���8+�Xg�'���U��3p{(�+.]�ɚ�1�C��Q�d�1�D�s��-V1�0��{��r����M׽��C�c|lr�����`Z)r��^�!_c��4�m+~��"��������Ş���<B�xqF��L��靄m9t���]$����ٸ����7���-�y\i�1	�1���� ΂�8$h�n�ISD{c�C#y
�@�=�Y�r!. 9��;2�4n��+�4YKbdl���,�T�s?��lć�����@��X�ܠ7֗�`���}�1��Rl�����y�>��ܩ�4P�%M+����8�OenR��|�8ce�E��3m!�
�5�d'�,����$����?`.�U�
�^�Vh�AY]��<��@��"��F�2���W�4���l�H-c���߰���6��T��Ƒ!��H|�UR�	3��x"�A�_R���;�2@-'�TM���a8T�>),9i��HuǴ��=�� ?�X�����r����Dp~	���pK&��f�-L���R_%ث��+ݰ�O+�$�8|mYzmS)#S<� �1&i� ������-X
�q7����L^����(��<�c
�ք�'䨜�N��EsUh�*��f�GU����)]L��X�m�>Yb��:�^�p���7�^�6@�P}�W�EG�3)l��0�*���
�"�H��?c��p�E�ۃ�B'Bk�p��O�X�`��LOB2+�?w��V��2z��Uj� ����@J���ú}����>*�_�3M���A]���c���p����y�U�?�"�4d.�Y������C�OO<�C��Ƈ25�CG_���;s�%�0��NsKvr&��2��׃f�`�B�����l@dHP�]a0�� yIz���P��+���؀�ߨ/֛�4,<q�g�|S�
����/Pk�<[�����ހ0�� ���|S�HO@�l�*Y��rr��+L#�m�	�b�X���۟�Vë�m��i58;c�2��&PoZ2�fat�+�wc�A���>���IM��h��;P��|�!d����d���
(7*��޽˵ˉň��� )Kڊ��C�	�W���?�^���)6$��5@�׎��`��C�S��D=W�ؑy������ʖ��	�->�1���RM���K�]=W�*+����O����q'e���4�xK�k	'|`8&���'�rb[�738ռ����6�qºUtvڏ���ɟ*�VF����'J�Xg22haU��U0�\��dU��M���pڽ�Ӑjz�}݇~:L�RUec�K_�^�Nx�b]��당��O���[���[<�ԖS�h���i���h(�1J���,851z���/�k]968�P�+�Ә���"��@v=`��k&D��a
5�����f�(�֚u����A��V�v�4����(��������6֦�"���ZL:j{m����=,��Lp���=c�i���QN"iM�J���O�ރq��;�ι�g-�Z���؁��Os��m�<j�2��y�V����8o~,Y�<|�(p�W�d��!��#{t��Ȯ0C{�RcNӭ]��F���z(^8x�[����%�n�?��s���j�l��4�tw"~���N���	��^� ��R<����~ܙ�;��6t�0*�S�Iv��&,��a����9�B1ʽKdĈ�f?|�uSܛ�ZnL`�7V�(8Y�0-��AQՃ�DJ����%�]F ���2�\{a�C>���He}��c�g1߿�ǚ�ln��u7�_��̑�9�b�0eW�_kMnVƑ�#�g�}�K�a_=��E8#�MO�0�7��YE��_��H�$��6#�7wF�WZ��Ꮪa��ř�ܗ�O%�:�����h��������LGϙ���xyw���yIa�gzC��K���Q��C����|��ٹuP7/e$�������{{�z�)����_���D��m*�?���$�w�������o��w{R|���C�����MCb�0�=��%^fO[���@��)
�0A)��@��o���������Ə��V�u�q��Ӑ[�2��P��Hf�m?J��+u�U�� ���l��.���M�@�i����\77�dx�=%��`�L��������4��q�׭_E�M;�����Ә���>R��u[`��tiP <\����z��_^���Ex��Hz�QЕ�'��E�ҳ��2�Y^��� � �[�F9��YN~�"9a]�"�;k���pUG�I��`�.j{�Cs�8��UsB/�n&yY�5|{�p��p�������?O q��B�X����	gƑ{s�E�t�3`u�H}M��=�k�W��qP�!��u�3t?�~��L����֋�mJ�mDFM� (;,�b����>��3
i��%D��x�O
h���
�|$oB4Ci��`�lE���6׻�����LIf�n��湭�R���e��/��R��6�9cϭ-�Q{�
��M��+/e��rL��I���E~�U�5� ��"E��2�p`zb9m�2��K����^I�� 6+�5�^�]�������-�TTT�`��6��k�:��^�KA��b2����=�V��m|Y���q��ZzG_@��D	d�@l��&�I���*8Iues���s��Ad�5��o��S[�-�obI[�-3�d�g�H�k��?`W�z��������:]�cF_��t��A������e�,*�&"���a�$�	z�59eh>e$��F����(����lpK �K���_��Y�;���9����k��vt�Lh����"��cJ� �r�#�T/PU]�	�&~��""8�"�1!B!���h�S2�0�;<!9�a�hO�0�1��O�3u�(a��k�y	5���ׁQ�e�J�\һ)��%�=7����<PEȶc����`{�]*1���t�*�(���K^���H��B�&�w0d���J�w�9$d?�Adt�l�7t�Ae3w�X'W���������&�Kcl8=̧FAQ`����HvQK*{�Y�:}�p�f�D���'�A�`s�2e��>)7��0���,*Jٕ��)��l��fD��yf}O���an ⊟Gc?��%�?v6j�'V�"�ۃP�QA�7]���_�E��{.�E�.F߬P��q���Lc�c�`	ժ裊�H�'��ΰ�ϴ5�����2��o�ڞ3�W��n
��#��T�`�dR��)��#S�Q�ӷ[����<I�����?�d���q�looK���$V������Bg����'$�yz��D$a�w�i�Ap�Ļ�ݥ'��>��I�&b"p)2)�vY߁Xy�y�����hs��2�~��j�J�	d6�L��'(r������yV&�����WgϦP����O�D�OS�C�zD'�K��P��=�j�湯��mX���BO(8�� ��� . �}����t�Kj���(������k޷:�م �#��3��2�����6�;Fy�L��S��l��Y��5�
�t���ȩ�Xa( ����Y���4o���9� ����N���i��)�����T���#�vA�^��<�
�Xۿ�[�y�����U���h���Z0�i.�d��d\o\s�y��8��`�q&��J����!I��?K���.$�!�.�彉�.�}Ms{EڡLu����
�I�W���[�8~?2��ʜ:�jȳ�)��${+��{&G�p�#2o^@7\+g�E~v�c�c����TV:c�k�3H��S��YC^#�\f{��}���ً,`�mB_�F�_U��f��������usM K�,-UǁH_�>H?^�y�` Љs]p!U��(.q.е~/*D��PEd�_0r�]��pA�����║k���?sJjf6rS���g�M��"s~c+v��S�Hɴ}e�r�m���aj�m2�C��+�Q��	�ϫD
_�
�����Ze$ngq=0[�4�z��<E3K��sY��t;�.�Җ�h�P+|9�k���
f́�C���kj��������g�V4���8�l�|���^��"����⭜d9���7���X{!�n�>;�̰4HY�Z.���8��*�$1[T�Yܴ���tF!���w�D%����m@�AM���A������	5���?/Sm.*�!I��ֺ���F��!O�s�a�"����3��a�B�z}h)={Dɡnz�ރ�;
3�&'2��/���"��L�ށW&ß��1@�aҶNf/���Nى7�B-`���ƬRp_t�3Y�?�+��b<��g�q$8#�����l)��:J��=���C	7�xr�-J��L���
�
W�ix	�~��8ɴVZ�cELb����cSEę���{��/���bKN]H0��'�d�7p$@�b�%X����?���r�<���aU������ݔ�˹�����Fd���i�������R�?ƴ�ڹ$�H�em�������{W��d���3�z���[hxR�o�TU�!��w�3K��4>3+���uW;7jC���G�_���M���������Z(��m?��{�}~��U�s��ڐ��� 	+2Y�xؑ)����N�v��K�΂Eŋ���/{��i�GH>�¥0jrh��@�R�xJk��{�23o`��)H'������B�\Jp�P�/�L��U���z�~�#/̡�i|w�B0�hxq�����\�S�@���O����ER��!!Q�ƴ�6�?�� N�7�EY�.�m�p��a$�6 jڑ�u�<��� W�f.W������E���Mt������@$�60M�W�A��OΡ��V�6��q6O�%����|F���n��X�`I��f+�`@���������/	+	�	&���}�D����F�x.�W�,&��j�pga�$Ht�2������>G��:�w��7�����S��'���N�[�۹����#�zqT�M��s�_Ĝ�*_~1Ci2��:�k-�-��.�^�}��Zq�˟�6,P�}��^G�,��~�լ�F���� +,;-9�ɴ
��$.tH�r��3{����hj��b#V���hY�&��P �-Y��
��E@��9��}���\z��ix��ˮ�j:%���;6�K��ә�"�-��b#G��$�w��=P$C�\r2)�2�3�7(����p=?��[�u.�T�j�2�%Z�<ְ�.\~w#3�e���l�n��8t��V���A��z�<����:JH���M��2���H�7M>;��#�;����[u�Rn�4��!ӓL;?;�T
� Ǚ�JTN_6�{2P��!�4�q'Bѽ�j�U�qŒ�ǚ�5�J(s>�̹����t� �bg�XF�b�j����>�pU�ہywv��?]�.����!��W`�� }K�w�U'f�i�N.�_�HYÈ%o:�L�E3Y�}A2�M6�y��Y�t��W�A ��Y,��+'�}3���xՈ�-� '�@f�2~�6k���rJ�r�F�G�e����`!cmQ��1V�w�	�Q}�zM7�X@���������X�s����m$,6�}\WHN��ƥ_��j�_�:*x/"O_W(�86\�S��|�jܛŶi��C]ݸ�[̓{���6��8'�_�]Y B�t|�4��K�� +./�-������!V�W&m1o��><@Ha�s�Pt�4�8t[���A�*5X�\"r�A�*24E��A]��~�)D��p�'��[��O)�?KhfCc6L�9.���g�Ш4��"*�GG��B�Ӄp�ɕ>�f��oN���������^�3\|��	�i��Nࠩ1{Y0a���Dz����!Ī��.�'�3r릫�f��=�)B.B�<^�Vӛ���\u��j��O<y+�ݸk�{\k�~w�ܿY&aF0J^�q]��x�xEc,x��!��)�N*䔘Q.: ���O�B��٦P��fMPT���N_ү��5g����IxЪX�-#IٗXG^K�R����2��)�gO�.�beO�`v�=Eգ�Z9���Ъ�cˊK��"�w5�?�H����҆w�{��oV���;�r��IK-"��p:?�A�!���,��p.��D�~��=e]�.�R�J�)~4�Կs{�\ڱ
��P���0KcN�ҡ�u��T���0�����r�5��;C��%�EY�� �ңf���|��=i�zCR|#2$}�q�~/&9t���?�a$~[��v�Q�����o�^��X,f����6�a�4�L��Yg��aM{�Ф��?�`P-�}O2��*��S|��84��wV�Q�S�u�W39d_JXs���vOR#���5!E���ԡ~޳mzn6�AYM{� T��Q����f�Ax�F8o⸛�U_�ͶF�b����\_�m��6�md! : nd\Y��Θǩ}��fO�2�QP��z�Ӄ�]���]+�41���Z�^\_ܱ��?H�0@C\$�cr�E��h"�+�gyM���|�{gdp��>
�U�jʠ�T��U��A��/�uU&@�Ss�����*ܔ�߿-:�*��a|L�v�C�׽�j�@�q����y�������EK�~!b���T^�2gKc_��A����� �v���I��<��82�ga-q�9V��Eoŗ�eЧ�bm!:[5��wI�s@Qm$BbV7�v5U���E���p��ɣ�V�
������<��8����/S�����"�,���q��+#���!���K�Y�s �d�� AB���Ү�4B�EhLQ0��n�Q�X~��\#��Ҷ�}7�X�ªGIՃ�,���o�����C�=�m畅	]_�h�Fj�� CNɸcϬ�\��G$ͺ]F�;��ɤ����~`7�%�m�9���ܳ�ul�J!�.� ������]V"0��ԊP�)Ug���TZ���v2�i��KDAF#^�d1�u����σ.&�2f��ߤ����HBg�c"}9�DZ��;�A6����X[0r�o��z�C�b���9�K���/����U�ɰ���m^��'T�w35n8ݑGYŷ����!�+_BOg�Gv	���V-V�agm}���^�����^�\�Nג.��e!���U���/j~0�����r\#���_������
��6Y?�V����hH�x��Ϻ0���n���+�`��z��,������`���Y�ד���4(-Y�Xö=���`�>H5�<�:�P���Y�r�����;���3�$	:՘{OE�O��,�c֣[�����ź��̢�G\�D�}����w����ۍ��n�����s8������?�#�ř�)���dT�͍���or�=*�Q"������fg�"es��F�f9�HYZH�1�v�J���](��@�f!m�s*_��V�J:�N�U��3��sb���)騎�:��	�v����?ê�S1�B����k��|4�˹{����2�&����pX9�x-
��½^h,!������7u�%}i�D�S�����$W%}������J%���� {�(��� ����r�EcD����nP��1�� ����r���R���7K;��k��6�머�Z�^�;����k�+�x�0 �c5W��i4�=p��(mo�z�]M|`�����X���Q�!�$�!(I���0��K��}J9|{o�NL�d#7���z��rZ��[�/���!ɬ����Pg-��� ��#:��3���&���l��^��{7� �����WΑs���;�������}֪d��{`EZ���7^ۥ�-N:�a{a����?�+H3z�����)�\U�
�!a��;~�:c+�J�CvBRGa��E�-	B���MT���s��\�����yҮ�	��ɛt�/�?��mG��XÁ��c�Ƚ�5 ?]Wk�P����.�%��.�kn�����'���`O���f(V=�c�vn��YKs�_2y�D�U���,
�eG�����Sf�w5�I�^-غ�� 
ij��I`��ڬ_0�n��P�[w��o����O�:�$gV��j1����=��/�Cd>���C]�;��v�������n���)":�<(�M�PIr�X1֜7^��	ya.��\]f<�yD�UL�h}�8��\S7{�ނu^�
�*V%a�Z�D�G|W��qu��P[�4i���3V'y�	W  ����ǰ�e�T_|ؚR�c71���٥G��Dq�/;R8βe+���i�=I�Jn̤5���'�Ә�8�Ze
֊zd��B���*ͷ��I�v����ѝ�����(�Ь�؀�q�����Rj�0+;�W۩��10{^��N�^�:�$��EBq�b�_w�ew�)�M���q�����o>����h��$�l'ae[���N�,H�m	vK*x�ϭ	o�/��Pg7l�k��S!
�5����=�3ˑ�/�*d2������#R?o�M��=uVH��a{zA�T�|�ƈ��=���-�)A%2r�E��f�]�R���]����z��t�޾��6��B!0aB��&�+п+;Wyw�`6L4S-����LV��秞���-���bصk��*��j;�w;���G�U8Y���-a�iȇ#��U�i�a��%�-�+��u	�5 -�n��gQ���~q.�f�	.ƃ�g��s�T����6���yIǱ�4%�i��Ey\�T=ɹ��04帪~�
6��`�F������~P�y�M+8�뙕Oa���5�=����I�'���s�a��س�T�Nǰ�4QH��y���^��9Y $�)���a�0������@#K��)1�3g2�B���j�,ϔ���Ʒ�iv^��s�;;H�nNY)3��x{G�Y�����{��	Ɯ�%W�_�+=��x���(���"��������])����.f�� �V@�
�<d;�*6�Q�\Q�W��\ّ~ގf	8�����
�@�a�DPO����,�3r$(���D�G���|fRP׎԰��_�S��6�e
tbe�����?�
���U�Ø��6`�X�c��2�	�����j���Z~c����ʮ��|�Ք�AD���Gt��H��B	�
*ڕ��+��Ba��Y�X��D�r ��h����Qn^�n_�gP9Q����@��xc�R���9q���޼$E[�1�<�)YPwp��N$G�:媊ӛx��I�/�$�eCvDZ��)�Uy�b/���6�*�j��ݵN<��pF3|Gƚ�**>ܞ�WW(�+�5f�p�@��L`x`�x�qǓ �.W:��!���]�����,�+�{w�^++^��CE���}Z�-s&lY���S�Ն���8i���[�8a�M�J��WAٗ�s��CLr� i�=����V�3�"�(܃.���b�~����7Dt�; ���� �G�!�;�m�1��!�!��-Nb��d�ѽ�90�c���&�{>	by�R��ΨC,�JkE�1q(�é�+C��]�V���*��"�=T���g��̐`x��m��bn0���>� �d ��iT�?�ۢw���X�]��L$�$>μ�4Ў:�� mm��6���C%�2����T�3��=%Ly���8P�M9�n���M����^�cЋ�r<�u�+����ؘ���I�AK0�w�ES���k�'�*���CtX���Zr�9����	M�H]W�̗�!h�E����vJ�h�-�0�+��
�8��	b�N����A_R��+�S�7�	"T��lO){-{{�������+�-6͵�G@U"F���NL��e�2��-��Pqq��**e�AkK�q��S�DJ&rY�Y��z��Xh����Y��Y�7|���@������Lsþ^(,@�n�96��!p���s��C���f��=�B�w z��,R[X�'�=U����l����cv0�:�з���(rA?�S��r(�#�%�[7Z��o?ήll�������<�ݘ�	2��z�z��@�y�B��Gd]��ƲbJ��'zA�w����D��i��NS����5�&Ƿ��#{���Xll����H�U�x�£��烔P��5�+=���	/�W74���1l�����[xi�s��)�,��,���# ��� P�i|�N�g�U���l���Fc��(���G�`�׼6$ȳ5�#4y-+�hG��KY)�F���otU�l��܅Զ�|�2�5�G6XpCj޷�̰�tc��Z���2�=�P	����Ѫ���,�B3j1$��ksOG�?��|�t�QYk��jd�_���ef1U��1w��9�XH���~L�{�z�4��B���
6���4QSΗ��������vQ��X�4\��I�$5�E(;E\y�7?�vK�d]�7kv��ˬ���˂p�
Qx�S|f��?��@���*_����?������n���ndx��'��z�"��x�A) mj��VU��Ʋ���@5%�ߎ��q�B�5�^cJ>Z������A�N��!�S����QR1�iO�f3!7��6�!����"P�le���
OT�4��.�����PxlU�ty�Q�4
�[~��./�5=Io�+3�-����2[�JZVt����ݳj�v;�̦��d�]RuE=���e�{�	���~�)�+.�@q;4kX�<�j��ך��,J���G~�G,�\�-D0��NBPk�̿�7u��u�/����vx�����c	T�d�0� eD��MA�W�9G�@RU� ��!P�,E��`�a��Y��m:�fJSga��cT�}	E�o��5�S-��7�,�w�9xY��ka6�o��B�]���8Z�God�__�^���K�Q�X+�m5%j�#5N~.r�t�3/�HuF
���UΧqu�ǀEK@���$Ϩ�y[��=O�f��`W�TS_�7˴r��kw�|��PI�[:ⱌZ�=�5C
06@P;V�a��zVXsH�����Z�B��c�z#ǟedc��?KO G���jػ�1����t+�����>�'K("�3� \�����2&^��F�'�V� i�X���s[�9�M�`m�������,`�?amPo�����J}�nT�E���pZ7�T��R�0xy�g|[(����{��_׽>3�ѿez���CT��U:�U�tƺ����:�s�,pdZ7>ja�!+gs����|����e-�g�V)8۪L��������̘�O=lO��X���6r��I�5(ݼ��z7v�
%���3�^[�ZL�g��Dȉ�ŧ�u��P�CF�����IM	�n�	lFϫ�2.��ce���۾/2\˨�h|��L�lM��t	+g���D��y��Y��)[+<3����i�̺��N_p���7%w������}<;�l���^}VF�'F��	���G�	h6'�pX5oW��2Cq���]�C��+��zD��:fI�?�M5J�X��B������� @ki ��gv<W�>��'�0����2F,
Қԑ�q���X��3�R�):�Ӄ�Εci.!e_5������_�"ħ?�'8
���.�gDXhw@{UU�<A{L��T����D�}#6i9���9-��ݖ����]Fc�c/i�������iX�¡�p��)�:��`�O6��_)u�:��H:r��Ƀ"��	���3B�MI{:��π�#<
ή@��>F 8�Z�QO=�0�:�8Ay/wV�~K=̀�������N�f*�b��K��_�B�6?��7:�<g}�V�Ўyu�W��&,�7ްТ���P>S�B������]�`py�$ˌ9daI���M��H�A�,���Yf:�ʹ�XO�F)h�y�{ �m-�ˢ�$�>lV_�����C����2R�{�p>g��{rĝ_g�p�A�bq�.m���T�ʲ����F�b��m1����)i��n�>S��֭,^o���<����CJ��F����Z?6ן��x.�qӉ��0W��B��n�H$7AJ�����펖���#ɪ��D_���M�r�3��b.����̷�j:�S~�5������l�6&+�924�#6I ܧWtj��@�����Bɚp-�Fu?��0��hu���8�O"��T|�jΎ�)D��Z9�05�(v����!�C��ax�\�i�oE�>oX�����4��GI���&�BR��v]Z��N������KO�Ȭj7~{�x1,X3�J}�ۺ[1��B���B���.?��k���y�/��#�{��9=הg�aB1vQtr�L71j]�(��+�(�|(-]����	�w1ۼ��(i!�񾆇�����0����%��lG�
�{���	y��;ȿ�55_]�����?m��T�4"�����d���O��H�:��1(EL�� �3k�*��OL�Ry~U�ŭbDT�j� :Vf��)���sgN#u�I���Fm�A
�<����c�I'��P߻�<e�ɬ՛q>��-�c�8>ڟw��w%����S�;��di��Q��>��
j����f��ڛ���m�}MD���^Ei�r��d�P+��I�
�|g�t�pR
���WjeI��W"��3M�qj����V}�a�..�+I���{���G�$13/`gOw&����ϓC.:�A`V�oqk}Q�0��6a��� ��j�]X�X��&�O���/�J 2%4gZ��� jU���7�����o�S#�m�W��=D���g	��ф5~}84�*�+�?7��{�������%`1�e���vpd��1DDskL�����X4�Z��ܻ�����cYF��рd��� �w��uּ�j1D�]dn2�ʗ�w�3��|F�pNh�q�D�ί��P� s��Z�]�E���#qp�
�Uf�.�
�)��Ҵt��߰MwA@r��h"u/,"���}�&�����U��n���$��%R�p�hKgW�F�ȿ�G�8$9'455��H\�V%�Ӎߖ7^�_�%-�$t+y�!Q)J㔬�(��w#������+,��{k�~�믲��9�9��Y�h{�m���5���͇Iy� �L�)1�ᇨjq9���SA)�������G��v�Do�^�#̓��	JmŠ*����t��`	Ru��η����K�!�h��$��#1�5%DM�ڠ��}�%pc����E�T�h��G��[/����qG�Dez��[-�yN���%�ݾ�d���O�0�݅7.�XcS��n�ڜ H]G��ru��e�ե�jiz��5��{���c�VUީ�ծ�~	;io¶o3��d�c�ʃ dp��b���6&*ߩk#�yfJ�ظ����!�W�AcO�5
���M�$�P�AV�{777��c�']���T\v��}@�C� bw�a�����cH5q�����b�~>c�#�����ڟ�^E��&%wh-鲉xw\?�\k��PmNE����RG9���H�v�� GC_"��EN���?T=�^@����w&Uv��wz ؍��)����=x(P��T:F��0%��.6-�K&'�`*R��_�q�$4�����LM��%o�������L��r/�]ޡڐs�➛P���/�=��`'k�C��}��SK�*�M�d��*��^�����)��"��8���Y���Ѳ�&�z�\S�k���  4��	�gh�XG���W�ɴ�6b�BoPy���8��%����v��յ�?��[��B�w�P���Y��>)��U6��z	�����nvYg��������O��'��OV�B8�)�Б��π��d`XI��*�p���L
�%&�i�G��)��@��dq�H���l3�����ƹVd�
P� T]�`+�ڠ哊C�v:��G�S���ի긽t+�5It�U��O%H4Z c�T�֜NY|)xi��u;��BTBD���	�ߚBO�9����=��`�8���\�����tRGX6qN��h��mݓ���"�̃{���S>HZ�À��rb�}�K��o��5:�VUF�%��o;���E����U�K��k��`�~w1_�q� ��O:䌮w� ���s�$��Q�Dkv3��:�ϊ��{��T��?�R4��'����A��/��[a{6���d3q�@���r�a�I������U��C��b�6We%��	���!A�| {4�k�Re'>8j�\�X������<��HW���&���SZ̻/����]���H�x�[�Q��8?�۴\nx����}�e�� &L���Ϋ��b7j�|1�ϥ���u�f��C{��P$~�&�脠�~�/��������R��5zx��)�a�_�!�y���J��h��'���2��i���#�G�
`AfX���*�v�z ��ϗ��￹�A���`�(�SD����K������5��,M{\�'oQ��_n�Y�ͣ�c�%i}m!��41[����/BY�������:Ғ`gc�c��7M�����,&�B�/��~[�#���
z�Y#�l���.�FҤ�1٘!uc��(�g�]��GM6Z���w'&����R˞�L�ig�9;;>g���Q�>H�o��j<f��GZ/}[����I����\�˻k�Q��է p~��ǾOh]��J �Fp[��z�EI��f����m^��A��Xg�oJ��^�?k�$cL�[���p��j l�&�7�A�����p����UY�%n�f�Q(h�����N�*���ė#��##�_%���8� !�*tX~�oV0rP|i�iA~�U���[��D2��y���+v�z��g�`��{p���4��^/�%t`}�j@l3=����()�;�*'K�~�c�#G�q6��;��0 �������yp�U���ǧ��*��^��x��I�Z[m�l��qi��j,wCo|��idR��U�?�?��c��>�JUy2�����#���$s7/���4��1�!�A�E����3:��V�4����9�v���3S1�l#�ae�H��u�J�	��U"��gw����7ʊ��M�]ϛU/ݮ{��-L%�	���<Xc��HB'� ɁF��\��s��?M���P���oB�L�:���_|�Q@�-�yu�Ү	���(�F.ϬA��U	�ç!�6��q��t��7 �Ol�QQ�'�{j��/~!\H�~�aJ�� 2����NÏ?~L�7�X;��Pڈ��5j��Z��%T��A�
�F�4���EK�s�_�{VJ�P������_-���Q�:�`²-M�0L�Ʌ�ź���^����M�7P���E����K�'�|����@������C>oZ+cQ��n4��Cn>�,]�rB�ܚ.��:����Y�$b��Q�.6�촿;��	��p�"��
��q� ʰ�x�J�/M,�/��q�Z����9-������@�shۂ�!u[�|m��P�$oX�1�����,-�����_`��KN����;B�S�:'A�[K�sP q�l��Efq1P�Ю�-����jH�vg �����`�A�z�F�!����6R�������n �r��+�i�>*U���m�tU=͹/%�a/�Y�À9H��m"bb�Z(?�F�/��=��@�k�+�4��2sxp��O�|�������
4�q�� �]�a��fK�b�8���G�g:�(:�,���t_���b�ɦ �I�G��j&t�aG�@�pH<\�\v��Ş5��A˿�k:*�tV��K`�a"=�2�u��4���O?����y)�Z7J�E˂*��d".�"�-�����ID���kRh+J��t��d�xWm	*���/1��$�q�Vv��O%J l���ȭ���ݶ똌�0�'���!��{��E!�����,�B��p�wR��s�P���N��@��ة?
�R:�t22~�>0�s�X
�$�`��й/�D�Ru���5k��j����C_`u��C�I���G�m"sRe��5 ��x~fO4�s�Ra��ө�u�'bl��a�:ૃ���9S�J?�5
�-ͣ�2h���*  �����6���b������j��(�x��Z`wW��/}�=�s������X��7:��?!�3��|�a1A�h��ѨY�q����(�l�$m��<�З��R���d�訂W�8�8�/��Z���ٸ�?��x.Dr{F�â;�`kO�Na�\��~��,�l����;.��?�#VCB\V&��Hv��#��3r��_���,8�ru��2�p<W 7d�0���� �0�瀠�Ϡ'?�s0��]+f�t�����6nN�hu7b�z��~V�8Lڦ5~a�F�#�W��ۆA���;mH�N�D�_&�`�����h��K��.��C��72gc7)A��k��P�5��_Lt51��%�V��ѯȏ�H�<�̾Ͷs���:���^޾�'�5�s �OԹv�8�GJ��Ԉs8��U~���U���`6v��(@������/��3�Ƙ=�Q���D�ZI9��D܂��У/����"h�8�~d�a-�oĸ����h=�5#
S�)T,�x8�G����Km;�\�Z�٧�ur[�ʙ�k�7vk��|7��\��Q.E/4B��eaʙS��hZ����Uj�^_^G&-L��Z�X��+��H�v����8rT��7ב�E>��C�ђ4����o(^�N�@�����ă�=�-�����?pt�����P�"R����5I|(�l����M(� �=���Yt�%��t���U#���*��߸��a��Ճ�9�`�$	����PM����`e0˗K>��9�]c/ͅ�(�Wr�2nՎ�'���"{�;۝!��Bjd��we��8��w�ac�V��I�V���:�Y@pQ?Je��iO�>};Iu�_�o�ƕ~�)-��U���>'����] ݜM!|��F�����=2�[c��__�-�*D���c�mi�8r�J�(� 4����{�m�܏�,���� )�a�He�ꀻ)$e��$��u6<A{����'�ꀬ��'_`���n"�	�j�]ivZrHt@7@b߇���6�`e��,�a�Y�k�e���5]�{�.b�^꣐r��f�H��.�������s]~ۼ��HG)�j�����C=����#�R�/�� �"S�:vT/;�%����U)����:V=F�&���_� ����¼R�}��_�-�,���n�=��wy,��F<���ޖ�ᔢ��GA�qHD�8�q!%=b�OZ2�+�ڶE�#��O�����K^���n��4a^��	�6� �!q&����ذv��I�D�T�E(� �.�=�A�N%R�`C*��;T_V]�v�7������X_�5����ړ�����m��I�ҭ��e�~��.}��O:�-g�����QB�0��ݹ"��n�z���XZ��h|���[|����k�����l��$(���s��X��U�Y߄F���׮����R���}0^��@f�����^պ'/���m0�I���X�dp�<=,��t;�%<;�,|���u��:<>L���KT须��$#�t���γ���=r�Ӊ��[b	8i�[��"MU�K��܏�k�7���Vk۔#��PC�� �-3>�NW�8f�.�ή�r�	�ه/l#Cbݶ'�ʾ���9�:�D�t=C�0&`u �hk+}^� *�WÜ���&���2�ڧj��TO_H�t
JR9�Ӧ�1%����.��E��\cy�X�m��}�OEB���Y��qD�PH�J�_���Uڎ�(���H��ýn7�Ћ>M��@Lo+�-zL��lm���x�8�1��r֨�C�\c��k�5�)�@��s����ƌkL�#�yv�rs;�=2��(�G����*#2z)$�s���� Zxp0��� %@���8�oD�A�S2� ��gmi?�o��]U~���b"�	N1�ul1�;���|�,oϰg<�A��9],�h��y�?�#��p/	 *gu��a��EH�r+��6K�:?��2����
�H���b���yOE���+i�V(�A����C�r:I�^-bØI]Z�b/~�q�X�X���PT����������VG�9L��q���Q�,�� �D�@t�>��z��P�Z��x��w�e�N� X��7b���lТ��M��=y��4������ /���okC������]}�	����+IX?��S�&�}ň�ݜ��П;�곋
��YF��Β>[���3��C��Уg���)�9$�k���N֫r�)	oUR{�8XOVy�u��A>��P����kg�Ϧ�qqof�E6j9x����$�18�mc�����D�T����z5����t�M�<���l��vrˊ0�S�=����.k�HL|�A\p��7�}�lۂA���o�W$��/6�-�J���+$<49q>�z��K8�OQ�?����{� �����g�O���x�g/�͸�,�τ��in��_vU%Ջ8�ʪ����N���*ǒ�'���&�JF8��Pr�K۽g�mG��G+a���r[7{��l��c��X�U)�`�*k�����@*��>@K.����+Կ��+ɶ5
�\\6�'�Z��A����)E�F,s��R�b}���MW]���t�I����b�wE �����,J�g���Dm��-����<�N�����Q`����?���^������3��_����m�T�xЬQ�G7�T��P���z��=�
�~ȁۓ�~ٹcBpu���Y�{G��0kJk�(0�����a����Ћ��^�)��2	�oZJj�u[���b�?~��Z2�<��O�5��;f���&r6���c#�3nΚ�|��2�f�ۘ�
�]j� �~c�׈uΡW�E%����N-km��)��ڴ)��aq��/��y���=h�f��y*5e�.�_E�pR���Y6\��Zb����������3�?/S�lYa4xՉ�^�	�5�1�/�V�p�4->fL°�Gڃ$[/�a�������� 
�)�qT��r��&�*C����{ �,jO' �zH�٩��m�4�^�c��X��N𓱁~�2}�cM�����TW�m�6AF��x"��Bb��<�.�Q�cۚ"*%���ix�$�:o�|�LϠ����2J��̷�>�g���2ˮ��˒@��>���'�/�.-�]���@�&���erc�-�P�Z��pj�&�:�~5ʹ�">�f��B��&���~ԯ~M8�>|�~O�����Yq�ǎ��刬��u���\�U%�tp��.�畊iF�r��7H1�.�c��Y3/_��s%ٿ�,�l�n2C�g{��}4�k1�%������H�5֚;Q����x���y�X�*'�B��g�j,1v��&~Ms�I�8 ��j�����w�U�(}t�$��G�N���b�8	�����3�)=%�r1-�*����q�[�*�{y��"
���W��o����W�'4)6`��:�f�v�Y\U�r`�O s���hK0���e-t��q���?�6
B���\�3�^�0���	���J�@6���3gd�*���i���z1=|����<�r@JD�t�CA����t���6�!�1��۟�ڭ�^���ZS�Nޑ-l��B~���	Ʉv�aO�pm��C�jiHI�蘣�-r�i����uq@��v�����2!Qp����n�]�RS�BW$��'!�갂�W��%��^؟��Z���s�ݣi�f�C�'W�aG��������[o=�!}���Ti�Ȱ�>hF�N�;&c,�X��*�V)�Cֺ�j���"����� ��kݓ�k�����`��Md׌3�o��rF�B��G$IA�w*sq���qv.?kP�Y��*�����(����硾��ծ�JϢ@�5����?N��s�Ir��B�Kk��N:��b���b�0���Qv����z-��i�&F��ª|D]	��i+����y�h��m��i��En �XV�e� ?���� ��j��2O5�r�/p\J+ʆ�����/=���R�8���lj�����fB�V?�L�Ժ"��`B��������ȗ�'%Mj�\��DQ=�U�_3�uS�1b��q(����;��3:�cd���bHx�O�	ay��M>�#q�x�&Q�G��7��*ū�C�k����^q���ؠI�K�VJ��߭����2�"����n���@fr_��z7(B�k��F�QzA,�����g�6�qE{�̍E}ymb�cN8)J��Ѓ��ag�>�G�O�p�0\
�J6�eI&i(�SV^O�í�]��!�R�j��tB))5���� ���g���Y��3W�B����u��0&|"��_��`9�H�2�\	�u������eXE�y^����3�턹t����@.��on����R�>m�aq;�C���4��Id������MV���Ƈ"�4��Z�u^�E1��0N�h�َ������izٴ���YָM�������]1-�Q0k���g�^��f��wy֐[�8o{������e��'�p)��+B������O���x�73���p�7D�����+��)�#S��$pl��ѡБƦ� ���y�ۤ��>LҢ�3�3�.jDi���b�g�./��ʂ;����pΰ8�N��8z� `6�8�M�Ri�Һ���m,#�҃;�P<�G�������
�>�z/����ȊWj�����6�S���/�NY��̵�G�d㸏�Er��ݯq�9"��&�j����E���ޙOHJ�3*}1z�S�1}�`mC�O����>��1�b�Ә��1�:sޟ�4s�[�*�R?!�y��(�W>�A�7�z��d^��\�ZSL��a0����}H2˻j��4_�'�]R�������u�; � 6����F�V���.��N֢
�Xʰ`ҟ��Qs�5�P��WZ�4����������O�F�M�BM!Y�;Ӭ�I$6������S��g�U�W� \w�QE�g��^QKR�tt*.���#{��������������Ig�%Y(ɩĿ�pê�aj\�]s�%�4�x���&'�d'X 1p@�L`* $��٤%6�H�C�x"�H���0b���v�
ҹ�S֫��\�*�YY|u�B��h]��}�=�.K�*.׬[[	��p��o؇�y�fT)$�ڜ�P|���[Kw�Zs'�Ψ��m4�SL"�?�yQd?R��I
N$~s�@�ҭ�� �ϭ�2�A��W��A��N�נL#�T ���O��Χ�	G�'=�� �mw�5�϶���t�S*�����\�L����z6)�{�C'�����ly�[�1�#U�숐���Y��V8�:�S�e����~�k�����R� A��.�X��Z�����7�c�t2R�֘E��1��s�J ��U�z۔�<�
�ï1.7'��j����	�Aϕ/�5�cpn�-(��uf�5��T�����r<�:�f�a�^��?C�Z��Z!ϗi�?^�2\��롼�!�\{��M�1߭��1���9�HE�!l�:{���+/��<%N�+qޙ�N�\CV(��l#%��b�S
�N�")���ky�*z:.��<���-W�y��&�����1��<�!��rW!�m���݋MS�诨%�c"$���4�o�Jԑ�9N�A�������T���<�!ZS$�U������d�K��#��5v= ���L�B��'�eR���筵�JЋbt-c��g-�1�|���V��,oPzސ9Y]g橕���5ϻ���1UOt�">��$%<%��Ì�(��SMe���n�G�Υ]��8;F�*���-�%��q���x 3cB@i$R��(�֗`Y% �-�{(�Գ�(٧A��ܲ��IH,Ƀ��9篢�_K`r	����ǂ?�9�:�_����Q�\!� �|��:N�heY[<J��{�,�<��g��	�ޚ��7��q<�j��b���ރz��D�i�����Jme4��24�'`�t�*e������æѼ��\&AI6uVÚ����ky��!t�٤i��SϘj������x
~��CƔ��9�x<��*o{U{Ɍ��u�T����Ԃ��>H2Z��z'���7�f���&ቁ�W�C7��I�8�3��W��>�[G��v��a�Mn^0z�J�d����s@�u J����{W��)n��>G0�-�%�����j�{��X`w#�;�t��N�bsv�D%M<}'ݲ�	�,�r�>������9�E/pɠ%蓩%G��,1"�\��	�VL|�/s��]a����Yc���kP�A&�x-�0�)r�b�Y����WZ�����ډ)_�\ʮ0�5ȿĜ�5�W9�U�8��v��eh	��E�hn:�8��Զq�+yi"��j�s��a��q��� ��~B*/�RB����|YR^[���ge���V���"�{|F_������Z�%�x���&!����e���[�b�xѐh��1�,Wrf�эJI?��	��4 �k�q|ҦIy��͓�f%R���.�)���cU��W�f�&P��Xf�M��(�L��}�
t7p�P�y�R4k�j҉[5x��O�z�ѯL�I���C�FXٓ#u�U�B�8�0r��L��C�9�����\��x`
������3'u_j'6y��?�l՝wF��o
5�j�9?�-���ΰ�ff�j�U`�hss��4��[Y�yEk��^�Ǣ�n����ˌhm�|��'�v�r'�brc��N��-�/�~�A����ݙE]��4H�%�eW	�AQ~>B�"��_ҘȲ����/�8H[�$}�,>X:[ʱw�_�{QѾ"���;�ŹYG�A)
m���\&���ǘ����ܼx�}`J����'�<�Z�D���r�A!B@����i�d]�
4�e��W,?��E�N����˶�5���٫�K�;6^������G�79�Auḥyi\���-�O��� m�g�~C��r~���ʈ�T���M2g_:jH�~��^�Yg�w+�U���F	W4|*q�9�� �)A��4��H���� $|Jr�u�WTg�>_��#Ҡ��8��6�QNۄ�vg苾f>�ሡ!y� 7�F7�tu=#u C3!6�ѥ�[]ť����Ǜ�֯�ö�T+��Ta����H�+���]S��N��&b�O��Վ�V�����8�n��O>-ťd�q�vRPmW��uڇ�n��W�&/���L�4���
_J��,���Mcp.��[��C�ʼ�ZQ�t���_�������"�"$�njSȽ*9D-2���.�k�GJ��M������9����ޚ�EӴr4i����ٲV3=(����vZg�z�&9"�m���q����f؊+�`������g�*3���Z�Y���`~�~K���}�u{��
�֘�N�X22�~_�ICʫ���U%�8扷Y`�{�1��Ʉ��U\�3���	�=��J{�,��jrd9D�7�$gchӍ�Jfײi�C�:����A|�,��`�.2d��;I��Ӥ6WWX�����Z��/ ¾¦(+L���v-Q�7�n�.���v��k?�Kk,$��ww��DNJ���j���?��-K���Լ@��'2����^�W# %y��뀌�T��^Q,����8h
]�������Bi��h�޲�����J���9M�[8!-��(눸��N�)����A�6��O�=̉J�v>8�U���Hl�����M�e�ؘ�*�D~��hT`��0nxwLiM�05&� ��d�g���ɛ}m�DPfjf���j���G5�Yv��N �$Y�>�,���*c��q��"��S��`]*�4�~���֒]^m_"�%c�M��T��y�A
N�*a=Y�5�y�]4����	�g�e�l5��&A����44���9���0+�E�\|�rP�-�;���Ѐ'!}�iZ�m�N��;p��J1h��A*�W�}�?d����A^�~�O^��$H
.�/�;0ӮN�١MX���m�Z�ن�� ���b�m��5!b&c�/�,����s�ʠ��tdSJ��c��:�|�b0��0�ΰ���z�Jd����^^���~�)�3]K�XZ���#m��@�v�Y�F����{��i�Xcؤ����t����[-Ab� 4 �
��|0�q/���-���-���S�^_{�����|]�B �je8>����c�"�H��WT�Kd���%�z���<]ڶ@@q,Dĵ���!��IpԀ�Y*@�Qt�Oo�l{��#���,�*4�2�p�XS_"��LV�hD��]8��Q���`-Y>q����W�?��[{@� ���@�6���ះIF��m�3|���1�Y�, m�M�u�8ͪ�奥f)���ʎ��w����	5F�a&P6�qm����C)���|	Á�'�,s�@�N�);t{r�Bg���<Z�%zj�,Q�u��]A�J������bQ�C ��6��2�[���%�����5E. _tT��*ìtp����iE=���10����p���ڞ�*�����3˷ ]���o ����?�X'r@e*�X�f؟�@��]�5�H.�Q�y[A&q�NYh��Z�E�W�g)���.��M�v!'mOՠ��
�~i'>/7,X��J�ϕ}�0�
�8}2��n����]pv��Q�-�x�f@3�,�1Eͩ��H���B۽y�3l��CY\��F���5w&�``>�j��m2�j�O����Q�"%ڤA���e@,L?4���pY���b7�&A%���#Kֲ�!e��>2=0(MG.o�洠��f�=��R�X4���7�_�ىH�v�B{�o��+�����3�f���>0�����)#Hi�$��~�A�^<���D���Q��@4(~5��@�=ϖ�D��4�����A�Y��f ���]rx�h�f���Ǣ,ͻ�ck3����
��C�ib�ە����sect�t�wKި�FCi5V�?��S�b���;F"e:�v2��⿺?�hFP�S�
E���b�?H|����}fl�>�����;��� ��wi�B\l�~-Do0X�Ĭ_����|t3�;~h�9hk����N�lA���s)<�.y�F��M���{r\�ByFT���&�n;��^�6t�Ղ�!?��ZVj:YZ�V-���&l��6s�:zd?
Ip.f"�����)G�H����#j�,�)�tֆ�D3W�����-���-i��Y���/g!ӭ�b{!��xZz46ּ�l����ޫI{�߂���Bl�ݣ@|��/R''���x]pW,*Y^k�:�A+�<%�'��3�QpK��a�u���*9�Cx[J~j �ZZ���"^�eU|�ä��>�	��4��y#�Gw�~�c��=�q�^�b�&C:���2���qQB�����\F��d�w$`�_���K�X���e��:���~���*�G�����y��Z�ɐ<沼���'%����D�?�`��ٻ�_�5�F-���C;��ByP��A�];�)]���p�B\�I8���R��m3���������P�H��!
��܈S�7!k�FY�� G�<pkQ�}��(6��ŜQ�-p�U0:��1�׀>�'_:oB��� o�|#2y.˭LI�����\T�_�����IiM��+�s���:�wE�Jgbq�kP��W��=۰b�"��R����$�Fb0���FYy����M�m���B=j��?%v� �c�����Gh�Y���,9SԸK��ƵxX%�4���m���7�5�D��|��_�=����R6��/y7�f���g"R�����ң�����Ӻ�ډ�>�UU���2����+M ��=����os���`��C��x"�&�|FTzb���f�1��\tQ�;�7��-�a��\9*�".Ĳ�]DZ$��Jw�;+�N,���5���a/�R�6�t}��ڠ���>@��0�s��Ì8:L{�����X�	W��C{�>_�5����:���u/	�������P"���=R=b�T��J�U����&[L&�_�H3H�H�h�T�2>�t�A��18�r�sB�o "�����`�����sߧY���E~��zF�x�Β�5����"�,#�p��uS�M
 =b�^�ծ|zc���T5tq�b�o�13,�J-YУvх�Z֑�s�s�R�\T#5��9����jX�������p�fX�D3��\����h�/�H�a�U���@A�$�6y�ADe-�������
���<Q��/X���e�o� ,�"�S����
�yL�Z�N��hk�q�������i;�!��R���U�)�Q��:���O�'�[�m�å��'��2G��&���%��!r��>�6g޾���]��IN���
��xqz4ǋ޾t��B����ɕ�u�_��<vy�&F	ͷ�q|�~��p��mi����z"G��Y�m;�5���O�_��,���X���Q2Ns�.$[@B�H+�q!���t����k��N�����$��X���(�P� 5��{��[̓��7�aG��LǓ�d ���\$���%�r��h:8�h�-ebx�mbxy.�\ �f�[ڥ^�7�8�X���*)!]������M� #z�ډ�C~J��VR�a$_�i1%�̙\Gr7�d�O��� �r�.^e�Zf��"�௑�BPV��fO4��C��d��$��m�I7��=�����rikt�/8�H���	���<����/�_L┆��\�h��6:'#0/)`���:&����_#�����#�9��}a�,8{=w����$�7���S@A��l����\u.�[�N8��J�x��q�_+���+"��i=�i9'5�QA�^ 	`"0技} @p��c'ft�I9��]WCb4iL����[��)���ǎ�W���Y��h>�����u���j�9'l/�wI#�J3�Ϥ��8�@��ӄm�?R���H�TLP?!=sa���'�ˑ91��ڙ�w3΄��:ڄ�Z��U.�m~�m�l+��`2���/��"��;]���/*��']�
��J7�Gqk�?�⳾�;�/�%F$��:�|&�t�M�4?�fTq�F}�?d��'�Q�d҈�<�g0-���w'~3��j�>20���������s�?��W��Em�O�GD�|`�W��gP��ѥ���*��ԝ�6�|ŗ�)$�0�I�΅����
���П����v�����Q��0���w�t*[?�Rv�z��}q$�0�=P*��$��;`\�y��1ފ˒�/��������0D�t;�ʒ�Ck�o���/1p��R�������u��&��酟�d(~2zE���:��s)C��/�t�1�n�u���u���:7���-Òʈ�*���6��6��Q���w���с��H�kR��T)�0ԧ[@��h7�S��T�jVm��(��z����e��2L������͵C|�X+Z<8~��¹a�H\���:v�_4�<l��T�_�x�Ū�e�t�T��PX�5�J�	�4���+U���n4Ŏ�#�2�Vq����∨��ٓkk$��e�*���b'G�����j(לQ�itD&��y�h�kn{��woҰV��!�?G�@|BE숗o�m"��C��0
���*Cʤ�Z8�p#%���KY�3*tW��������	r��ͯ��2^}�P>����ީY&��}
�W~3��vQ�e ��VK�
y��C1J�$��4������6�Q�����ZďE�A>ݓ�ቘ�/3�+&� �ۑ8��	�F��?w��X���y*�]�P.�*ur<���\O$Z?��\�X��8:�4�5]C0�Kip����閉�N��S+='I�k��l�����I��.?�6VG��w���G4Ґ���RҖ��2^�3�+nu�9�R��1��gm������.���P�󓼏���}��Gd��+��d�0ӭ���p9�ML(@���k����Ws�8S�1@V�k����������Ru[J|��4�K@�ҫ����2�X�T3�<Cwx�;{s"�{9�g�V�'FG��Wf	~'iޑG;s(b��������|���'�^f^1W6���p>����Gcm����n4#��]
'j���l�"��P���F2Q.��ˏv
L�}M���:x�0]���,�_4�ʢ���)�bA��X�n��t�2b�_�qs�����(��H�\gC6>����c^£c�F����x�)];��})o8�$���]�%>hi��v������Y��2� ���B6���>�ZRF%
�ʷ�lOg�{��� (��{%Df�b���'i1o�e~�w���y�<V��jq�tx���:�cz"W�u'Y�y �_c�Pl��ؖ�Or�G�a �����|�	�k��?*�l����x�6ܯ�g�C�fD���j/���S��͉��G�W�#ū�L]�[+�	$���Pl����e�0���.p�-;MjЉ
�Ou���(��AM��]1]6@�u����KҤ���D2�R�4�_t,�I�';��UI��?����ȩ%��7��N�������%�
����x)Bt��P�VJE����>�ͻ�^f�kO�}��{l!�%���%�~%�:��n�����`5������Ǖ:��U��-^ɤ�����`�}���T���|��:�2%����~fK{ӡ|���l�:^����~q��"�HBZ]���tH'%;���L��[%G�o����^\��g�M)�]��)�J��qH�
јL��#f}E�Ҝd��K�=P_�k)A�x�����AA�x�q7��(f���'�8�;�`���E���A%���d�H8��	: �h�Zfog�7[�զ���|M�T��쐅��1a�'��� �+��F \y�V���,ت��[8v(���{���7,�.Y,8�&-;��Fxb�,D�w�}���t�c(��H�]���q+O��� >lu�r���c�ўu�m���,ާ��.'&-@�Dm�h�Ź�_�A_�ۥ��E뛂!3�]H���oJN����6U2���_�Yg���jX�F�=�83ă��|���X<��Gs���%d�nT�}���>*�'��4���N���`��_���X��_EĕB�?a��J����&C����j!rme���M��b\������P�	��Arg��ĝ��D~'27�B1�\b"�8�67�-~oze�*��Q�P�;mL46�8�����\�@��=]!r�S��)�a��B1' �њ�K�l�ڏ-�ݎ�����t�"�ٖw�Yj.�]�fth�gkI��a+��P��`N�$C����~��Y�������R��ӷO^A}��[��c��e�W�dI'�\ʟ�C��c@�rΤ���ئ)p��L�H`�T{����qP��`:d#с=l#�_Ǆ��S0c�5��}�\a]5�x�����n��@�=�oER{$�Mט�)�#��6W
�,�䝷��ߝ߻?hD|���s�p ~��������4�4ZQ0b�K�xa}�Y�P�Mͤ���z!��x���m��X{��wA��u��sW>h�����������ObWY�s����c�s,|<������,�;��╢�~��a^����+�����
�=��.�ΣZ�W�@@���iֵL���t ��|���,�N�r�E����:Ec�=���s��t��[��wɵ#渹h�m��=��n�W�Cx;,ߠ>2iy����Q����qx(�����e��sF�.;$�?�O%Sp��zv��G��^vۍ6���}�t�o�S2����������
�z��wp>�u��!W�	(�^)Y�o&Nk4�k�q� ��-�n�v�.Xh{���έ"._�`8rÃ�����U�E�~=��@:�ӌj��[���Ő���.ӱc*s� ��Q�Q�R���,��F`�vY�׊���ÁR��ٹ�N%y7%�|p��ƣ���pf�k4� ��ي����JX��aT�%��6Ր[�r/�_�Н@�1�
u���� ���!�͙���[�
�Q2�]ǫ�xٕUD�d�21M�d�Z�����@����coDAvr�ԏ-�y���r7��ry��~Y#�(���n�E�V$)�~���ԝn��/��F.�-њ�̭�s?Dφ�l
(�<,�"��}��o�c-�wW67c�'��c(�!+o��a�O4b�x�0�����Mz������	c"�<��G\�(�+ ���;��B%(��Y�����w]�ۏ��2��Tp��,�j��yN������p����� +�&	Ob2�簍��!�ǽ3�/��Uw�t���\�h]�$���&���;�|��AJ�"�:�0�7J��<���m��CT &����0.w�E�+	iLg�;bdBm
�T |��s�B)�S(}F���d�ŀXGw��k0��2�t�D�A���Hɳ����)(����d Q$�e�eGb��K]�\i��������׎\��۠��N	^ĈOjN�稏��IQ
��S{c�	!Dd���J����1Z���4� oke��O s�p����L�c��ЅDð��s�-��:RV��c6��z���a��V���_�rz/��5k| ? ۻ�xQA�V2����<�qk��N8�f�*cQ��[x� ���*Pa㗖��,�E%z|2JX���ib�� �;=�"��Y���T�,B�5l��'�V
�*���,k.q[���W���7>����?xq�c�A�U�3R8�5|}\��OL�*�9��~^����+4�2�[���e�;�lU*C�,*�Bwϑ8ZÊ���[��0c��b�_+��h\3��:[#K��L�@�MQQ0����)�ߖ�N)c#eW���w�n	 ��#�&w�Ў۞�vK�,1 vh�Y`J�쮡/�sTu�F�Jv���oO�e49d���z?3�0�w垾6��5����J��N��P�  A
Aқ\��ǥo���A�_�Q��,&l��������Yk�v(�_�<�?�0Y0�9��8��'��z�� �4�I�VX�}��XQ��ُ����L�����q崣���Bgw��၇�G3�v� �;�УI �<�^�N�:�~��	}`�9��>����� 2k�(�\����6̈́��{]w$R�e�1D���5�h���.�i�q}!
.Ť����6�p���"Rk�i�!��5_���dL���!2X��;��]j`)i�dk�H�{/��̦=<I��b��Eh��r�F��W�G꼀^MF)s��4D�%�+�$Rk!�]�e1�F/��Ȓ��W�<��nʃ��J�k�`|ɖ��h�+g�f|W���27����ܛWL_˾>5 �8����C����������.�!���z�`t(�:Jc�q�
�4b!&����,��D͎��\�����:t��L��u�)���"�݁'�⹂`����`��cS�������!���� )�O��:`�^UC�L�����m�
�)_�J@�G1�&��ު�M����{0bkv�> t�\��5vw��`�|N�x#�R�c'�ؔ_��y�:�ϟmӚ��H8�謍��D�*6���8��4fa��f/�܈���fN"�&:�!��r�0(x�O~l�|��9hg��r@�X�r�c�cH+")~��䊬�z��mZ>���g���GM�;���H��uGs`#mن�7y/�LGҙ�n�?X��gXڈ�hh�T<]���#�>��T������y�i��4��s�XJ������ z�ә���O�x�)��L|�r�)�"gʭp,d����.�3�6
�iζ$	�w����<k^/֓� �)�f��=����Se�>.����HT��C�l��!���AV��}�0x�`�Vʃ5 ��0�o�pc�v��=�)s#R� ����,]���O���cX�h�8 �+����R�6���.ِ_�Ȏ�%�.ҵ�l�#�+}�i�R����
�����D�)2�y�% �� ǅ p���,�pԃ���Z��j����7Ֆ�5ϓ�ß�����,����!�qE�.O�9�w�	F׽����"~���I ds� ����mЅ�(,���� ��p(��H�K��G��ū���>%�͢:�TEN�\�l���:{a��-��&��Й;|�Lt]:_�!�D�@�1�1�0�Dс�ut6�L��2�L�E�nu����XU�4��d�=3��ʆ KCϵ
�f��cw�΢_\Eq���Y,И�yA@�as%�����X}�=:�w=vx�.z�Y+�y�&�3��C{M�PB�1�ѢCX�qY~h.��ڱd�^����8:���s4��a��v���Һe�_ ��h驷o2�ud���zv|�>,�թɭMD����5����eZZ,0]jufF���G�j�B���$T���BW/`i�V����\ƨF���Q�~�B�+�XB�*�Ϊ�,/���8�	y��[a�xq�r�9[�E���;�M��h�Zb[��Yz���n�!�7h�@�G��/2PKy$`�4G�˥S�����v�w�m�n[
��:�Z����U�\����X��R�	}���mCz�Ylt��稴hY�6���H�&F'�[�� �E�#{�K�ԡ�b4 ��_��]���^|!�+QwK�=��dx*-7�P�����t�ʪh((
/�{��d#<�&�`�t[���J�3�	�:����$@����:�A�3�Πg��3@�-���;�	�9q������K���������H��,���KճX݆it�$��?��,3X�@�U%�aʣ鏁�#$�
xE�iZ�������7>�yqx*�0�}�r���ۼS;� �+$�F�&��)X��X��i�ק�ܘ����l\��GJX�z�m
�f���M�yJ�/��R���1c�M�P�'|�}-��S����\�4�
d�Y`R��Ȟ�f��#_���HL��eQ�lS��Z5P�d7�n�YQ;��5Q��$��k�,�ˈ~�1{�B�J"�����]�᯷��&4M������/ J����G�ۼ��T�g���)q b�'�n�.�x��! �½�§,ȅ�:��Լ$�C�f�-�=���~ȑ���m4��S$$�kq�N��ą�����(�A�y�
�(F6�W��W�zZ�6��]�K6{"ch������3�M�	�S�un���NjJ1��z��l'�'E?
���碀Jg =���W�Z?�t�f�o��#�#9ҿjb�x�l�C��?�,��y|���3T�;=�g��g�ܗ�u)��	
"X,�,�6@�z� "� QyO���8��w�4��H�ґ����g^B��ez���:�_Ѧ._� ?aO�I2�ӭHM�kQiE̚����0J'��W@��~V���4��iy�Vؑ�2���.mA��D@.�^��!*dKͧv�̸D�PL��x8EyV�
I=��,�IL�!%��i-e�A���`����2Iz�����h�I�x�X:7z�iٖ��6
��'�u=�����XS��ìEz�בR;��'@uI�p��� }���l�4�X���f�RA4\dV��q�u{�{%������چc9���ZNr嬥�o�՟笌�È]�\O��)7fa�:Q6���jM����Y�`���tcd��+��@��k"�/�Ҡ�(*�|�PT
�)��T�7��둸5?;�,sگ4��BX��MI]�D���&˳�� �����m)����k�3�4h���ogU>A�Id�Y�y�/HL��� ^)��^#o�t+s�$�-�D΅����mwR�j�� ��`�2?�;D}E�{i��|�Vg@���뭥��� X�y����[� v�)���,a�aB��TH�"]�nesR���š��d��Gjk!h��6��)����#��%�V��{5����v{x1��m�w	𝌣�*�,���X޽eMs�0��뗫�Ϝ�{�]�$$C7��n-����@�*&�r���Q\�F��kЀ��6O����;g���Ey1�:� �s㏙H"[L]���Sqw�?�FZ����+�p����V@�NS� bU ��`��W}K
�S�i/v��堯u���Z�/Uu�!�i��1�c�� ��EpF~%#��b9a?��d���2��z�j!�ȒU!|:�f���ٗ��/��p.ү~I�������%���>2dK����X�`6V	h\?���a(��l�0s\�[D�C���%}D�<�� ���<�L��������ֻ��B��?ٕ1(L4������3}��^R���Ir��4Ͷ��%:�r�� �ya�W2[S9wZ���Q�.N<��ق�]Hm��	��3S���i=[i0�dE0�k�?`?�^,c�a�>�t��c��(=;������M��Ě~Y@W�0��6���B/��d�-�ıJ�>�`��ÇΦ.iI�?�J�b��ϛn�2ֽ�#/�
��q�bd����� ~��Pz#�mM;��'�0MW��/�cd�}��D��'�u��[�Rn�;���>i�� ����D�*� ��d�`�% �`�[hys,�������g�Y��z���!�5��_˹j4$�~����4wUIRR5�FN�֮�ү���������c�l]G5��Me�Q�`o<'����{u�~� \�����#��{_�UR<��$�M�	q�Ǩ\��fF 
�v���	�Z��d=k5�h�5 `}���[�k�}1�w��Kzo�T�N*��v<��ީ ���4[a4@�dܹյq�R�)�
4 &�uR@����2p��������n�>[��O�W�#$�ٿ�_��D�N����]1�$�������i� ��:g�'P!��\4��+͢\
�	��X��Hre�|$<��Hw��_堒��6�؃"{o��Me�yJ,^�f���3�]����fc�s����x�y""�#<�5"c�[2]ɵD�;s*ʋJBj|�����@q,�
��@�'V�)|
��ƲZ�j,c*�-�'����/��R�M6hP	�=�9�S�U����f��d��5�^R��r|�&��G��،�q"UF�ܛ������r0�&����&'! ;����J[8�r*+h8|u�O�
�����.¨4�!�$�v�Fs����X����-?���/��j�o�yR�x�}����@�\����w�媨*Gm �����a����P$��cn�p���RP�'a�Kx����<T�Sқf���[�;�*��޸;4Lt$�Lԗ
M�������:N�n�bw&Z H��ڴk��@�>���K�� ���(H]^Δtg�:Ũ�S��p��KY�Q�h�Z�\�J�?Z��6T����s�Yތ���y��P�1�bB�i�Y�&�1���_Is<�U��h���=��U������7*^D�s~��}�@bY�ߨ��%OM���+�Ok�`Rͧ�N�@���[L���g��${�R߆�Ư��U�[;j)�@���P���[�o�����F�_�϶e	���LZ�s%kx��ڶ��6i_�B��%�iۜ׬�b���j&�w�T���T�1������g*+� ���\��{�+�g����Ĵ\�z z Y>c:!f|B�"W+���I1�v��zx������<��4.�p�k�\����}� �l9�R'�STn:\v�H.Ō�@�L��"�|i�Z4>�A�0��V*۽q'���6��||{�$�(� ���<�uJ����bCM��|���s>�0�k��{�/B��V��0�@��&(���&O�c�����;{Sp֗z/6z�A�K��3�x�1��\��������/�U2��t��?A�\H��,�K�]�a	xK
vQ��v��_[���:(Nd�9��ct�%;�����	��hLhai�����sT���(�q�dIjM���r@/4���;'.��[N��%%�LP���I[�a�6L�G�NQ��kZ�Z�nvi�>��,�j ���*z�(�v�
8uYS�&_t�M��G	*�Q,\���Ru�b���xb�R�//N���WM����q�Vm��jM�_�"N�xx��X�ǽ�D.��2 n�5�7�?��t��!phw�ND�3�^���Ie�
|d�I���e����L6M����`��=F�h�JX����s�=S�d��ud�Y}�'R��>� t��9��N9���TRF�|S�0�7WJ���u�7�K��r*F"�biq��W���>��<A<x(O��I�OcP�;�Q��o.}��6\ף��#��������ި;�B�H*����ˋ��	� ���8�e^�$��Q�?��:}���_��&�ۦMޞ��Ar�UI c��(a
i
�ܷ�LZ�~>F������	��F��DN�>{�Ӱ���߬]�J��̫pQ��~k�*I?סm`V��{��h��(���j՘zh�Y~þZ��9@W�݌�ث3׹<JdZaJR�'V��U"�b).mӒO����z	���.0�{\s)xL�Z�᭨C��za+P=�`�%-��t���c���TF{��>]Y��������WȦ��S
�]IݶL�e�@V��Z�T��pr�������>�T��} �pk]���$�uL�ZΙY��g9a�����u��bE��&Qʰ��g��M�8��h���lo}�$��~�[�M[�c/�I�����SO�S�5`pZN#�����o�N�_�B����]��;]n�'0�m�y9�Z�'V�M���G^�X�hW+sw��5`�rʝz^��~n�.�zlC�9H>e��uJ����Z��^���Dj�
ݻ]s���8Z�u�o��5��~������u};��W��	O<�Z�*�y��t���n�g�KZ�y�`f�mL�$�����)�S��� �윞0�0 .���`�^d�e<�Xh���M�#i>f�{q����ѧ�\h�1 �}nsۑ��y��L�Θ�O����ǒz̗T���tz:�ّI���!D� ����E��<�� �gj��A���CD5���cx�_�?ۈF��&���`Օ�o���NxyۑRb*�K�o�q���?Q}ß>��>P׮����2�Z鍊�da�=���Z�`خ��X�!�h7U}�Yݡ%�Д}[B��(��Dhy-0�#�����5�<|�+>_P0ƍ)q��7�2s�L	��o���wg`����d5�|�ǜ[� ��J���h<�"���/S)v����z`L�H��9��H��Q�?���N�J�ws+�̕�<�3VY�����"���Å�F���s]�T������&�\��b�n�%b�0��P*��<�2�:��޽��B�N�E��b($�O���l��|�*����v:N;��\R���:2ǭi�Uſ���c=��՘f~��Z����+����S2< ��{,��BqR)�d���q^�t�i?�?��ӳEn��`ѭ!����`�d^� -(����¥Դ[8��0���xFZ���9��aq���@M�����>���)gM�L�{�7ԑg�oY��3�G��9*�R�ڿ�F��o��q��4`"�ǥ��_ղF�x�[U0����E�AYgTݿ�L']�
�����60�I{U9�n��h��d�*�tdJ�D���Vn: ��ѳ�c+|?T�>f�~U��ԧ��@�*)GH��wF�0�LZ<*Ŏu��n�Le^Ni�B�?ָ�d��$=��ȗ Of�#�u�=�m�&7�7%?D}���\m'd�1�>A?�f����VD(JX&����P�i��3cbxi5
�z�}����.����������3i�=����'��Kܘ�/�U�����%	�Ƽ�C���P����#x����;�������$c�ؕ <{9r��%;��ukbH9�Z0�HN��g�����-J���bڀ{�o#��=����`��b��Тg.6�/�ޭ�`/��O遥�[�p�#H��HzCE����p�m�т.�q�r�O˻�Ȼ����(��H�':CD0����Ŀ�O>.#:e\�$�k�� ����ρ+�OTL:#l@Z�o#9G��E� ��3�w���w����V[>��V\�m����`=�g���`�`��z�Y�6j��z��1ߠ�R]^J�[PA�$O��C��w���*���#Ug��\��L!�oS�x��s'����b6������������=�>Ҥ\R[U�C~$d�>Y��q<.����*�.�$���� U�`�-�}��C�m�-k<��WQ�S(ۺ[�K�K)(�f�˩�@��=�����R��iC�I��}�*,r&yq�hެgqX�X�F�����zG�'mw�����s���s)�"M��Z��^I�YaU	��jV�T{�FO��52'dZi.�"ٷ�Əoá���0�Lz�����|�]I�D��($�z�݅�'74�q6��jw<�&uQ�n&R��bf�L5�,�e���,C��l���a;�Q |�Q��%���>��M�7DO�\���č�Z�#�C=F?�?�G��"�i���-	%'�1�A��;P�e�Ei�k��鏨�e�7X�̅9�)Ҧ��Q*�
�#�V��=:5n���[A�̉�E(F�]w�
&������'ai����4�r� �L��uA�|K7	�Gn��6<ܕ�w	�$@@sM�ɞ�DB��9t�i R�ɐ]�0���a���2���i�krT��lWH�-M�zA�SevA��Nx
��'6�=<��9]W����q�1�>EW�iEG��oX��m���팠F�޵����L�$��U�o�;�t�����Q8�ج#A����j2}����:<f����h�N����<�R����M����/�FK���@���_9�u%�5���V]1�8lm�l�"�$C`P�,�L�#g8E��_��	n��x`�y�qT0�y˞�闎f�Ũ��RDRBsP\:��E'��7�O�ѤRb���*$�'Q�	�p(����*0��׾4o�F��<����>���*ֱ�#Cy�秹8�!.+�(�y��D�g�nf���[nJ�_ww
����>�%	�2�X�/jn	� El����z�Sl;D|u�j�[�&����%W�=Va�Q%m %D�Q�[��l:�������^6n!�kҧ��:��D[���Ѳ�y9��z�hh�����EޢM�d�hj�J�%���{/�FǓu��A��Fȡ
�U�/����%=�V[�����y�A�w*�g�LM���ED7'W�N��*���wӅx�IB�L9��__z�g-]�Rov��-]n�"�jX|`,����l%��޴+�څ�{���#دj*�<!���7X�#�y�
z0/s�	��)�����|�z�_���W��x>["�:
t>����/�'��ij�<�AT���B�E�0/(`�z>�8�X��Q0��#�Б*�5h�z��i1jB�9U�P�0f�
-1U��B����^��I��{���uOlNAm�vދ|�����^8gj@^����.���k�+���	�p��<�"�g�7>�'3>	����X���O���ӡ���G�i�x �R��<q-v�\���ߙ�� 9��Iٕ����!���w]��FD�� En'�B�"��|o��uI�*ݣ��f�"�>���y���b�|��>����F:�J:�D���L��I���_���9ƪ9예[4� }��{�,`�*%?�i���	���>��,�����u5��$�K�Ά���0����M��`' X����qR���b*���Q�QM��!�D^�Y�hV�*xln��|��cf�8E+��)C�KY.��ϖNp�ybγ�z ݱكq7�8��("[1\�xU`9*���kQQ���T��c[,�Ǫ��	$���J5�]ʫӞ�©.�����`ӭ�3�yR����B����NB^_�S�E���C~���r�]��|��Wr'�;8��lP�}'�n������`Bϴ�cH�X��G?�,׎��ܼ����)���z-1f��ў��\i��/�ݛ���Y���g�f]j�1,�K_@S�։ �;Ɔ�G� S֥�`94�=BҲ��υ��� �*�8�ޚ�+�<,��&v*�<U$/���y�9y�׏���h�f�r�J�<IT�\ f	���O��4�s�ǣ��RX��dH?��;�#
Ϲ��:z<UM��XOL��0T�fї5ƚ��m��E�Q�
9E! 쁄-ǻr2>��ێ�\$Fu����1|�i�ٔ����"b�j]@���3��G������G�Y�o�H+�)�&x=m���Ο���V,�_!�ɾ�?p�
�QMB�"�]�c��ú��g9ȫ���V&��ӇZKq�f�:(�%B���ۻ�H  u���k������(�� B��Pi���6�ч�1/E��
��+��^���@RϺTҨ��K�~���U�*���bs�0h��I(�q^	�H^a<{�\��OՏ�"��SL�f�bSS:�"};��q�����ľ���Ł;�d� �އ"�ӵlS��˟���rkDr�]/�/�������f�f�`����a��k��|w�$fq����N����K�hm%��軤H��RS�.�ܮ�\gcN��] �+ȇ�Rx�7�����S<��\Bk�&hb�#Q{�b�e3#�F����_�a wD��@H��y�֑�jݐ>N;��d�8���R�w�^���r��s�E��p?���3��/��퇫5�q�P;������מ#�Xyؽ�?�w7�CO		}"!�]��?��d&3eKL~���փ�sL_��AC�^Z&���k�?U�~/ �Ϳ0��u�g%��J��y/[9˦2�o%[&��"�&u���C8�k������k:S��>v5UUŃ�R�2S�&k���b=�0 ldz*���6�N��O^���x�|�-�Z���.:QĲ�Ղ��X��A���	/��]Vm��Ṹ�(��@f�!�B��4r�Oݘ���j��&�H���C�����_`�8Ń���� �}�ӈu���i��ԼT�}� �'��	����-�q�%�{%�;��EA��D�5��>��	i��XԼJ2c��H�ND:�7�]b�"� 3�����6��%����9�� ,���Y3�9-^����C�c�m�F<ǁ)�(���W<&-8v��\vOzr�, �
�N("�Ip�3D��,k��i�v��M����m,�ɼ��������d4���јV��u�R���.A ��㓗-i(8*B�<v:F;����嫰*�m�S��rB���c{m�Vq��Oq�Sv�P�;�7����G����_<�s�a����ʗ�G4�ę@����'B�ڧm�M�@e֠�"z�zyε�{O7��<����8<���@?���M�`:q���mө	Hfp�Z$���h�^�ԋ�!E�=d0YnV�8��إ� ^<͜5��2���%A@gT͙����"&���e7�k��qj�9�xv7������R-�=��-�j�mw%��/�=�sκ:=�[�A�AZ��Sr���n����~���?t�m^	����S�~���!`���j N���<?L�%?��y�}Ը���&9h`��u�Y1u��Kޥ�����Y����ٵ��a��l#D�0_9&��7��m��X����>��-?��	�+ZV�[�7���6	�P�Tdb3��K?��U'���!#�	)�:
9�脬�2�����ґj�/*�1��<�q�r��E��K���H�
L\��¯υf�9y��R���g�O	:~O��G(>\�9A��Yc25U�n ,�Ce��oE���t_k�j.����Q����K[K�����Zy�(�bc�j��-ҡCe�@&ZgU3Ý��-a��z)KQF>	w�Y:�s�B�xF��'/h��Y��d5Q�=/΋�iS[qjl �<�߿�gؑ�Dh��ܩ���8�fٕ���Q��@��rz�J����@�*C���Sآ�H��CnT�o�`/�N8���uBI2d
z8��j�`qao��v��_�٬!�7&5՛Ӎp7KQN����W�=c���������ct��wfK�v��ƌm0'7H:J�)�m��X�ܬo���d��Uc:�arh̗�� ?��n����-^�#�MS?l�i��}7es�B�v},i� �����C���-�"G���J��\F���e��%�1-�{sL�GT<;��\â"$�?(��1Fd�t�����א�	q�ڳ8�궥ʍń�-_ۍ������O�j�����5p�${*LW+��G/&��xv�?�\;�z�8���!��_)���k�A^�6:�;�\���E}])y�[&*J�Gp=�ޡ5X>����rbu�0��^7�(��y;zK���Q!t`�e��6BAǯ5oU���F,�!ϯ��<��7#�s��|!�pG���H;_c`F)����7ց�XF4q���B;�v�����kO�/���� ��] ���͌�Z��
�`ꃄ�~�����gA^��6�,��Sz�wC�)�#�y�8
e��j2�M��J;6���V&@�K���@a�9m�	�����*��-��J{�ٲ�x_��1�c<�*xYǖ�
�� �'�6�tsO�T�;�w��)�9s�$pځb���0LϮ�R�,��t����k��yP�D����}���_��3�H��I"�d��Uu���ոٱ��}j�6^teR�oҞ�&w�!4��x��\'�	3��w�Fd��J�$�p:��� ��_A��ҷ���O��7�	��l�d߮��J���zH�����Cu\����Ŗ�G��a­҅,� R:#_k�23��s�
�������[�����z��ƫ#�r���"�"I��jΈTG��83���v��]���@ߑ�gK�W�cd��t5s:W���j3R*�5Ȁpl��޿�����n�Щ�X�Y���C�މ�-p�]�]�4��RVճ{�a�P�ʋA��������u-a��x�M*�����p�,�|P_R*�Pm�������*a���ej����	����FF�����f1OU�'���X����������7�MEU�'y��	��*MҨ���-[o��ۆ%wFl/�нYc�'S�	q��j���|v~@�:�k�r�*��מ��k;>�����8� _�T���%X�S��b�Y���Oq�8��EE"d��S��L	Z�S�_�VC:t^���o֖f�M��$�a}�~aƏ�����ÆA�	�T���|�5����7m�Q��(L#%d�z��S�T葡~w�Z�8s��(�������0J	�wO�-��C6&g��s_��jx:*���p-4��bJq7 �"n:�;�/R���Oϼ����_�����������t�s&��O�Zm���K�\0H�C�~I��%�f��������Y*%�y����N�	<�5j|./���2p}��B
i�ܸ?��"����c�a�h���`<;�!�L
���v不Y)ϵ���XTu*�����N�k+�X������Z�����ݷ�|\�.���|�3c;����-VjF@e;\�D�?�x@J"�;:v�Q�_�%d�to@�U��dB�^h�*Ӫ�>��*�&_=��xBPZ����Xp3�A.����X;� |J��D�/���3�� y�(�LN��vu�X6h�
���Uo��5�NA����4LWC1"�z_�)��eT<3�!���0R[}f�΍᠈s�&3rN�Z�h�B.�t�L@�'G�̨!��w4"���3�w�+(Ů�4���4��w�I�
�ѓ$�o����yFK�1Nq�������9�L����U�����9�/�2,d/v��e���F�{�l�J��P,�5e�gZ�]z�up�N��c��>���c�(�e�� ��׊_R�����C�z���$C6D����	/�-C��Ёfo���F>���.p��l}z��� ,GcW������ ����N%!��%Z'r��bppIO��OFI�!�4�և`[6�]��1!�ԳsD*JHU�R�̳+sC� 	m�g�gʏ�K�{�n��^����,k���DxϦ�n`ڥ^��ט��[>�~Py�V���ꎘ���c��5vYkN�_z����0�;���d��z$��u��i˷}����yRt����|}�g�.i����4ZD������9�5�/ ��H��������Ȍ��2����݉��"�(uL��#�$���,��G��:��ʕO�6�4���WQW0.�>o`���3�s:��p��8����&!��3�>���'�|x���"rY��t��-�lf�vf�O�z�RxG�:�y��֮D�s�u�po���3���sl��������_zy�������?�`@�Y)�"�^H��I!]�cw���U:B֩l��o�p*�\N�nF��i~�+]S%��_��>~��3ƓO���![:���T`�B�����J����~����U��t�@>s"�S6�,΍�"�`��W���z_b�
��i2�
�E�����>��E��/��b�o�&OO�m�0`a¾P,+�Z�~���Z$9�	A܃�Y�s�F0i\�!�r�I��SI����m�m����Fu�ۥS��˵�=6�����u��Y���"��R���\1	R�@��6����c�9���#e�0�w ���ըR6ы�1Z?Є�A��W��}:ZӅJ��+	ײ�֎��PX��~ŭ@�H�}��KjQ$�c��g���H���P�pܵ+=a���+H\�`4C�dQ*F�K��"v�0s�0$g^ܬ4�Z��N�
����h|y����Ʃ2�����Ac�d�U�3����ܲ7�i7�Ih���jڴ)�4��r@T�գ����e�}��\��i8�+p����c7|����N�����I�����3�i)n�|�.z/����~a����%�D�1=m�.�}�e{=��g�=��L���W���si��T�� ݠ�_��a*
zjO3dw�ڠ�B8��F��ۂer�V-�+���k����
���fe�z3P�<�5�
� ���| ��Q_�Ko	�"�����Xn�s_��
;����D4��[��͹�;��$�(K��m�%%*�8���VK���\�~h̵��maS�4F������ˆ��BX��RU	��ZPE@�%}j�HHm�[pe@�\,*�pd�q�y�ce҇ |R����:*m}ށ-���g��l�X^y�Ľ+Vq� ���ۉb����u
�^�Z5�<*�T._c�KQ��g��9i�\U�����~vv؆Uq� =��b1�ݓ'�Ϝ7�6���?���՝�o�[�q��i�s]&�נ谶��;g��u���)��,�w���9t�W?2�;��)X��5�l*�36�;�2X�FP4�U���r��BSءq @u�䳨�<S3�/4fQ%��UU�/�|d�ʿm-C������6|�7�v��~`�ܜ}E=��f	*5�	��4�ܬQ�������-�&�4B�����Ö�3P��ˣC���(�����Qr�]C$*��\��6I���V�������<#O.{�M
�R =��l��c8eW�,ׄ�sl�Ƨ3I�ɳx�	�\`�0�A��a������R��`)�ϟ��bY	Dk������}k����E�i�bT/�5 ɶ=�}����)?g�+���[�"�}��2!ϔn������ސ�4�	��^�b���b��5v_G��Z� ���ӂ�qvH�/���3_,@���;����1d�[���=7���eG��ʊ�vuo�=ۿ�	�����D҃
��.ۨ��^ے`� "||8|��2������/q�4���`���
�eh�"e������g��u�G��zb���ɴ��H���,y�\�#���P:�|N}������/��-�b���Q�0�kl����y���Oa�no�T�"� {�Om:^���#�-c6�f��a]�c��[�#ׂ�
1K�K�~�M��K���7�)����лR�J�ߞ�F��/�`6��ao��u��av�|�A�.�?{�7n\tQ�UyF��Xi Ҹ~M��z%�p\��f$b�{F��_H�⤭�$���6c�8!���_�ҝ��E�ܘ�@Z�ڲ��c�#�O�\+b��aS��Mf/�j A��sL;�bڍ?,�6?y�Us�}��N�r�,x���hUu��Rx�L�&q؏"��!�7��Q4!sٰ���*�J*Ź݁'�����ә���Bߙb�pCE��ʉp�~J<9�7%�l����ɚt�S����kZ{��}E�4b��U�T�9����)	~ 96�2i�a����N/<�ɐ���ԲT!�k�+���BL^�	.EO�Jh~��5��J�(�g6�V��6��]qZx�n��w��s�e�����m��:�	�o�-�ߠ�J���غ[_p�^�p����n�:pUl._��NMZ?_{��!(��}�A��_/[����9�lL5�h��B�<��S���h{���i5~�LhM�Cč�n����O��h�:��c�k$1S@����E�*C����&�5��\?>U{	��u�P�ZV���M#�~?�B������yL�-!��)j�֕��+c6vI?�s;W	���j��50�]��`� (e��r�i�|�+A��+X�>s�L����?cy|]�i�6��MV���Z�����gr!��Y\bT|Ŕs��-��6uu�e|�*�W��@%Ӆ����c��C+�`�Q����oS�����iu������	�w�!52�WD�{a�V�@�"T�o��^	=y`-αxR��q��E�I�ȷ�4��ǅBz���y�����<�-Q_����r^Bdъ�K'��9ާh@$�@��>���ҾV,/�[%�I�GP1�u���p~����i=�>��XH����P��\���7vM�}P ��G����1�ȓ�ˑ�꯱WJ���V�F�P?��Z-�؆x�j�l��*.�T|4��I�]�	憀�O� ���/f������[/ONYa?�G�E4�� ˛�����d�t������H���z��I�:�Q�lԗ��M�ч�r�;�~g�܃��EbٱD�%�':!���ӯ|�8�SK�'ʀ�w~5n��Թ��R32AW���<�Y���"�k�s��m��������?s;�͈��h����DR}Xw1�k�O��h�5�iRމ��g"^�1 �j��p�{-d�T_\>?�f�M�0���|��HHALT��IP��n)��j�+��qE���Z	�m�����2Ah-I"I}��GYq����^6�g�eG�j=�S��s��į@�sE�?,Ake�$0�U<n�܊�i o�3*�O���<���;�P��;��� Ef�i�	v�Y�'lv�5�E兣�����Ma2t��_p7�]y�����5�1i�(yTw�OmF���=h/g�B}>�eJ�w�pw�b5���8+S����������:P�� �Z�9	�ζ���`C�+ݼ��n.��KG�v��b���	�n*�|�	{�T��	��Ӫڊc����m�R~|�2�4�uU].�'=W`�Z����y2_<�FJO����j��� �ir����В��uJ�r6�ui��.�4�KW�rk���r�y��Qvуn6�i�x팂����� {����j��5��<"��
]�Z����AF�VVZ�f�
�Q��/ �Οg�Q��Y�۞�H��J)�j�&������`�j���W��il�edL#���W���(��9�6�kD�Q�D�܊[�����֤yU�'��]ѻ�A�|�wz{Zu[A�l��yM3m��i��1Ø�MaS�\OZ����:P!�Uι'R=���}?�pZ��Vs
x�hŔ�"%O ��3�-V[����3w�x���LQ�ͻ�>А�]Y���Q�r�{���"gҫҏ�b-`�,���a"�o�_r�㩕gpw�V��I#�s�cʲOA
\;�N0PY�"��S�"�a_��3���H���k^v��Xh܂�6BY+ﲧK���>�S�S�dZ���j��~�P��2�UB�~c6>} �nW|K=������t�N�xln�M��5�0c)S�*ɣ�ky���? �9G�?�Ѷ.4���nOyP�mٖ6�@��*�!9����5�"
$���-��������o��A4/�)6fZ����|���7c���t��-3��e�I� �M��?Ѡ����g��4�}$��e��,�ph1��@qO�ڼl��ٳg��3賏iznx�N�xŧ(��\�a�L㿌��`E8�I�Zg�5lt��-���Q���D��G��`�q��yb��E'�ք��6K�Qx����R�*H�����-M0G-�-�#H`FY6sC\*�V�5�����<�a�>L4�����U� �K���x-�Ͽ���	g�RQ���ys�0è�	�u}G��d�)Á�e,m� @�A���OA4 ����&��XؚΣ���~�V���J59�,�>����;qW^� �_�{қ�2i�Q���4Z�0K��'Y [:[�	���g.@è��v%ȸh�h�P�J�geм��K/�Wl���t��T�jcy��l;�|Q�g�4d^��c#ľo(vk:_���Y�����Z��r6��'^�A	��}�"@;)�P��9�����S��G�^��U1x�v���vҰ�#
Uɢ���#��F.��4P�s5�F�ҼP�٧�v������}��ɚ�>�w*�6��!�<�0��p��?=�W����WMoO�irD�؅oZ�	���!+�1�Ő`��{_R�Έ���	���b�IOV~�*߲�i��2�ȷ�[V�Z�z~nJk��)�V�W1��$~:tj����U�L�gS�|`�|ߙ�}��9� ��@7U�n��;E��F�/��7�$V��������=[.sat����,�Ǽ��Wx�c��kD�H.��K������bd�ȅ��+�腆'����_=*��2����(�C�:�)�Cm�p����@\4�g�~/�4�R�I?EF���a���EZ�&���SQ���Z>H6�o��`���y�?c��T��>��C�ĝ5O�ͺ'�Н4�����
C��`���� ��w@��$�J�|���)�Y���ئ�r�*��G^�fR��aF>Я���3�&stX��H<���g�/r�|&�;�jv����A3?�̊��f������|ɏ\`���"{�X�)�j�:���s��,�r�,0s�g����
ބ��_V���؆w���%N�"g/p �\s@������?a�!�*0l�+l=B2�N$�Ǣ��@���1�_y���L��E��d{��H�BWҎ7g [9VI<���n�����m�)e	�_��퇸x;�^���	>��&{�5�};���	�6^��`;"a���
�Μ�/�n#�¯!��]��Rv �m8V��>/U�]�pʽUA�h�d��}���,�;�UD��e^y�����^��*�밢�[�]� ��W{@:����!��eU�/ �`ʳ� �+�"�c!֖0�([K���ns��ZG�\����Xr9��'���ȑ���O������l�N����:�h	�Q�Z�7N��,/�F�r�uK�~�H��w���ry�>FQú �]<��5\����ub@���/�	�����by(6��'rͦ���,�*T�t1@��"��5F	��L԰R�Ev���}���{��Z��&6�+�:b˙���Z����Ý&L|�t<M�Ba�@EA������x�KC;e3n"\'�y��}�4����߭�0;I�d�ыh�� *v7t0h�p���4��mX(g��aJ�ɳ��?�D��M���	5�6�7�S�>6��R�8�׳��*��0f{̼�᫕D�UNݥ�=��5^�%��]&��"�B����i���M��tU�C��G��"J����f����tWy�ۄ�J�q?w@�H�g[";�L@����@���ұ+���'���|M(���a�d��'� 
����%Y��Pw<.�������|�t���o���H	�`Mt]��loߐ�Қ=�C�WT��{��D��֦��ۂ0���K���7�5~�k��c�/rsi��FR�,��4d��,:͸ 乷k�F��F���<"���#b!�''S�``s�d�� �E_�8�F�s�j��z�6pn'7�HY�	��I�a�4�1ݖ�;c�G���$-ZF��5��G+d�Y��
(6.(��#](���!��>�XL�9H&����ã�y�e <��P��z(`2���Y0am~���>+��N��%���
6��?�/"$Ғ��4���-ِ�w�k	�u���g�o4�%�"���*β�w�J��8 �v�%�C� ��E����hwܶ��r%��>�x�'��	�1�ۋ�;Ө� T��N�/L�ِ�KF��x@7���d_5�3r�=�JpxTu��.[��/��+����<�D"�eʿ�����@KU�q0��uѸ��c�:J�4�L�����᷸OZFo�!�T���7#���e�D�'w���ӎ��]I���t�[Z{兩�a�E&��.�t��R���j���2��1�< �	�(�Y���ҭ�EE�����݇��H�Q#{�(��?�#�J�����Q\7�2�7,���\����{�����Z�ˊ���-�>B�
�B���^)H�O�-����t�:M6�c��蝝T+$M'.1�[�-lzM�l�+ք�ۍ_�d���gv����'9��0J��[�Zұ.Q����s"ad!1���Si[pI���M8�~�ϚW$t>����N��AK_����N�l������Ж���<��ཏP�*�EY�'<�M�Rb��X��ͶT}�1�/ڊ��!i�kr�c;�)'�T�������KXv�/ٔ��s�ܨ�9H'�X"��s3��e/���
�Xw(z7w&i�B����پq�x�p�bv�y�������-���{��ܶi�ę��RX�S��L׳=i���LXf߈!]�o"~�z"a tx3A�t��bb���� �\`��h9�0� 7���	{�nMl.�x[���tc�~�Q��I�A�F��A��ߑ��<�����$���4(�ޣ �1k�3�O�[ŪZLl�D�QwLd.Epu˘�ڥﲣn�`F��r�}��[�+�M����K#ڹ73	cl�⨴�D��I��O��z���^B�Ъ(��#���`S֗F�?�(�1���"y	�ƺ�T2ϳ�bU���H�G3k�b�c�ɍ��{ �-" ��_���B0�q*%��ant�|*��SV=�`XYfI� �,���=�v���QS��i���W�`��З�l�vm=I��+֧;�bXob��v�Ma(;�yK^� ���ҁ��3"��>7Ȁ��	G!�?L=�_�ɒaye`�)!��9�׺��c#4�##h[~e�67�m��g��)�VE�<1�����~x�|��z�csV7.2�ykY��^ޕ�h�/@�'۝_J`�p9�+7�勂0�PNz��(H��O�8�܄�{����Y���-�J ݿzwø�B�ɦ�(dѾ z�����)����	��A8��,6Nr�x;�5���W[:�b)��hB��߰{n�w�'�@@*!�y*�aLD�K�%3lP#�<����3R���[��#�s�Vy�8�4ӝ�=d:�ڶ\�#<@&�M^�@^�Vj53�gJܒ��J���+�J��4�jI�Z��d ௺�Yk`dz\��t�4�!�Y��h��sd$g��ݠ���Qd�{ZbN��� {v���~��Fͻ��(�R� ������C����~�G��럕d��w)�Vk����[k�M)�<K-J�@ڣT���>)��<��;z_�6��Ħ��k>FC�Ƙ���3��:\�56�!\F3�:�E
G�٠�I}:(hVj��,�uY�H#����+���7�H9#�5j?G���/a]�$���SM�4\5����jό�fS�T$����k,�z�\��R������Vjv��洉��GHZ��D���*��*DktbK;em�r�c�Ve���`$`����hic���RP�G1��h�ЗՏ�r�[���fu�g���s�����vQd4MOW�W���$"��&���^�{�;%6E�4e�94x�L�>ƴW�*�����˳���-CQ�?�f��ЧD�}���\� mz"�v�^�*Lp��H����@�7q�D^�w{�;����e*�����<��Ӄ xI_*\E�X�Z(3K&L��B����k�ȠVY,�����
����:�p�;V~��:ˋ���
�J�o1�˥!�kҠ���QQ�dd'�
�F�W';����+dI�+ N<~Y�uqǖ�QN���y�ni"&7{����پ�0C�+r�sۨ�}�#~v%d\U�]�"������n=�D��}�[��b��N�Q^�AF"��K��H�X���*p�I����W!�,7�F�w ��5���KT׻�kn/��H_�׆�G���0Ԏ��Ĥ��H��є�A�6��_,�6� �O?H?m���^ l'��l���85��T'�Ĳ�)�	q��&yb5��/,q!�%����y(�M0����j��DI��uk�In� fd�1���="�\8Y^/��8������nK�'�]��t�Ӂ��SG�s*2�E�.����^�8\���JXϡj&��,��O�s�_��A���Arj[MͺS)L��2)_�[����4�
 �υ�7����/q�f5��B�X��i��2���)_XI�U���8����V��6�V�=��3H\%$�(?��E}��U�ouE�����O|��37�`2�p>ɳ9�/3͏Ԅ�'�������~uRT$��_�ZF��We���ؕ9���h�k{j��]'�|��ɛ�~|�Ѭ�A����l��~�$�Ffb�`�fT�}d�X�i�ֈN�\�3��	���h1�0l4��8�%E�U�e�k.8$Φ�����=�7�8V�ҽ��6�Ȝij�2s���\V ���{����13�V�i�I����� _�=�U�lb�@˳3va�d m���һ�6���O�&�30�=�݋�ßAp��c� <5e�iΥB��Iu��;E�K+�~�/���<��h�U��7ʷ��xx����s20�n�)��3LAm�z�pv��q���vQ��2���U�ib�����+��9:��8�Y���,w�Z�A/�TIq�b��r�"6P�xF�E!O!~�0�yƣ�T���̧�����L��*�� eu��g�;���L�6oW[W�-l�ǹ]3xBL���t�8�,%���@:锅���Z�Y�}��<�޽�PK)�dcQ�R�c�N3�ɺto�f@����xZ�5�����p�a��_������	0���𵧝��/"�(�1�|��3U�_ށ��{�!�x���9�� �αV1�u]`ᓶW�D\;�n_;�"��b��W��W�>V*vv�5�#L:9'f>~{�u8{#�0���j���ՓT
W	"�0�[v��eh�5��y���o��(`K��ݓRZ�Ew}{�:9mV)��`7'��	�������jPN���(���m)z~�\���̍a�ڷ,�70�Ēd`^�.(8�+���n����dy��M�����y�Ίu���"B$h��%���w�čE1�k�T]��1�2b�Ep�I>�f����4���7�^R��Q6܇o���1_�ԣe�_%��zx���tʯ6�o��D~:��?`�����6�w����_�|���OE�!P����K�'��fQa���UW�:o������C��P�����=������_���[�����Y��s�y/J�ԑ��ؙ�h�$�����HL��m,��}���A��it"Rg�\tY=�}i����dʷ�h��̮� V�G��������c��}'��j������ T)�f���HY���M�+6���VR{ߨ*��u���fd�%فV�u���¢��P�+v �HK�%��,��j��E*>�;@�Dbu��4����i�Nw+j}��;Q�����I��ɰ�?ۏ�%����U��X�u�G��x����[c�i�����s�>|E0O�U�c~���I�7u؏�
�D�n�qi��C�=Fvx��*����qZt9�T����;PܦK��i��HO]	��=���4i=�HK��u������0����i5��w{iW:����je7�P�=��ulد��<��挘b��MM������=�2!g���� �o�����0�࿆��H�Kfk�������wc�駕�7"� ���M��P�"��	�1�I_̻Jwޝ�]6��>udA�V?|�a��ٱv�E~kI�&裔ca&��c�@L�K����4£[#������ЃPh�k�\x�����1j��^t50�U��sx��]^p@~2�N����+��ʃ�ر,�� ���A��Q���{�S�8�A��F5QClnc�\����O���x���FǷ�ڟO�ő������Ef�a����->K(IT�x���yGO>X]&QJ�.Z��îY�
��Ʈ��xXo��G$J�GP�\Q�r��%�����z��-��>E�;�-KK�<�= tFA��eLJ=n������c����*|���Qa*ō$�1"��ؓ�i�ބ�rc1���+tgT�x^�_&;��tAUFF
�Zv���������`M~�"�v�s� �C�!Li2���C��2�����ہ�!g�*|�5!C�H�DɪT�g��g�u�ϰ���7e?�+��W��̨*��Z����2�C����=��v����kBRW�[r��v�~e���0�3�;��^���
7d���`�������Y-O p�u��
�ùw�_l���C���~�]���m�*�5h�4 ���%D\��P?��}#Y����C�ONw�M�k��݌\&��O}�z���F��R8Wc{W��.�v��^��~eW�t���ͻ����:���I=Z7��O|,�� J�u�������i��?�P�5�L��O65�4���v	PP8�n�65�(]�A��
D���}�H�e�s��1PԨ�b�:Y�k"�{�S�@�3�tP���`�h�A�?����q���f�C�E5
2 0���Y���5�EOa*VG����i'${� Ή0�����T��"س�)lgox���>;.���>O<?0��s,���|�����ȯ��R�r�ˡ�Pme;ry�$uf{3�V�?����ˢJW�&ɜ����;���@�{8��)�E��KJv��Trh�qg�*��<���k�"��X����e,�JZ���Rm[Ia��d��G��������l)탑8J�GKp޾��a�-J�簇͗��p�,G1n~�;����j(���e����^�/Y�i��=�;@{J@HO/A���F��R�T���E���ٮC��={��5���NckE<ɽp^eۃ�Y��Έ�c�L�vK�����G5 ܼ�'y]����}��Չi۟�Q�-a���7�5i���R�/V����	�7�p��O��o����E#�lrgb����m
?��np��@}Q^��ƪ�yƲ�u:�� lH� ���Z7|p���_�S�U���q���%�:�.���c�o���{..z�\�#�xi|V���ru_T�v��tƿ�96��FfMɮ�*;��=���Ɨ��у�yf�m��6
.Ę|/*T��T��%*D�,�OhjK��oW�J�'�IyE.�}C�����6�N���T!��D��5�h%��s�^�)�ȍ�NÖ�1��r�ղ���3�_CjOZ=�������aĢpF�-����BW`Ѥn��z�%�m�+E��0a�!��bi�`�C֒����o.����z�\9����X�#3�B��O��/U�(;�I�Lt�2ma �6�|��)�4� �t��^Wt��*N���������B�3����g�|e�J�M�"���D�7mjK9�;H�9oF�mت�Q�9�5��앱�t��S�C]��7��Ū����ͻ|c9RI�6��i��r'C�:�������lu��p7~:�S73-Fj�n��?�G��x��Bg;���dXY�/����ܟQ�?��<?�"��-�G��U?C)'���5P'���
�@#��9�'H������ڐ=���d�ͿTq�痮���n��P�s&z<*6Џ:aki6�f�)��T=9؇�ċ�����#��Mi�l��$�yY��'�>V����oJ� ԡO|]�|�s�eߣ8��9({��BJ>��\#9�p	v���G0�ԗ�G�F�i�m���6���0t�Q�]�:��	_ -fl�1�VY4���>0c��ll���n�>m�Hk^�P#}4�!~=�q|
p��a;3R]�yR�Z)��Lm�g{����{�yft�P��bMb����Rf��f�����\OGVe�vIvznDQT5z;N�Cd��W��v���F����ؑ�V����+��0�8/�/7 ���8s)����7hc�y��3�g6F#�땚�*�_���;�m���#Q���Y@k��;�́����')T,�%v�+
z�r��U��fDp�j�>�i0����sO�^���~w��;(OrW�!e�]�	K�H�Z�x���b�텺[jtv�5+�fH<�����yl?�f�y�vQ����o�7�px'�cG+e�a�V���m��.���)��W�UK��A	��	�S@r�w瀜֝��$no��D�V��9�F�h��֧�L�]�R� c2%@O�b�&�K$~AŽ�i�����q�q��n`��.��ν�����>�pwCj�)1�⥕Z�0��`zBS6ӷ~¥{�p�LXwо�ԧ���ׅ;�^u~nE�m�*�$bcoꡝ�o�)�)� !��øLO��)��i���/"0���r2�M_�d���|2+ē�Z����g�HP�s���/�0�s��{6IW��1�6\?��]�*2%�g�Z��ع�/��.��ƌ�c��>���<{۳�,�װ�jz��&��;6�R�jɷS1��-!�9�L%�C��M��%�@G](�{�-"�n�I�OV�-'8��U���q��M?k��-�@Ju���]�@fm�d(�faI�(�-�Mk�b��	���uI%3�Vw g�2��(�����ش��~Æ;�b3�Ws����5�c�G�#�+Y��� �9�$ }B���.�u� d[bg�2|�+Wq0x@�|������	�����@���ǸIJ���+a� ���=�[�)"���mODF����ːeVc�X�׬�q�*����0�S�"�1dpC�J�8v�zQ8�j��5�����訖*w�co�5��+��#�Z� *��i���܆�-��}�7��˲������d�U!^�$�<��{Hd-�D�`�ݴ���~� �䝚b��i���������WKB3��%� �v�)���U�&��/诩'�I�4Vލ�/�9�kww~��8R,k�Qa[���A��9���6���cj�(���e�]QZ�M\f$_�j9��2���u��Z��4q
�	m��]���������V؝�����6
�3Y��3��!��<���#�v`N���و�ē�.vn�y�M�i��J��?ʳ�����-:js�;)S��ώ@4%f#��0���mT��<\cJ-Kn��@������1���	�]^ڛ�x$���}wvKJ��\�?	�j{�׭�S���������
-���o��:�b�lZ���Ɣ]jt����3܏{����Ry�f�5�!�J2���_�z`�n��LE�V��8�/���{�K������h�l?�<IlF��� 
��򽚨I��s��m�����"x{5zv�-N�'␃�QY0��b�gbcn�M�uH~ ���#��V% �;�	�e'N����A!Eg�ҶҫB�`����;��3�Sr��#�7S��,�(��=�����)�ٯ3��,˺�#�A:���_[���e�m��q�Yd4�bi�(�gjd�1��~�WL��*�;}R	1*�4�ۼ����]PC3;��>H5f+�M�2y�J�����X$�S9�9
��+W�\ϺG�	e\ )DX_-��_Em��yt�<���,�f��Nl��xms�r�y!g�G.�V��E0�|��o��f_W����R �Q4��p��Q$�2B���ěT����ޢ��"�QHF���_�G�b�RΠ�40gq��؉���CE�ٹ�T��\
S<�?,8�����ZB��$x��]�s]��k~B"�u���Y�G`U���W��̡"�Mx��*�9"X�+;��?�&d�2��O�aN��i4��.`ฃ��KKw�������*����t��U�l�� Xя�3�>^̮�>��c����I۸-y{i�Y�Ś�Y�L8�'��zy� �G�.����
�E?F>���T&�S�I�y�]%E�u��P�Ț�ň�b�-1���l��sG��h�Q�����L��pv�G�̬{o�UhhBd)��ݍ%9d��|'
�b�Dč����GWH�OՖ���7��*��J���s�q�[�	"'bϜ�b����xf3���C ��a���1i�
P�t)����L��Ng�.�vǨ$G^\�=?g�c&����� ˘�ъ�o����Dh� 2�V�\�9�.eY=��u�W�QaP�"+7�]KJ���s�lAȱm��]���8}�Ƽ���U6?�Kz��$��0����=~N�p�Xdk��| �CRA*��5U�2���y2 2�#~�?�]j���Z�z`NwHxP�,Σvr�Q�����8�;
/��y��y��m=Q�(p�H��H��R��t�(m��gy	�{�8���sp�{�
P���A�2�G��P)OU���b 	���[��4��l��q�(AT^��73��&j�8W����v�nY�q\�S@��+�h��v� ��/\�M����$V��6� ��;��b�}���WU���uK������S�APJ�--)�� W�[���8VƔj�shtt�D/݆����EqlC�0��]yJ�`>�joÑy��G�U�沉��
��**)�x�{3YS��T��<@� � �J�[��>wPiFBʉ쭹�6�b��A�ɘ�#
0J�\��b���
�����՗=Ӎ�z���r!"���I��̔2�v�Xy�dű>LtLqoMX&-��>�Kc��	���x�<��N��G�H2�G��#���c6J�A�RJ�I;1��^��74F�k5�D��K�Ñ9�։��	�ܚ�~���9$�?�L]�*e����l���	"��_��#��{��?����A(.6���x�vLl�D	|co����Lm���'Յu�M���[-+���"c@��/��N�*l�)��Es�BG�ؾ��S<�vk��U���|0d�����6c�ڴB���rb�$|"Q��iNA��gĄ��=S��*I�3�UQl�%���1��أ$uR�z�"���Y�$#�S���P�<���$F�j^KGG˕P4�|�o�D�h|+��y�T̶������a|�0+�(0���?gQ=����{V2�>�����d�h����R��9�`�j4�����[#�n�������#�Ǌ.�l'��#��BB�}�o�%LB���	l��~��W�Lr�=�a�?�0n<]��:~���j*s,�#�v�E6���4-7G���\��'f�$AF�GJ|k�Y�H�Ѳ��?<�%1Q:Ap�N+I�a8<�r�-m�4Y �����AU�$��:&m��s�&��Ⱥ�<C�~�hU�̧�B�r�Z|&1���V��\�)l�B}��յD�F3��f&߇�5rYY0���	m�L���L�c0F?%���&ǫ9����y�>b�&Rs��@��a�0�a��9G���(���<T_l�_�2�>0$���[3�.�Κ$�����>��7��8�<�7��%�=���5�̷x/WB2/?���h<	�BﴌB���m������}
����O`B���\�tޢ�Ok>E��J��m�!��&�yك���(�ᘲt;ruk�쒰-ӷ����y8���%C�	��z-�"l��m���1�Zt?�m؃�D��Stm����ڝ�-���w��jT��T!P_A��Y���������ƒ�X0|�Z�tm�[%��'��A��<��ĝBF2x<:D�l��[�y�Xd�JW���sY1�Q�����,��+�axcy �s.ۅ��� ?��\��������c��ŝ~4���L�UĪ��S�g{'=��[M���[�E��zkU$��ȸ<8YC��آ��B��"n\����2LK)�qS
9���{�'��j��GR��?9�c�%N�D��ت<�"��b~Ƨ*���;�2>(wb��e	b >
I��PN��l$?b(��d��B��uQ�{B�p�wV�������V�Vy�@���b�HO�H^FK<N�Ǐ�!���i��31�x����@�(��m9�o��,��
[0F���v=�f�`�F��`�6�XѺ�����3�h	1��R7��_rs��7S�X��]t�z��? �=��i0|Og�U��A}���';������5#[�8�ۙ8���[V�{�|D���H(�q���&�K����&�qQhCi|.���_���T�\GM�H����ߕvcQs����ȟ�<:Ҫ�N��I�����!��
�{�)j�˓R�i����r�n5vC���-�P64�k���^,k ��W�[R
��s��!����/�
s&.���{���I��5z(Hs���g�	Eօ���A������K�<+��_�gXt��:�m, )Do5�kb[�W�X�o��qҘRI��ي� �H�,��r�c�iI5A����*�p��x�h���a<�������I�,���ii�r?�z��� _q�Ri��/S�����m(NnBF�7o٥�����Y��FF(��'�W�Xu��>I1EJ�@�\WN��|2�wLy`�f�do:��잜p[y��5E�<͌���6�����#>��&����=��'��ĭ	���@���[��2�Aj��鳾7L@AwU�v+����G�A�J����-�rT�79�vc��V����ܲ�z��K�.���uW���GBq�- ������	�ρ\c��3\ڬm�<0-I�K�_����F���NF��?â5j ������ٻ�C����`�&���2ɽ/ϾD��|1����J~N�逅�
����5T5j��c���?ű��U+���w��c�Ga�9�0��ʇʿ�V���%�,�i1���;����=����LE�]ʚU���}C���(���EWT=��u?�mw���>)$A�dt��'u���qZ|�i{���8F>k�]E�+e`���F�{X�S�E�SG����6��V;�UH��j���dO4��*_��ZIT.��$H�@i	r/ӭ��{Y��aF�a��i|�����'yy��*Q����w�pi����"1�����|���x�](�Y!8�zcn]Bk��IYNub!�*��t�za(���`��4l�^���8�AEB�����騸��,P�m�t�d�~.�^���ن������Y�X*�G9���fU��JY#��r�SL),7�h
�1F����y�D�|u*)���L��88C��hp\��@+Jł��e]�,�l1�H4�Im܃�S�=2�Uh�/���`�-c��s�VDTq��I��d��v$���T0|5(�K�7S4Cj;�5�^q�W�0ы����_N�5�+�?H��hL4�ȱ�}p+Ѳ�;���J��������OKv.�̶1{mwB3z�H���,]��()�2����AD�����Za�d ��ӊ��058Y���s:	��}Q(���L�p��j#`^pJ�̓o6�ު�9$P! �<��t�2��-��n�;P��<x�NuL�l%.�9������BG)7�-�Ju���rb�:!L�*���P5Fm��b�h�+�0⼸�IFsU���nm����N�Ź��-��E�Ң��901Z&���J�l���)�m)F5�}�|�l3�	}[߅ Ӗ�ʏ�Y�/�lf+�s-�:��0.�h�GLi3�3�%��0�xB?.&T�H�+�ĕ&��v�W[�"���L��%ȋ-��!�jձ��(t=��5���nX`�К�� s/'� ���Yz�;^�OLOwr5�.p�&�E��[���t���a9�{�
�Q��O�폻��`�߄"��LJ�!��"�\�	����,�ʗ�>���`��)8�+6����=���R���\a���� ���!���p�|`͒fW$������]X)�$|��-��~i��ʪN������v�"s������A�)�&䰳p�V�gv��c{�G�R�����ʯ�b�rv�fk�C�>Q_.*�A_�O�DSEx������5w< Sc���"�6֟Ď��Af�0֛B�枼lM��t.x��;���hϗ�(�RRn�]�ͧ�x��L�G	C �O��AYt��:�s�7��N*�e@#�%p��3�V����#w�k�w�fc�ZL�U�܀�P��\���]�LÑ���k���\�1�;�Of�����zmؤ�����nx7��Q㞟cx؁��!�|%�!�v��/��^7n��烊�19�SHJ�M/��²<�PNm�V��}/�&9��������N����m
:�3'���Q�j)|4��<?_<R�菫��tR�����30��wvT�>���^�ĸN	
K�%QQ�-�@p��u�`,�
<@4I���ޅ��iƭn���c���
���`�*m/�	�p��W!��80�!uˁ¹8�7���\E�m��+��c�֭���]�M�*L�dSL��,O��0����#�������)	�"�&e����"����6����||��9��d�XT��9P12ɛ�eB���j�|�Q(�Sǲ!+�Q�,X�d&n�|@Fx�0�����%��8�$�rs+9彫�q��`�b�>��X�x(�O�(��1��?S3����q .x�мӵT>�����-���p{24�|����l��պ[����ӳX��xXV����O:OGhD�4,&��w�i���U����Q.e�)m��\��U/K?���eJWCG���Nyd�K� Ά��	���-��=�u�v唭��>Lg�aĄXKZl��c�H�I���
ÀH\I�P.!��n4�a��8^V_4�����nẬ�S~�a��d&��ϡ.�X���m�w����	��h��s��k��|��Wa4;�:R(dZ����dM�ge��|M*
J憘��z�\��S�QG��-�`�F`��#-��D���I��a��Ӹ��N�<���O0ӹ�������1-0P��y��ĎྰC�z���DݬZ̯"��Qa�^C�`}����4Z=����PG��'.��y��y��*8�"�L,Q
�vrH��åқm��b��,9^�`�Q���ZNW�MLB��]�Ӿ7��'"��R��!��
��Y�4�0w�
P2+R0W�|�Dr��
׫y�6C�4�D[,$�K��<ã.r��Tw��v��I�|PHZf���3���[�n���-p�����u7��XzC_1��罡]n�t���Y_��ً�E��)
サ���J_Eb4|oG� ]2S�xS�g}�z�������sg���_?(�,��Vd-IBl��	E9���N-H�Y[�
6��E�<�=���4���%��-��O4��{}DaE	}���{6ý�2J8<���rf�G�WǤ/q0̎�-��-f���5�+���@E.�������P:�mr�򂉾ɵ)6q�]�F�4�-A��lξr�F�)�գiÀ_S+'	�S���f�$�Dg�o�<��q�����B���%p��n��+��
V3=�M61�{8T�_j߆�7��,�HB\�r�C`щ=�&w�`��"TH%�>̋w��Y��8%)��G�VK���>%Va��f�X2���#��[̀���I�ƈ��Y0�R6:�*W��jt\�pqmf�E�g��#��}�0�^/�`���c��x�`��rrU�g �-#9�=Ga��}5�}Y·Ɯ)��ueQ8����C`�=̏�a;=0�"�0!�&g��k�!��[��+�^�b>Wb��u�Q`�ڤ�1��vR7X��ϔ�F�f�U���{����y���	���z}����o��Ws�31�O�!~��ףIA��ű����a�"K ^"p�~z��dJ�35��cʤ��te^*���-�jo8;�$���F�����G1��!I�����EK?��s:?q�ۍZ�uR���GW�[��ڞ�k�������/}���� &��]�s�ς�K�M�"�H�׍���_+,�tK���8c6a@��)(�yț �(�ϣ�ٔ�M�Ρxَ&� r�ň�)-�l�H|hN��+��8��a!�"�#��q�"xs�>1�4�x����Iir}Cȧ����:�����Y��x���+�r�e6�֢��,���C��X7�e�p��,)� oX�*�H�I�����Ѷ֞[�ݫ�`Ցh۴^Y����\���J5@@&�8����h���(��PRVqyt"�����`�.�����h�2�|�D$`'�W�6#٢s�0SI��;&�q�һ�T�Z|��hYp�zC*u�(��a9a\��	`B�3θ]��6��~j�;�f���J|(ϽD�I��|��;KY�9�>LD<�"&���eQ\m���ѕ�?������>����0K�q�v=y�K��c
���Ж��X �6'����mzZ�T?̯R (,#�=Ŝ^$s�=C����<&��b�ha��^��x��ܚ_S�o�1 ����������J�pɴ�9Tt�����ا��u�3gΛ&i��?�����=I����5����8�&�X�@�%���z�M���q��d�W ���XNX����m�^}�+H�C��:�T�	2r׾n7�zb��J���1r5�I͈AA�-(�+*/��L�	.���"E���)�1�ۊ+N��Z\9Z�.xln����>|�,���1?aq�*�l�|D����������V�e���֜\��7U�6��ÿ�e�`��?m��nUf=YG�Z��0.�#��q�
�6�Ҁ�xՌ)�x[O���6��j�H�2ĥ�<�,|���ҋB��7'��@��y�kdBё<#��Ƶ�q��B}�N����� Z��k��P�� �t�D�ДUVb��S#"��b���㑵o$��l�M��%�ǟ�J4�L%��=�Bs�����b /�L��O�6�+�&��@�X,	����w��}lk�N`�U����%��I[�|��� �7��A����l�"����%��\�[~��w�%jy��P�	����Wp����W5�D"� �������T���+֡�p!%����G���Vɖ�����*]�@�i�C&Q����˒�!�m�������vϚ)&��h�&�Ǟ