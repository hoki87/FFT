��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ����������h�j����]*u�ޚ����"v:\���r��XxKP�kٞ�G+�]|3]ڳ��b�?(�K|Nc���:Q�����(K�P�;|Q���PuZ�V��)mD��qd	�}�\��(�v4 �n��9L�l�"����}$p��Ȧ���=�_c	\ʻ�l�A`���wj`�H\D�j����-�c�4�����}�I�%������і�]��}�mvt{�m�Ke���$�j�q:9��jG2LzY���_��@/��?z��ޘ�����o�FOއ�尖 OwԜ�ơO��B�����C̀߁f.���2 $p��Vnz"�Dv� �!իዽ�a�h��F۬��ѐ;�=�$��"=wm�{�Tz3S�Y@6g�I����G�>��vZ��o�H�f1�t*�+猗�4i��-V<�-���L�қ9����u\|�
�&����t|BaA���!B��Ѡ��:��Cf���VK���{߲��x|��A�%`�H��j�K�^�d�=�F2�up|r��-s,���N�����t����,����@g��M�R������'��� �W�M �Z|8��bĮ�r�S�*�[��\ƃ?N��NOm$�T���x���d=/�������V���g�R]�z��y�=���q$�}�+b���Z��ZC4�����ދq�>�l��+E�����ߦ�0�z�P����2Q�SE�n�����"��O�+xS�� <ql˚�`��G�� �����M��g� ��.�ҽ��=�S�[���s��Ǝ�}$SA[�u��\����4���0iRa���}]��ȨG��ix���}���S'�Ż����)x�ʍ�3�������ʴ�V�=.�#ndI�a�@@����b�/Q}��-��HCU���&��O�vKPM�{)4eG�xH_��b�=	Ej��b����2�lf5o(!i��CA�Nw�� f6s�E�uf���z�G�R�,���VE~���ڶ������P?��C���/��j84�4`�
?;wF��AԶzNsM< ��|�UJ���y�㣳n魺W���Yn!5"x>�N�6�*�P]^Vl�^Rɀ�:����Or~���B�9bȋ=S�j��[r}=��u�D`JFʓR�s�{�R��5�`��9
 �I�`IHְc��ʤ��7<��˯�#�&���W�� �Ө�A~2����p���
�KN��iU���z�2v<���~7]�I���BYo�ײ���؉Z*��Q�ů5�� V4}��o�n|����ĥ�3�C7z�$agyt���0��8��C�蚮���C��:!���~#�hO޺v�H�Y���z�g����AWY�6��7V���/���@�A�_t7-]�,�ν�O8/��U�Ը�rg�C2A}Ma���t3�\�^�a"=��&u����P��b8�VMB�0S�Z(�?�P����[Wr��C\�S�z�Z�M���#<�O���Ȟ2�>�G�$*TLp�zZ��N�ѳi�{�si��^�JU'������W_oU�A.N��ń{F��, �Hw�
�l�v�]��҉��.M�}�ǽ���mj�3A�Y��A�y�%��m�����q�פ��ٺ��Ȓ�j ����e!�c��x�p�h�Y�����GH!sZ3��U9=
��Dv�"�K|Q\�w��ˆ͹kl�;6!p+m�$���m�8Ci*-'yaӹ8֓���<2Q ������M���tI���ԏ*T�i����{U���둖��1Η��҂E�Y�2��PR�N���X�>a����W'�3.��:����6^q��m��='�d�N5����L�6x�pTM��C\?��Z�=1�?�I�.j�L�>��S~b
��x�|��ۋ�v2|���'l���@����n�Si%B�Ď���@�a��K<W(�Ix��^A`|EɁ*�D�b��&0�^\Xj;A�]]�+�w�����r�.����G������$��(��b����Gq��	}��1��"���?������T�W>;L?��1���C���%'KV�l�Yt:n
7��E�h�PЧ,���ĭx�-��藭5?�w�\"_�q*9�����E-�;��@, f�}�0hJ�����&e�./�o�X��y�r�9�ȷ�]�8���*�w��8��Rd9�m2(���$��!D|u6�r�\B*$Az�jt ��O�Kl��e�,JWb�o	)+f�)t@b����<�6V�Or˛���+�*����	s�hŮ���o��,�x�t�یz�}R�@��"�u�e���,��|מ�q)�h�?���.����Q�w�O���燺0�K��"N�l�	�,�����?�BO�)}�5}ȕٲÎ�cJ����Ɖ���"g9��m�R�8������D��u�=�'��2�^�B�?݈y�僡����"ޤ�W�\���� �[� M�r�=�,�;�/y��4�a�B�Gס-�����>�\�bw�Go?�鞍1�M5^Zj��[��C�e~B�K@����Ty�V��WM-_��D<�3d\��5T�>E�B��E�"f���_$�o�q�������Ld����$�n\��Ná^IC)<��"FNv_u c�b�wa:N�-P��'�q&�����m��@�)��li9~�=�>؍`�T�K+�Ғ|	�L=�W[�<TN\��Iw_�|%w�%8�a�0�2fZ� �e~	�0�gl*%�L��C�ـ���#�nλ�O'��!�+�G�2� �{�F������p܀,��+���߁�yN����"��ΰm,�����yp�v���b&l���D�i%obrZ�s��J��q���!�#m�o\��L��LOH�;x�U8��Vp]n�c�����%1�~����(����-��y�b�0��Z0q�-�4�o�X�^�r���c��V���`KhV@�Ʌ!S��2���R΂�	�����I�|�w���H8Ej�FK���ד�Hsw^+����v�?1W�����V̾��ö@!?4čF��p�0/e�����R��e�b��`l��Z=[΀�MI��o`�	}w��������!��~|ȓFe�0W���-O�>��2�C�Ky-��+"I[Cɵ���0��L�4��DNr�����LsO*	��	9@��c<�?l�A`,��p��%!wȲ�MCҦ]�_��K��¬�6�zo��TO�ؕ	�H�%���]b��`�J@��1��[A�<�!J{3����˓؏0$��N�?��J�6���0y�Ni�0s�+���[���釭�T�6�4�ɟT�rK�9zr�R��{��a|�3G̴a�S��o�>k6�[ZČ��~�*�b�aI�k����a�cH�?���;
��̏e^�� H���KU@�H��V؇��ʿM5��D�k�E_�������z����h�DS��4���n��$����L�pI��@>�Kg}������ֳ�����b��h��&~�f>���e�z�P��F�}�+Tra`G"k�ڀz�A�|fnu㍅QI`(}+d ԂI�����O{
'����r�HZ\��Z�4-7��y��@Ei٣�r1�z(����%O-�����S�����B#�D��Z!�rV�����.��pY���o�Xv7�dV��?�6hYFc�^p�Pa�46��r>[w1J
c]V�lO�}Tfϫ�^�E�[�W����F7x�����\��z�@OL)"�d�v�F(��/�`�7�E� ����1&�a��pڮ81�K�\BޜCv�M��{����_^���=fZ��zh�f�j��M`$H�G�;�MiTo��"kdqQ��Ց�bb���+�JB�2�b!
bI��Ws4f������X嬵�>yC�$�z�mHy�� V�U��_>�i��oղ�c�S
*B�^�dR!ݡ��4��s�ٝ�Yn'�M;ȿn΅7����_ؓ}<��M��wJ��`�y����	���D�)����9'�!P���Gi��bi���� �t�����e>z��l����iA�뾘N��r6�G7Z��KC1'W��^��q�W���fÖ�&;�cAL��n�`�)�'����fA���M`*��4����-9����4x���ջ^��X�F�=����[�}А��폌_Yp��LU�O/��z5�S�A��/A~�w���~fd��� ��c��S�%VWK�tX�M�~�w������Sӻ1�Vk�Tt��k-	^ J}� W-�������tQ�o�kO(S����bus�Rw����D_�tB0� �lM��:�V�@�¸�d�{����l���4��RO޽�����#B���H���x�P�
%.��p�p� 
J�W*x�Y�.���x�ɴ��¡9�a��8@+#����ґB#� �e�<�~A��K�2�h,5 ��;�b���e�
w����_+�8��|ey��}�W`;B��C�}u�41�{�<{��@_���LM��߿��$Z�}�w�[P�H�=�����/)���$�E�z��(�`���=�X10U#&���J|fQ�_��H)y��u�{@�Z�5�B�Dp��jTMH.X�9\���$�"<�j� �|.����y���Z`b��%t3)S�(k�N�����괋j� �$�yR$J���~@2�&�������a��_���΃��AW�A��r'��}� �EQ���J7+Tu��F�xD/��� �O���>��@v���� ��G)��@������t�K��8pY�4؜3ʾh:��״�	錿;M�	��S������#�:�����M�(� �M�+�"~�|	b?iZ�rl��U��N�6���R�fQ��	����R�?S^>L4��:u ���,�Hƴ����q����_������B�8i×2S��*�tie#��!��d+����OY�pA���7�V�Ϳ�al�#+)g{��4��nP��)c�*n�&�MM��ن����R
&G�oZ�Ke��TD϶�Ʒ�;='���p�<����2/n�NqlZ����'Vx�X��TS�G&�*2���˟�����;�Y)�>� lTq��:�A5����v�e�x��:Kք�,F�$�s��L,Y:��:��z��|���ZZς<�!�6������"���BRa�z��_<��X~�(YP{�b���j��灖A53��PhL�������7��7i��c��0����c��\*���㿜�)�uL�2�::�z#��8w8|��Bo3�#
+���f�c�p�/I8����v͐�5{{%����AofA��w�眲��1��`<ly2�����.��x-`ZbD���oY/jQ?�[LGP��e�N�~�C��oLߵ��������! X�������۝���h�HoC�Q����|�W��A�H����m�%@��>l���J�0K<
�WX@z���:�
�/˝�CZ��*M��ea, ��F4+זa�	��1�F�y�J���B�+m��TY�kY���ޡ����.{�40��Fvl�?=�j��Q�o���3�ϗ�P�͐?2�Y���J|Տ����D�����<�~F���`q�^�l0��`����1E�A�L�2G$t9��~&"�ގ �ʏ�*pk=؈s�T>ɪm��Qa#R��������%D���ȃy��M��T��+(�h�,�od�uΣ㎔�"C n��bv��As��Ѝ�����L�.҇&������V����p�R8.kN�LoFRj=���"��v������ �1��A�n�u��}Z�⪝P��Ӊz�/i�����;қm��1����k��
��`�a�r��nL6 �#E�y��WQ�	��ζ��.WY �A�&��@
����V���(jk���Г�w�,ʗ%''Kڠ�S&.;��%'?B!į�� &�r��]M��]2��'qM��_+T]��
Nk����ا���m���_.�,I�s��[S �9_�o>:.S���A���<�W��MI��p�N��8�1(59���(�n!9X?s�&�W������C�̩a��+1:n,��y	A)!%���L�����&w���ȱF�7b-	��kBz����x�.����Q�,S�� ]JCul];<�.�V���2`�D�g�Rk�+D�K���8�M����Cj� ����.��b��j�\�����k�뒡#���r������\��NQ��%�i7�Y@­o�u�[���R���5٧������k� #�O��)H�f�����\�Ƕ
ZSr�@X�:cNF	W��"�*h;�c&9����Н��%�*��H�����}�H�F6\"��j*�������,�=:Gc�"K�_(�u���~��.�m�ِ�n}�i��7�h��(�VG繪��ύ��| �d�*�1��u�Z�9�w(]�ݬ�4�ʳ�̪i�SZ�6-{�ĥ����j��?`�e�us����Nz�t�7���4�Z�G���, ��$,�Ou;��n���B�9i	�)C�qW5�6M�[1d�P�)~��(��i������}K0#ږ�_ �w� O�5f��y�Ͼ	��ڞԫoJ��F�,R6�ѾC�֚���Z���8��}�Ķ�2N�ɧ�3�M��f�eQ̸4��'�L��;H~��k4dSz1���As���D��4+�M��9�