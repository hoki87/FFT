��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ���������B�N�-��)����!���NZ����p$`�m
1�&��8��C)l��?�{[�������2|��ݽ�]�#[v_4�!r��Q��/��%K�2�[\qu��j��ǣ�uP]PT���
�둽�i*�n����p�xЌ�Ǣ���9|E<�oD|_��9jlbD�~(� �,�!|��q�_�#���f.��}��nIW��|�Vy������*����s��W�r��nB���'�}_��9�����"�R�f��
��]�v����9�+���+��3���s����~]r��u��դ��ذ2>%�G���Ŵ;zV���uE��qt	���v��ۥǗԗ���⮢���QΙ�\�?�9gv�=���$˭-��i��A4�[��'�
WX�(%��j��	�4�wӨ�������%!��@�wW�KP�N���8�UUs�4N��3���f��XD���<��ٗ���O�	��+��>nڣ߾P�6O�{�0�� <��&%�uM�[h�&�crYd�K� B�F]�_�M�:�>�g����bR�I�(=p��9N~.;l�u�\E�����9��C[-��^��vʬc�S'Z��<��[�)`�g�YU�@O��+�H����ZQH�ĸ �T^����a������K]U�"���*S����b������G8�M�t��@�=ÿ��`t:�ݢ2�h[��čsň��M��r$���|UC+_u���Q������H]1���L\�s����9�N��h�S�"��s�w>������f��G�ėc ��0̟�G��]:��RQ=]à�����~P�>1 *^��t��x�.�4E	�9Z����?˟��j,��s��
A�s<�	� ��|�S19�e�_�f��W���ԩ"�+�x�5����*GJ��}R�q�Itu@�9�����U臰�Ȓ�"$�9卜� e��/�d�6����`�,euP�.�Ȇ�e�x�`m([��I� ���֞���#��V��4)�*�G&�F��纍���(x�u�]��0YY��^��k��hp�������@3Mg�y���7��������j�f���|W�ʩ�0^7���2_Π��j-4@�a���~r�4�*�u�0���e�-z��pjַ�������4Z�*������#<T]��xX�D(ٰ)�>�F,b��G������t����������afK	���#�@Ȟ�����[#nZ���O�X�iۦF���y�`�N�V�-��]frT ���gR����n.�L#���<��2��2�}����Z��gK
9��	�t��%�$d�] �1e�����X�������y�I��Fxc�j�KH!��j���[D��S�l&*a6ɧ�/U���/n��FW);� v����	�H�� ��8�Iz�(Q�GN��/h��םOQ\��	L�V;�}]�Z��ؐX�߅��"��x�2<r��Mɚa퓄u�|�6��'��*�JZ���;zտ韦�;J�(�)�Eq�C�����U�K�$��Յ����PI":�R׺d�/�}�U��[�T��x��NߞV#�#��-aS��%؄@�m�˽�h$z�
+��r�% �w������h�mګˊ�S�\��q�J=�݋�����'h������l��u����$�
�*������V�d�q[;�'@:�SBlȞ�pc�\���z0�߭]8���'��!�'Tuc���x�;0�eKk*�����S�<y'oɶ^���|K����J3�AC{�srK���߫��]��S9��W~�y�
��6 ބW�hZЅ�4�<_WƮ@�t�|$G
]W���I�g*F����K����]�xvlݎ���t x�m�)�T<��ML1#��4�A�]z�q�ǴG�0�U�������6Zln���JKj���hګ�աNb�?��K�|	(�w*8�V/����2M�<���vڵS�`��V���8ʷ.M�(@d�M����$���B�גZ��,o����m�*N�K�)u��˴��W��߳&hhet�h��`ځN�
��EAЏ��Q2Fx�
BEg�~�HP��1��a�x�����\�KpO���nC�T�һ�rx�Ǆ7'��"��6��S!��Ƕ�<�hU��B k�ܑq+p�c�v��T4x0�0�$�� %��r�Ͳ���*�_q%/Z$���5�v�:7(���!;]���|)�?�_#"�h�й<��w~�o��V!�$/
Z�J|������S8��</CI�+�78�᭑�=�f\.�Z��~B$�wi#���+""*�A6s�y��2��M�����؏T��ߞJ�(�[q��#�e�͛>��ӹ����S(���0�T�-�M �4���������ۗhp�m�+?��r�r�*q_�����~�A�hZM�x�?���Ф�w�^I�M�?:�;	�<F�ń �Q�}�_g�T�����i&�n�����~��ۍ��91T�3<�R��Au]������ł��ݦ�˖�￤�;�c����b���V���;8]�:��Y�i�]{�e9��P�vK�	?��%�d�ݾ/�jŜH��]��앇2Y�F@W�
�gDcWE�� �6b�F������A�ޚ�Ǘk ��/�����y�2=��;����Ȗ> %�W�g5�P���ơ��:����qF��|µI&3�#��� "i�U�?-��'cs�,��C���5I�F�W3'���wW�և�XZ$�Z1�;��3������xWl4�[�=k��䣞ϯ��ͨo��L�>,[T����, h�#H���рY��k�����˙=0���b�U��˧�m*K+@�*O�@��$0�Ֆw�����Sbc0��r�5�b�NP���$
�uZiο� O�%{�	��,ӠgTP�/=�{�P#���0>����C_�CV�)k�W�j~���5�1��U��TA=�j�"�6��g�2 ���=v�r�����V��j���B)���6Vb�vQ��ѱ�9�b���,S~'�V\ȼ��+���2Ǫ�Q��SL!���3�)������
��g��d>y�`"L���M	K��`,e�ߗ���8����snuMJ�[5]�џ<*|]6�0���5���7kKX� Jl4cΧB��"n�#�����U�N��5ѵ*뗸!8��D�D����F�b�	�W<bSťԾoZ�7�sWፂ6�䨓���&��E)�dX�k̹4��#�@O�I-2�d�S
��
���0J_��I��F�n���)����^4�IKȾ󮗢�dr����ڨ�x��m�3���C�̈⃼j���8p3?��w������8\��X��(tRۘ@x�hi���2��b>$���h0�x�g�zb��xz&v�	�*�f\N	1< ���p�`��"���Ǵ.����kG���+nr��3c8-�5���Pϥ��$���:1C�%�È��t�Rj���GE��f���o�������,��H5��υǗ�}���Ee���:z�[��3��n2��P L�Sr�[̣�"���T�-gS�e����p6�=�RB��D1�uy�{�R��)�_�G�a>����6�N��n��
���^g�i���TB�6x�+��P��]���m��b.�$T�nP��3������u�����398�4Q�+bfB���n�l8�`@���������tx�l�$o��-ّ_Mx1�!H3���L�]���Y�3(���a�EU����G��Wi��P�
�x��N,B����hP�H��9�*��#�!ed��N�#�"к�)�Tᠤm�;X�>~�znqӲ_A=�^�*����"��9g���}���o�iiY���[�;t��hS64x�K+���[�� �&�t��Y��`�v�u�n�L���-��@[1��&�:H�r�-@�x���������I[���0�q���Ĉ�]m�^��>4�x�o8F,�gi��ٓn�N3<QZ���iB焕l}��Fu�ˮ�Z�($#.Ibhќr������z�-��3o�!�X���{��9�,'�L�����g��۠	oN�q����D�����C,S��r)��^�1�J:´��+���vgҋ���t�NBA�o!�S�� _�ֆ���|xrW+P�������<��sP>3�� ��j(j� �U;B��2�N�R�q!����C,��}X*��N0O�Y�~���.|^"c��	�i����n���ç6/�� �݈�Z/�y���`�"���tfW�a��㗴�G�Q��=+w�%XM��i������(��B�o �z?万YW�68Ag�����*�v҈�mW�۷��=�]��mGi�����ŋ��l,N^�͌^�X��>�+�a5�A ����ǳ���<��#��2��/S��y�ޠ�L �\�
�Xal`���`U뻉!�c_��SQ���ӭL�r�/�Zb�-e��,�]mA�#��5`�6���oh�Bx�)n���ʮ��94��D���-����I��ˁ&�I�IA�=�5�>��������؍��N<�eڶ7��k�A�+8�ż�O����*��H�:���B��!H���u��-v�'\���$�-���*�G��vc��T��Pp���oUȹ�?{"X^@��@� ��i
�0�F����xh��T_!���-�ڤ�d��e���K�J�Q��U�,���-	S�5��槼b֪���kb/M�����.1������n�3>RO}P��~H4��=���?kR�!���v����ED���KA*
�F&����$������lXA?�5�|�f�u�zL��p5�K�$�C	���Zt>ϣ�0��ػ�碠<�!�l�wUď�5�mT2�\���^srO�(�8���:@W��Y@��ѻ��~f��`���JH��i�pݒ~��Y��i��UZ�#؇ �oz�����`Ȳ��E�?���=�����Tk�
wϧ��aN�������p)�����J��0�|�ޭ/F����5Qe��4���c+�d��˜��;��u	I,k�4#��7�ש�L��j�;S�_��<ݨ�7Ja9g�<��¬�i�'�^��� 0��QM�IpJ]A�lAqL	Ҭ�T=����)7��Ř~��#1����	�vfZ��F���X/F1hP�2�%�5�d��ࣹ,(	���S@w�;���o4	Q�9�C1@PP�|����,�*���k�~C�� �M��x}`dΟd2UW�j���� !T'����kJ�g�%X�\8��u�X�M)�Y�%�F@��Ε"á�LF�p���	ä�����M ���	p�H�r/�����z�e}�s��}4����́*���D���Oi�h��"���0���e�Kl�P����/����u(�Y�Fj6=�V�fw�,,�+3���� յ�>��q�N=Y֓���9���_a,9�|./[7��7LTT@Z�8���A�6�܁��:�����f�댷�7a�sh�Vl_����#�Z���kfky���(��k�"�e���#4�*>�z�58i��u�I�~^�0�wtZ
.r�s$�+c�0;�:'�w�^sF�ᚨ��_&S�
��*䷩_׋��ƖS����=�#���YΛ!d�����Ǔ�����H��9���?����|��U���m]�]� �5jl��K�-&�5=,2=h����6y���QplC��3k�M�x��#X?J�u=^q�6��6M�j�g���'b�>�)��
�*���U+:�s�xO�������a;)�r�/c;@����q	Ã�o[3�J}�L�֣���B���c����6��Z�/	�eX7���g1Ww���ku����`ڰxP���A&$L����H��lV�j�r�0������6�� 2�S�����ve�J�Z�>���@�G[黌J�Q(y�r'_�_�+��`g��^�@����2A��6��&�fם|P9�� �(D3!�+B���g^�D���L:̒@�'�75:�|�S&��hy�`8e˒��C�3`�ʭ\q`/<�%H�r���zܦ,���|�}&���8nҴ0pp 
["X�Ү�j%r�E
��9�661����3��N���น�l� ��xT�z{��N
�%����X�Ƌw"���ë�"���ʩ~Y���p�S�
w�"��.X�E<�������`�M�~�.�c�s�����O����%ye�A�%���v���V+E�"��Юl�X�(�R�β�v�2�8�oʹ�n̔$�TS��;��ʓ5��yv�`�-�6R�ڑ�ɹ?��{�[�>$_�~%� ���j�SO�6�s��������S��~z��2xM`���.�� ���2�H��A���]��e؅:A�x�������`77Ď� ����Bлz!p�b�d���W�l _��tn0���3a��l����p�+8�x"2�{d��� ���mVZ�_��*�'G�'ݖ�T�lŲ���h�+�M�\N��1�*�W�~�*#���;W�����Dq��o������c����'[�A�z�t�*͛�U-�r\���K���e'NҰ!Ȩܧ��U�Qx
�RB��e�_��EK����&P�GP۽~�e
gAkE�O&��De��t�5+[�߳�??��y�W�;�nYCJ�E��� qW�K��90-�`��O�Cָ|$L0 �GJ�"��XS���Y�s�&����U�d�jmMA��|�����!�X��\d�s6i-�Fn���T����v4�}�w(����I�S���dp}���g�ܖ��V��w�#c��⦒�ǌ��YU��t���n��2�g�hl��Ņ��,�9��S��H^�e	!ɧ�����U�g� &>=�O�� ���R�.���iFO������L�L]ޣ�/{k=�A��w�B�ӳ#<����y<��FCef�����|��O����siF?p��CnܫV�jL������@�����d�h�[����|&G�?30Y�O2��.��1)#�/��n��S9�]���/��Ɔ	L�J�4��'����C�h����!(�˃���hT�O��S M��HU���Q�Dq��$� �0�."��U:���w�nt\�qZ�vz�@��a"F�2�90��w����X�xY�� n�WW����,kP˜��)���v�t�np.�:W� B���.#c�k���Q�X�_��l��}��Xj�D�4H=�Ꮳ��G:�#�s̤��I�G6PR�P~B�2�Y��Ż4�ܴK�!IޡF���e5Kz��6��(���y/�j���L$m��Ѡ���G�ؕpҙې�Mxޒ�9!�4�WP�_��J����ڪ֌eO',.�\��9,��4/%+�W!�B�ڜ(	fǩ�׸\�0��F�1I�LD�̏����V'ƒ���}-|bAPe��Nv@���x�C"����+�T��n:����Aʫ�ح
���Y�i���X^��4�+ܣ7!U�(�sU}T���w�uRx��#�\�ǩ#Or`����J;ajX^{/%��`Tn'�r$ݦ&�@[1�KƤL��c�$x�ʫ=�+L�MfW�R"%����6:r*��>�o}�y]��_u�o���Z8�㪁��[ɒ��q^��7Q���b���n%#a�
����k��g�	ծ}��)4�'��^?c�L���]l!\�4?�;&jU��u!���*?�OQ���9�ܚ�5��$�{rƠO��L��D,�r|P
Zvc�ts{#��%�_n�^�v��3�:KT��0g�ME��[����Fw�K���>�S��z�� 6dB���"p��F1�G�/Z�_*r�X:�%9����}���AzޛX�:�'Ǖ��>�h�tP��:�E=���4�UT�:�[��#]��c�li!��-%�xb-�ZE��0,�	b>{�'f�R��~Z�J�[5.�*���6��-U�9�O�����_��j'���_��A�+�nǍ�9�Rz|���~2��4Ff�vY��\r��ǗC�����%�#�D%�#�Z����'�G(��(��Ow���B��J�����]L ��ob�(p�����n����^TTR�ZR���/����
u� ��2��Y��OC��l��h�nE3b�� ���T�h��
Z���u�5�L)X1�b�n=fnk�C;q�(6�G2@�[�(�a�K�ʉU��\y�\�G]glʙ�k_��.��/tZ�z~��N���*c�վ����\G�5�l3�5������*>�؍�1ds>)V0�^��	�L�o����|?�"��܁���[AY�ُ��E�-jɡ�F̄�Q [G��\�'��w��7��G��l�H_��Z�% ���yz�7��R���n�;#��n�ӃVg'��
ٴɸG:�\_[f��?�zǜ1�Lk?p�>�/1=���f"媜)UT[��Q�k�͏Pb*��t�&�f��&olv2�%�w�X�����+�W��.��'l�|X�S.>�@y���-�-_����˳��y9Q`�|�*aqTg�W�<t��
0�n��_�zCC�0X�Xl"�[�#>G
�>���+�Ր�m|6/Y�X��s��[� �Y�r�jb������⼿��l���+�H$d�*��~�D��f�jy�0��'���3���13j��əj�������{�cG�dt����N�ST����F�C��b�$6�~�!&V����4�M�'T؋������O��XPT\�^��?P������j�7 ������������8{L&��wX���s(h�HZ���$�T�?(���Y�}��dd�$;@�7��ٷ4�0�Š�����s�_zs����iG'�T�p��$^�s{�<��/^}����o�m^�c#��C�k�q\�Lb������
<��{ӝ�y/�C�i��8�S%�.S��:�-�|��f$Q�H�O��$�m�kK����q�O9ގ�um�w�h4��M��Dpl��2ɇ�/�wd�*[��G(s�)�L�'��Ǎ?�W?$��*�l�k��^�jb�����7��+����=�F��:��ޅ��`Z��|\�BO�[�\`�H�/$I
��\��"������Rm7��E� IR��A�v!�6���꭪��\�-Z��	l�i�N{��y�^��l�������N�摫>���r�9_�x��Ľ�G����r�O'd����&�)�9�P"���r�d�(�����k�$v�G!	��i���(����;f?7��_{�2���X�|*w�јN�P�j�����7}��i�M��/ko�̑�V���/��Y�.��ڽԭ�����Kf��'�kj&�8���2�j�8�?�?�a�D�R��9<�͵�WXi��P *o��3O�,C
XB��u2�9+�L��o�:/�0������vM��[z+��c��sH�#����T�hI��r���=�9����晜e��9����8�9R��|�"N�{�����uY^|����.��E}MC𢑄�y3�B�z�;G�'�tL=�0���P�a��n�-рn��w��dJZ0ݺ������m���R�넲����'�hnќ����l0��P
/���
9�L(�>�P3MD1�@��M�G�G{RQ|��^�����7g���'�p.nށ���0i�]�y�`U銿%Pi��t=I0�����w^�v)�� ���"Wk���_m'�2�"&�� 7��f�Mܺ��L�MT����&�;X����;, ���.1�����p�EQ����"�hV�K��}��\��4ǈ쵓��+��E�{�أ�o;�<,��>�s��B��������Hs?��EN��E\��˳�DO�TS�����`���2�Z�W���"Ɖ��s,>�.����ڍ�H�ߖK� P��L<퐅�����N����(7�ʑ|23��'uY��� s����oww$d�J<���Cg�G~����O��C
"N+�u�8z����ٵ��uۻP$�Us�`kF��BB�v?&O�H!i��:A�]m&�j%�Ae�,�`�� ��߫8��^��\Eh�3H���(��}no-�ʮ���աWK�|ji���H
xb	4��h�	#ZLw�|3�Q����\�+���� �������<u/|$�9�a����z�m�7o+)��zpрh����֣D_@��5�DCliU��U[�[��(��|�b�u�qH��H��q���c��`��!\/a��\()
��qm�~��`�18atqz�8\� S��&b�Բ�ՂX�*�z�lI����<�{�,0O`8�>�m�X�<e�j7�k�}e/�Lje��u��2=G=�/��*�; ���~9��H#��ɽ%���-�&��Jslk�Z�[�S�*�0+cZ:ٿ#Db:L��BO=��A����R۱����|%�W9��jS�P<��l���s�E�0"�!����8�a�V�w[�99�  ��b�R�[�CG"m�w�Z�1��0�BƸ���1.��̰�+�u����)�p#[��>�B���s���ݧ�*չF�0kZ ?Z�A�צqs]����{d	g��G�z;�
*��O�#%�����Nho���8f:��6@�I���:c�B���z�'�� o�I��Ǝ��7Ô>��D����A�r袎ކj�j�u�|�kYD#T�,���j�N��A=}%���)1��g��B�Tת�����U�� ѫ��%٤�n0�I��c�O揓�aU�����O:���3d*�Q0�`Ŵ���ɳ�~����Km�.�C�9�K}���Z`k�y�}>JZ���:��	�6[܊��Q�nmh��z3&R��v��*+�9���F.�CJ6ueAX]�3�ZU��nr5:�<"�6�}�JG�v�
��	o[h�����LM�?,s
|�p�;Y�T<����e����쒚	�ed��1s�+i��@�X1��<ʚ.8��B�d��$x����ü��x6N ��qފ�/MV(����H�H����R_CL;k%T�F>��}�`9�H^˶s�ȝ���4`�q)H��gw�f4i�^SiU!Y���l��Y�9���J'�j3(ne�`MS��}(?C�9�"=�1w7,A2��?���an�Mg��㶙 z�i�o��L��o-&�B���?�G�
���$ԭ@#pyjP��b7���ܦP�4l�44o2i�VV�}3)���
��}8�H�0�fVhI�j��t>���Q�AB��Q��l��Ձ��,H��6�"�~W��P��w�%&ە�Q�O����ճ0����ʧ���y96Y�^7����Ck�c�:�ᝦ6~ȂI�p.�P? �:��t.Ngl3����z��͍� �1��O~7��]�[����"ڬ=G�=>��wq������pFgc�s�nz?�ru���xݮ�`7R�Xq�,]��W�0�cy��l��H,�q�d	�����#b�ޅ��5�Y;yL!�n?x���W_�e�*��K�N4�8����E3�V~��X���E�'�j+�Qx��pM��ޏ����� -3� �Jz�2�7��9I�����U�w���,mx�w���/��wS�*�}Ē"���W�~��n��'��.�S�m���5��R�n@�>�ܒA"�]�"<��!�C�"��y�4q��䄄�b_��j�D�_��w_V��9�=�?n�����5��臌�X¡���/�����U�z�AaL���.Q�������L0��}E_�5��a���Uڟ���<'h�_��%��e�N����W?!��sbz��8t��N,��l옮�chY��p���g��6Φ |��\qu����F Gx\B���O�r��ߕ��L�H���L�_�������[�Јr͛�m|��7�k<ܽ���e\&�*xH�tx�l*��f
( 'C ��Skٵ	a��$P~��v#�D1=C>[�$�b,�����y��u*��VN��!�;��0��g��L�b���~�r��.%���a���7�u�����O�V�����o���W�������������*�(r��G��
}����xY5Iy�
��p{�x�,�%����3g�㧈N9�UMwf�+44����v���?:�m�����7������8ӈ�/���IC[o�V1�������[�aΏHGQ�,��j̞�&�5.�'�N(OyL���8H@&�_��:j��If��ԙ� a�����:�P��g�O�O�����1�`kۂY��J`7d��.����A���-�7˜�H��p}���N g
CSn�\a�m/RH��!��OCj���ys����n�Zd&o8�0�!)NR�DW	�o�ɬ��,�ô�0tD�ie*{�R(�u?rP,��|��|(c���F
���@����T����u�)2.�����^2N�N�%x��!z������=9���x@<7�@��(Fg&�E�A��u�4�>E3 �j&�妼|�}��銰q8n��Ӫ���%.D%ѳ����b���T��._�������=���A�͡f�]'�tI��\@;��p��̧7��$nqˈ>kI�L��j����.u�݃�b��i��v�K%�����
��"����/!pA�����?�;��!����z��w��(eb���Z��0Gw�H�Y�&W�9]�!m�WazTޏ�[J�h���o-T��X{Ҁơ�b�p��@�)��(ϖ9h$d/�(0Ha�j�\�d1d6�	�����h����$���^�s��Y�U;��u�t�c�w��	C����%!�����9ݴ���BW=ɯQ���a��x����+o|ν��~�.�����q�j��k=�Sch�9{�$�BIKp|�a�93�盖k�$��w>�Wj�G�<m���}b]�c�`�Zl��GLV�V\������	{�o��[[�s�qsf�������A��tΑ/�`2K]�O��G2���EtWҀ\Lf�i`_�\� �"��w^�����$ӟ�t�o�3,��i�9{0��-�6�#�&�Zb����sa����9������(����	���a7E�ІrX�U��\.D!��͇D�>�J�	a(�@vϏ�C�U��/("�g��4P4z��q�]v���/Bo���4 ��=�� y_���kčăpZ��GC�~?��D��^��(�	��t8�F�|��&Тp8�� ݟ5;_!8D��wvK6�Uh�����<Լ-�C���6"p'㫒��?���)G|��o�a�r�L����u�c�5�@���uT��?�Voh�t�ɉ����v�r
�/6���T�Y��T�j�P�9��eǰh)*�{��jH�Y�ps�$�n<b-> 6"��J�G����I3J*���`���o��hĊJ�#�d��$F�����+���,�}f�/I�us�T�nQ�0�A��.ղ_"FR�:M>�AD�yY��P��uX%0��[F�ۍ��SZ���Dx���B'�^�1��������L[��a�@!��ڼ�W�+�~���G���)��-��f��Pb�Z�_쩅a�V��iX,ħ�(��S������aL��^��${�\�Mlz�P�D��
�D����Mv�a�Yk,�D�Q�C��	0�B�O�dh���(TlKT�Y&~)��Q�Cl�9�C:�	2��Z�,�z�}��	�n.׉�H�����uD�+�n�߾������ f:Ew
]Q] l����fV!W}�a<4��)sq�U/S���yD����{y�v]�S��Qi!O��$�x;�K�y�TBfG�k3���M�Wk�ܑ�	�|��rr�lT�9YQȠ�w/��v��k����gI1�W��x���Ȕ^�����@�GH��`S\������`������	�2�����K�۴�(˞Q��S��-Rxe�Q��t&L����4#h*"�-�w`a��7�q��=:��Е���ШSēpqq������b�p�$�(�f��{D���f5�
� �ի�Z����k��#��r{����@ә��B�4}W�f�ή�9��+��3L��"RO�y� ez(���� k�=�<�����܈L�b:�N�d;p͉۩(Gx��ɾ+~X�00J���H���*��'����<���5>!�ju"n��^�a��i��8e&L/{Ӿz�;o��*P����0�\�s��C��ޯ�qŘaA�н�u��&��UF�E����[�)4v�� �*��I����.�mG�ŭ��	�*��ELj˕�𵈒�(2^��6��[p51�FMζ���sg|������J�5���6��m��;�za��%3�2&���J-v�p� {��̣�5������P��@�f�"�ej��$�~p��l�HV�G�`�lV���:�_���Yk}y�_u���`H)� '!�ܸS�$u��8;��(4�v�w���#�*��璪�ߕ�P�8: �&�&A<(b��=;���&�`5���_��ء�):��l~*fmY�S'���2�+)��@4P�UOD$rC����-�>��`7�*_0�(�����b³�u99�.��R�)�~1�n�2o���iL�c7��:z��o��l��Dw�$V���E�T�ֲʊ�C7�M��~� N�'rq���m�	�����3lS�m�|��KO�����]�.=��t�B�xݗ����e٪Ew�-2��]�`c�6�(�/V�7�u�-cWۢD��)m�_9�}'zo;�B����%k���X��"[|�c��/�]��N�Wp1ϒ��"���\R���s\2Q�'�'����UdR�D��ǂ��e6e�%K�[����b�~��B�����1[�#�+��S�)��,�o)�b�o�c�W7�*}>x#BZ��\�Vr��ں=2�0kk_<��rF�V;�;Z��~��|%��
���P���kN���絭0L��ݓ$��N�Bd3cǛM�����3.������+n�哻���n����i���x�z�W�+�ij�l���?6L��C�tCV����*7x2�	��'ia�͎��E�w_5Z�>�2���Ɠ���=�ؐ�H�OW����uc�2ᘕK׿V�L�<}�=��Iʏ�
D�:-��3�¸�an�6��ڳ���!)6��WB��}��N^�/Z���(~h@�'����/�����<�Rǯ:�@��|(����� 'J�U�7d"�t��T�jOk�ԉ��PG���!V�cDH�v�]��2�LO8����?��	����M���O�f:���{oE��T ����,����!5��,.4��7��z���D�"Ԣ��Uƌ�����`�b�p�W�УP�LhԲ�i����}:�3�
Ŧ,������jȽ�u"?1F�+fv{��"[*��KW'�}0���B"�V+���,�Z�O�'0��Y��o%�t�y���KݪK���e1ܪHCg���餭O�DIlTд�P����[�X�կN���~�`�f|׿NL�0
_���B΃�3�G ��!ГS�Vݳ^�l_Gk�x&�T�=�:Q;V8j�x�7����j����^J"�P��[��<��eR��<����$;c,j]ˍ�-z%�=��璒l��	�r'T���VAT-}k� T�ǻ(k�U�fјR��h2�FJ�[������fP�65��B��vH���p�������'.e���s�ʧ?e�ܓб���W�]c����{\����mDt���U����4�G�¡3q
��7k9��>߷�Ӄ����������)��a]1���os� <:����Y�o��j�CR�͟D��̹��6x$_b��,�^��2�;6?�C����:�H�I��I<m(��B��z���<J���9Ճea� �i�ٜ/��iUP�~�>�eΨ�,�n���|���#��.r�R�&'׈��l�Ȫ�a�����x�P��o��� B�����,&��ݭD4��?��`Eԥ*�c��N�%y��`��"ެs��tܭ*����cb)'ª�U} �`儭��BR��O=措��Y�+�x�e�ol{ק����c��:�u۲�^i����\�?YI>��Y���|�j7���Hg�[�S��HÀl������y}h*G֖�d	�a֍0��rì�|�a�hK}+Qy$Xb��D'�|��+����֧Z��G�cn"�����\�ip,���H��d$��';C
o��.J�g�Q�K��f((4�M�~Jިj^��-ץ3D��c�܍ｍc�'�lQ��yc���4��%��=�b
��c��Kn���'A�T����J�Q0$�mMT0ikI���,}F�� ��!;+��4��hڕ���V\wD��&U-��������=:=�?*�G4�o�~}�s�ݎMs��s��栍���K�̩~��f��&|�
/���Y��|�Sɑw�uN�<U��S��<BG��@�}>�s�z�Ugu*W���}�^W�� :^F=�[Ҳz�i��T�B�u�V���ۿb�o�s*�)��`|��;�:�ȅ�E��A�(�܃�[���&^�L�惘d1Em��F�m�ߡ;� �F8�m�9v)U�c8��K�@�Oh�C�����8>@	����c��i�È	S&���@��2�?2C�	XZbc�!�2U���IY�ø�k^�6������f<�^�BA]_����#�:�T{�l{�3)t�m,j�e�� [��〰zET�ږ�G&�>��y[�(+8��׹�t,��Ri#8�014J;;e��tF�v_3��w�-�(�{�GɂO�'�s�4�'U�!E���[UH��8��]��>g�`@�OCo'7�	���T�Zΰ/G�e�xl�n�~s�X��E�/�}6�j�(ӟo�W��fZs�7c��P�K0Kg&�-�l�v,p1d!��c4"��^g�E��c�n�/0���!�XU?�1����@2���W�\/e/�Y�2^�#�/�����_��1�/\�Zl#̘oy�.,Y�A���`�_���Bm#��B�;�=b(�#Ю&�1�%$�r"1N�R�JPp�[� ��i��u�~�O�z���9RZ�F���Bl�� ��`
�K�8p�����ᕗ�sG��_Ϯ�p�1^�^��Z�њ���E$c,.0�W�zSmj�����pV q~�z�L>`(r2P:0
�>8*�X�h�S��y�P����/��8���� �r�`#�"5\Y�K{���9��~��I�QG�xb�-D&'pʣ�#�5Q���0�4U��{��r�j�����3��-9������p͇X�!�N+�f1
���H�0!>t<.4mmLhj�1���0A�?�+/�|�V�_���&�L3 �xj�~�V5-�S�����j b,�i�8��H�*$Ό�<�J�7��oǷ/�"l�[�P$9M����vLn�Ec�|�	��W�0^��_-e͔��7A8�iφ;�J�'�Y�0,(���y��Ϲ`�_����5�ʫ�Zc�ѹ�c*�`�^@)�}�F���V�����4~�t��0!l\(�����\_���M{+k�X}���儉K�Lib5.�C�����S+�n`�F�t[��:=,|�(�.�͐:N�!��������r9�\�%G����o��X���?XXփ˜`���{�!2����U��	�r�� �T��,s*m�:l�¼��+�!��n]��Zݖ�f4�<���V�Go��_	d���f̟�B�n�y�q��K��l�/�i�+��2��,tVm����6r�D��JX����FO�i�J_�R�D�9m��Dڭ�g#��ې�//���|����0���i���J��c��L����(2�uĻ��T���v�����v�\��A�ɶ� ~����7�W��{n?�{U�z�UQ(<�R�&0(I�"6P�8�H�K'��v�Ov+�`���6qs����ގ�o]"+��g�K~Ɨ�1(b��_&���Ea��mą���#1�QR>�l��p dxṆncTY��B.ʑ�.�?p�&�$Rp�F\�,:EU�d�U���la�UW��e"�Rt��m���� �k.�N���t��&M���F�&,D����$����㷣�{rܿe�f?N1��Y~ YD�-��a*���+e����Y�[�+@ LW�`P��jYo�1.O�E��$����޶))�^�p��Z{ŷ ���G���6r��"�FPrG�@:�<y�)I,C߫�%	m�1�o?�q�u�}5�P�Zp���7y�*SD)��x��&ƾ?������%����;���oM?:AN�ﶖ7�?���M����Zxz�J>�c�:��GP �{M��$.�y~�]~X�Q�?<c]iWp]����B���T��f~I�(q���w��_?�p?hrUͿ�Xi���<�肱�U���t~Kjg9���1���Yd��x�V!�S�����`߆�C���)ؠl$���X����Z/'D���������ߧ�x�/2�����Ѷ�[�I������J��5)$�VmJ~c��,��##��p5]�X��V�29mcD	�`��OµS�=����Y��;�<.{b����A�p���6�ulM�N�:a���f�&c@�k������9����P�b_e!������ϑf��${Y~f�=WR�8zE�ݪ~���J��ƭy�0�l�_H���k��`'$����2rU���R`�2p��r F�^�������r�x%28qdƎ����Z�l��T8�;���V�x��z�=G%�/kZz+�^��o��Q��ĉ��W����q�A3�����=>���=�J9��?�Z���C<�U�X���x! ��=�V��v��!��!s�*�@����6�׎�U	��n�� �4��*T'$t�8�æ�N����֕mz�l��`�������ʡ��rh�x`�A�c+�a���V� �hȖ��w�.�v6ڲK���T���0��z��߯�pM�����oAؘ���\���� ��$厮y՜嚭.V�Z�qP*Fc9���+8�AO�'a`(>r����w1�yN?s|��d2���Xp?��j+}�� Tx&/���ٲ�
�A�e��JZ4a�*��3�f*K>,-�#y�;�
�� �Evw�r2���ݖ��j,aӝ���8�:��Fۮc��e񹶜Hx�V5 8���)�el����.���Xl�	��ڙw8?K�Y�A%��N�zsL���^�v>Ǟ*�@�>��漾2&0�T��`�H�^*�����#+=�����,��� �P@�c���i'f�I#�r��8��Q�m��&�;�f�7<p�6_�bjSa��76�e��?��^0*��-��ʡh��=⅋/ʱ:K��v�l0/ă�{8�����Y���c-��!��O�m%�&%H�?;�;3{�|�H�	C�2�W�����!
�ii��Dx�u���;�_o
E�Ua�g�� r�,5J�{�F�Lv��uj!� �##`-R�l|?�[�5,ÌM��.�������5>a��Y� ��(Y)Ƅ�dJS2���qO���p��F �	I/qq�_��TK��N1�$�h�E�ߓ��y@��z5`c� �(�-q�JU��6,����l(�ݹ�x4&�7t�-��\�fwU�lo�:d�uo�"��������PR'*���u��w�������U�UY|7zx����(���
�t�I�xEb�pI�Z���H�Ω]Hj����_nfT�5J�*L���q��G4�]�-�T(��D=EC��%e̳,tf嶾�e�<U�Z����9pd�g�����ztz�L�ja2��r	lbBYa����m����u�0~��%�8ã�~a7�&�eeK�S^a���L��I�wc��y�q����:��؅�H~n�q�`m�-�~��5mT�>�.����
b����� ��=�1����k��N�ú�[Y�w>�'z�KWx'���2\�ޚ�Ti��L��7�F���O����5��_��7��O��(A�9��6��j�.\RӔ����&�� tnx��|�\��n��Hx`S<���kҥG��F�^>������y���zE���I�:�l�����(OjL?|�w)0?��������Q��>c�=P�$�2�/��B��>��Vr"���"�:��;kQ	��I�;�qN�6����.dyy����A�h��Į��:� 	��-~�C�o����މ��;&���� ��I*�Hn�Gɱ8_y���,-�(���oo���ڗ#��*�,�T����[�EU�E�a�X���i���a��M���iU �Wz�ͮ%�x�Y���Ob0��B��+�^�)�ެ�MQ�S�?�%BX�`A[��'�K)sI���"�b����NdJb����/7�%y��1��6ɳ8>l^���ԟ;ot�����	�v/���cP)� �㦳#x�R����p�[g�

��{D�Q)��D}=��;�Z(j�B�{���2nl �z�$L�̂S��K���T�����(�m��ܜt���WVt���j�$���B�)?���Df��d|;TYEX�#��r��0�:6.���)�o����lU+}������;\$��^ŝ�'W��7 �������3�/��̐�h���?�&���J�����[�P/T�$N-h��O�B�Ja��U]|(��ں�P�A<�����[tgD�(ܣ��]����C��*G]�:,d����1���6�CW�6f�2s>z�dV�=|1�:�q�0.�jŀ8F���^,�k��'�!�a�Kmh��F�ݾ�ͻ�FХ]�z���F^�p��@�	�)CIm z��6�T�}Lm�����p�D�+1�m.�m���x@�t,X,���<� ���.P�ҳW�ũX����e�V�;�9��f���Y?�Zo�XN���� �������so�A��=��	A��nv
% ������<�{�o�'�F�%�~	ޣ�A���%�kSR�p>�k�C�R3�V*V��,��mҜ�'lEw�jY��,J;��|X�槵�̠��3��_�0W�! V�\7t���iw�L�v�j�pnn+K��0o��/rʠ")Qk��.v�r�I$;��M!�Uł�QTI���|$�{}.��fǵ�a`SDk
(���M��FP Z�=D�kn��� ALT���@]��s���ݤ��HA�1*���Q{�h|�b����+��|��٩H����B)\+���g�H�R�S�2~�<��V�:oyg���+�L�c�R���^�6��D�7N>G�k�B>boo(l�l@-)�|`�Nt���9��5~9�Y�e��;E���Aq6k��]N��Ze4�bY����L[o������~����f����m��6x�jR�;�G hk���MK�Ux��Ը�$������~�� �u�z��� �	6�1�e�7�6/��T�1����8s�0p?r?RJ�ʹ��n�>��8M�%�U����,U��~�F�v�ӖA5E�'^����ֿ�5Ճ��鞨2]O5ˢ���V�����f��]O8x/}8���)���
t��h9����O �������dg=.�$@�T"�����hŰɁ��$�ҧW�|¥�̿����*��t3{rZ�����L�`�����f�t�΍��.����[�Zi�@���~N�q���!WaD�#�_��83�ML�����A86�kl��=y$Eo`��q&��a��=��iP �eN9y�j�,�d6�nY ��h�hr>x;=V���*��܉4�%�
�p�w����L��M^n,�1��]�5�����<����,T�[u��Ԭ�_i	���R�σM������e�,��@�mM0M��gܫ�s
���2�L��g�
DNg��{��+ʫ����LQD<�M��D�m5�@�ǧ:�O��uG}�Uo6�C򋛐�Ъ�!��XU`<�a`T�����\�������/WSM��`PC���M��"���j��G�{G�EUac���|�Սo#�V�JD��?_B��Pb;x����Uhd�t�ƂaB���Ɯ�
��i������Ҁg*(��Ȟ5��%��75L���T��М�y�Q{e�9����]C�?XrA�"�mz�z�:(���m�5�`uu���3N�3�����6y�q�޼�#;ӛ"S������.���(�N(�6�9�9��qX-�|����rw�\:�E�6�N�X���[���������]�g
+;��̝�t��
��rb��\��AJ�����7e�kfVg��jm����e��P�e_v�3k�lذc���:,����)�\2zH�ҳ�ɟ����|�\�\:p�nK-����	���ء��O�R�<
����N16]�����i�]>���9�eW�ӫ����-�����Lj3�ak���9N?Oڣ�_�]3���P*����Y��_������: ��2u�$-�G��W�[��u��JA+�+�Sx���d����f�t��1t����6��#�K/���<,K�� �&�C�ի�8J��p� �f��]�,&��6�g�A�-�M�1s1���Y]��4�0�Ӄ�?��`�a��WZ��w�#���[���Vu����
=o�鐯�G\H�?�����D��I�Q2៕1���Q�}�%`��r � Q�ܟe8��$��R�N�ª�ʐ=t�ûG1����*�w�w �D^u4��C�c���L,HP:	��h�H )�h�4<�������T���ڲ.�z�J%+Y*+�/��E1��׆����1�3�%π���>��N�J!x@�;n8���r-���b0N��;�j�n�`u� ��1��|-��q�y�|�v��wx6���;Oo�wɍ1';� �u��w~,���7���oQ����`�'��Q.�k�uSS��kc�m�(�&*Hi��;a҆`����a��4�ñ]'Udo�u崠dbrD��P����� Odk?�d���@��UB
&��nUkf"�<Y�q��������|�l���=qB|�F3�l�o�>�qȳ?�UWf�í�>�~h��$H�d�#��N_Cs9���'���
��X�5me�{lz�Š����+U�&�|@
b���ۦ����}/����Wh���_G���H����z�� ��ĺ���8��S�A�
��R�5��f�^%�'!�\�$d��KG��h��d�����q�3��;-�qp����h��g�Vۚj��j=�|�P�%u-�tc_�~�e�X��P)�h-���@�d��ݷŃ���˽zt3�S^oz�sC���YĞ��c#��aö�"�	�Gl�H�/X!SPg�±��m�-y��IG����iQ^������4������Q���t�֭��	�;�{s��y�����*���2\��Z��E\�2�#Z�����%xA�2vpFYUvl��Nr��4�-����VWM˭����|<ธ�^�5��g��9OeC`����	�^�N��<���|�dC��I]�3��C��B�2\���:�̂*|F�)e>xe�i/S���PS��o$(�<7�������D!I,���AI�m�r�n"�>k'�D	ߐ��摭v��iy,�.�"��>�X�y��}��pQ�
0A�ܪ����E��UtX�kݟ�%g��%�BZE�:����Z���>�Bk;#����z>�z��S㟛��a#�1©��=g!�.7�)��#B*��֡���^��%�����O�g(@��4�y=�����f�:��#�V�noW{�T#����c��u�@������=s�P�� ���,pۤ3��R���,��W���6/�&�����6UQq�Ǣ�hR�:4$V,fC3R�C��6�!��)i[�۩���-�8��$�7���n�&L^��Y���5/!����`�$:��S�fF��>���
g!�`��ww��[�J} v�\�'���9� �s}g%��u���YSI[�q�g��ٔ���ՁAB�R�,��Rc]d�b�Xભ˅�@*$c!r^��I!���
��@c��<��	^6qA�Ǝ�ha�C���m�R�|&i���HǸ�G��
Uq��hK�=�(�U����z�hR|����a�A���C#њ;[�����$�@�$�}9}�K��i��«�'v��IҲ�\�	 ��w��Xa�r3(a�P�����xk �L�x�]
Q�Zk\[ծ���8� !K��w�#}�ߎj.g.��"�sc7hE�A� �i�BQ
G�Ǌ�(���\��fn}�k'm�a�ke��~��IC�{l� w3ӻ�f�}'��pC�����?�l\�+�g `�iss���JI�H�p��P�0�%H)�jI�}���RZ�Qf4Zsut59H�-���o رT����S�g �g��\�.�o�NqT�`p����mz��ˣC7}ҭf���M������Rx�q(�Y�!.J�9�[*0GZ�1�\y1d���CS@���&J����м�7�(A~7�j��I�Ѿ�VKl/��-<�1��D%�d�q4nЧ��[��:+�M�,,pQL)��e���K�5t�⢕�n��)i˧�1e"�@m����E*B�,���ݫ
�GC6�SE��q�(�+�ͤ\�P&Jl��KA�8F,�::T�Ҿ�ڼ���cN�� ��xf�N*;i0RG@����x��X}U�X`^�����+e��x��U���L��5�7ΌimE2&ʵ]k$r��{/Yf7�UGQ��k�
���o��x�L(�-�? ���a�VP+�/��r��}E9q}Fe��MC��Jκ&B�Tj[>�I捬D�	�d>���)���3�V�婫]|a�v� �X�E�E�0e�����pܱ/�>Sɝ�_cX�n�K����(�>L��*�x˗��u�����=��`�|+aɉ�!G| |{D���Ygnݷ� ��
~��Ѐ��Y_��H}`	��Ղ�?����9 �O�~���^�63;!�M��4���� w+
����Ĩ;��h<G�=M-Ҥ9��w��B�g�/a�N��-s>,���
�!>m7)��}�����W�U�36��$�Ӂ�������A|}?(�<�-���>`�O{3N�5���r�-ƺjݪ��,dU�ح�[�Ç=���λZ0�ⒽY�>�^���+wl�m�^hQ�K��mO:�(��P�U�tV�1l<]�T��'o0���C�j]J�|��U�H7q��1u�Ci�!75��f���jWL� ��Yw�Y�ˆ�7� ����U��|A���գ�2����h;j܅������ \x���Q�m/<Q`Q&��&�-����7�[�����k��ܨ�!ر��j쨅Y���O��H��� �1��`��s3E�̦�*���c�����1�yЇ�'	�E�,�T]��[8ջ�lʒ���`v\9L:��"a���&��ñu�,I��}s3� ���.Yj�{>�e%��w���G�	_��ץ'V�+y��:��i�FGk�*�gΪ��������06�U(D;��v�n� �]�N��Q/�H'/�#��<l�9dV�R~�+� s���t�A7R�vѺ���j[=�2iJd�s=c�z�k�}=z.�R��?�*w�'��+be�X��(q�*��8���|]�i�.�:�K���I������?�(�79������K��=��A�$=�5�w��ڜ� �5�^'Rf=�SO���Y3�Qg�	W�.:
K��W���˵����m��ow58���q�gaTB{z�Ͳ�Q���CЏ?ˀx�y��!��?�֟�cV��
�ԑ�]�D�W)2I�df��"�]��{��7:u*?�5/@�7j���B� ���킮�$��qO�Ĉ!�hNlȋ3���m���������5�>Df䝬�P���+��]�@��6B�^bW��e!�ޯ����`��������W-Gp�]��rR/G���2#N&h2RR������S����K6��Xp���*媣�w<�#�m���ۦX�yW�Ϫ!���U���:2O����m�Q#�Ғ����	<�e�@��1�
��w�z܋�5k9|giB?���&��O8�ߢV���x�V��J����
4K�.����%Gw��3�΃�9|��}��v�ڍG���?��`�_~N��A�����Ч�������������~E��Q^��d����	;�s�>��`�춵��^jq
\��~Q���~/�Z��}�q��]0��8�t�9b("�l��bUw������Ai=j��T��h������N(\ [hw�;]'(]��^�=d��XoԦ
�C�2��v��)Abu��X(>G@ႝ	a������o���$�Y[}1^�7�?Cw"]u�f��M�� c�?x�����8ֺ���a�\UW�����{�~��*ų0?;�3��)�o(	�,��t�]�ÀpEyK�3'@}d��Y�7@:Q�*i61e$h܁��N�ߙm�ŗ@. $�1���~�LL{��I��m;�Ħ�r|���f����y�vV���F����>G�k%VG�q�u�sĮ$#Udp�mLv�һ/��f+���okm�nj��'Q�ፍ�c�ݺ7|M��$�k16�z�l>`z#����P�b�������t��9��L�� /��G~��h?tt�v�6�F^��<%����i��.f����P�ȓ������f�U��=c�Qr�Ͳ��^S+쿽��S��M�_�~�j�/��T1�1��� �� �5�'7scM[)֞I���@�3(�,H4�YTO<DW�]��=�3���N�72���B��r#݆�J��E�D'G���5��/��z�.+�uO��'M��yÒ8Vbxx��%m�"73�޶8��D ��\`�o*;q�+��R*ّRq�v��94�)��X�q%i1��:ϧJ�!�O��tp$�����-����-��4H�'j,������F�������M�Z�z�G^��o�����Ps��j��&^Ug	���Rb�.��"2X���Ю���`�U���r��Ҏ���K��p�0hXy���Q������X:���K�ьf�[Eg%;Hh\�cg0��4��S�޴��px����I�V�j$�@x�c������u���,�<��l���p񕒗��E�*b��+qC~Ґ6�c��Q#���B�`��5(����qU��� ��a�ֶ˳���M�H7�}ks#"��82r�L����HY"��ͮ�y��ވ�+��	�DǢ�<j���P͡���K %L]�̎sݓ����D�@0+[�2�-�J�}�V�3�@��|$��؛d�DC��J8�
�:/s�̥ �ʨ��\��|�!Q���fp��Zu�F[�*g��xy����et� &��oD����a� ���C�R��K���J�7���~�M��M�������������k�O�F��_�w��=e��z���U��p�ϩ�K����ͣ`�J&q��g1��/c<�t���%"��	��5t*w��EY�~��`�z`�B^�S{d���r5�T���R���� ��,����T�]r�!������F�PГ��â�و�C�U��Cx�-;��arW+�,2�_F�N{s�K�{&S@=����>m!��G�P]�j=�ՄGi��E-���w�/s ٗo��]��ӄK^ќA����%�
�g�����.	)������衔�mjt9DȠ�J��t�r�?F�g����xz �W5�����q|�G���Ǻ�΂�\������a�����;��"2O	A��US�)��*�g����c):Dc���\�[utL��"��;U��V3�Nӡ3��5-�<����/s�%Z���=�|�.�y'��Vd%�TQ�R��}x�=��_�ͯ_�x��������Z��o��@b�r���Lo"�s�&���Tj��)t�P�7��J�@p�Nm����	]�V�1�O&���A?��t_����������:(� ka�8����|K����#p�C�8�5F+�*����!;�Nt�j��[��2�{Ջ6$��_"PĂ>g6�n�8��23��Hgcئ����TR��kᜤݵ��p�0��Ϳ������ް�C)��B�)��c�����dt2?Tx})�_Y����7��m��*�1�L�Fy�	#?H,�0��	�����f˯0X�A�"��i+Țh0E���88�q«�طB����U���X.$	8�=7RAb�O�*_ ���H�no�M�M���
�X7t��'rxW0���$*��?�o�����<h,�z���es:�%E�]+�W����@3:�4dj�ㅊ����!�ԫY�Y���3m/C��2�&�Dih��L�/'���o��8AJ]_��R$I�$��e���']�'H����T-}�}���Ş���_���NAڂ�@S5D�E=�Z
tх�|E\L�Za"r���3�,��;�A�ݯ�f	���Qu����8$��!?��0��@}8Wu���gJ��>O�_�ȭ0�-"�7�6L�l�EN���"V��D62o�{�������Z�!{E-�된�|~�4!d*�O|��+W���Ҝ���p7���~���5�&3j�D"��|6�<�.��cb�u�k�����0�;�聴�A�{�����e�} 
:�1,}��$J�~�R��<ˑ;��e�3x� ����C�3{��8�9r��G$��1�ͷY�v�1���3e�㈳�`����w��y����&YΩ�.�.�M�!���Uy��
4S�Do�5�6ZC��Gѱ�B]3u��7:e��M4ֱ��aks�
{�E�j���X�B�e�Ka�]�����"|%r�w�.�}�R�xLT���hV}:�%�
�$ٴ�����|�<qÝ�K}�bN>LGm��.��b�C�	9B�ӿ*��VL���*����� B�H�ӕ���B��'ih^l%�	��x�Y	�E^$��e欇����S�LW��q/Ѧ��צyQ�����w�d�`dl����B4ǝ����.�b	�O�c	��坸9dK55,Ý}�q���e�r�:&�i6�%�v�J
&7�8i8��'��&fr���B�]1պh��fU	������*yK*��j�8�ꦝ�?qı��j��Ѱ��m��xr��M��۳��R(H���Ŕ���t��,�dH;6�Gh���~��Q-��H,��yGa����o��;�㌔�4��X%�Y�x�Z�t6��J��F'�c���q�85�S2в�?*�3St&����0����h0iR�0X��	��=���s�Ӡz�q�����`�uc�8	-�̆���B�-��r�U�0�Ҿz�ﭠN�}M���$8�*��)a���<���"gDh\�C2�-�X���\I�7��g��!Æ��k��84�'[pb�˿ �y�����*��|�V��*X� � h1��T��d{p����Dd�ibkX�m~a[߈�y.�D��'�4,�{Þ� Q���Y8�R[`G �6���z���-�;�Z��݆�^�����={��oz���r���^*����]<��9�Q�L����ڸ��[0w.���~���m=ᇿD��p$�O�Q�J��/M�'��X������ ȧ՚�mH�~���3F[A��d��^҅a?��L7{XYQ��T�n�մ]Ð�����Jv�l-a�z�%��盛U,�=��:*�:3	Ǎ����v�,�k��X3S@D*�by8�q���H�5��c���Ȉ�\��Q���refչȹE�DQ�D�QN�1D��v^�'��Ȼ^���'| �����M����-o�zo�e������͜�L�>�RW��� �?�?��	�D|pP�d��ύ@�2Р3���?u����WH�����dU>��1��O�&ܥ��t�q*�W�XlJh�M<�k����I#A��YIg^"�耧�Q*�Uoѥ{� ��GC��%��G��Slm�G���|lkz��%C4�M�a1λѸ�yG@H*���#9�G����`(R8�t�V��K�-uwy����n�)B)��ϳ	�hŬ��%u�&�n����2o���l� ���7�I8@���+PX�}��]R��L`-/�yQ��b�������f����{0�$��:���o��NcgDL�_�f�r�]"����+�r�oKN�:@��^��}(A=H�1�E{�3��U{_s>����]:��XH{�|w�~O���a�Z�����k�0��C|����f�y/r��3�ӆl���r�?E:��N6����В&uwtHZ�F"*LӂɃ�	�T�W����$�� :���j?O+Lx�
�-v_���7p����ŭG����sE X�סk69�����N��p���1��v���!,A;�T���`�ZA�"�]>�ʬ��!��$����ہ�4;37������T��'�e��@^X�rA���1��&���7VL#�C�ns�oU������h��r���]T�M2�.�7��(?U7e���g���޺��h,S�&M��;���u����\kO�4Gm_ҟK�̖�Z����6�oi�Ɖ�w�z��d%�3�5����ܰ 8!<}�X�~�̼9�b���%1م;����r*lu�>���m�k��!�E�T���㐄PZ��>��$,�ݡaXo�����59v`�F0����Bݤ����l�������|P�#�ƚKhr`�D�6] *��svY���f�(��2�g�_{�@��!6$����z��-Ìl�?��-�EV�sr6��<a��wa�0{�����[wG����Q����9Pz�/����[�Qڝ�����l�z}&@�o����=����VeC�nӕ����PFV�ܒ|��`��1��K,�{���C��]9��HCs�8�xH�e�Ѧ����ZE�3�sg沀Gt�nW��O&�j���S�G�,4���|�����O�<��l°�+�N���&�p�5,Ʒ��C~���
�Y��.�����t]톋w#ҭ����ƴ�$�u�\�-��R�̻��x���~$L-=Yt�LD9><z��X݈n��K�2 Ā�� �^�p�	 ��ˑ����r�t�dдvXm���zR5z��AIB���M j�z�60��a3�}3�ӱ!"�zf9C���C��I.��n�P&AOq�F��(O���P�E�`��l���#7.��"Y�J� �3���g�H�E�$i��\����o{�]Z�-^(�8��0��C�>=��D���<W��ơuhO|&�O�,�WrҔ��?�r�*���:�-/����[r�b�C�\�<U;��^��@aE:x�ܳ7�O~��F�a]��; ``&w���3[R�B��ׄ�4������Q�}j�fo�ĳ����Y�����{i���~ܨg�5��Cׇ}�@;E� x��}2,\����av8X]f���y�����eP���7J�T�Y������.�c8tՄ��P�̓�j1�vA~37�[6��&|��N���Fx�q�� ƨ��G6���po�+({�k�ҙ�"d�>!I����0���ooO��6�/���4b�W\#G�J)V���
�3*��g�D1�I�d"�hAy�l��Ȏ�\�/�rmll(�W!�c�>2T��Md�&��A����䃗Kp�G/��I(��N�#���H����7��������쾺��:���T��J���)4�g(��s� ��^L ���6|
�)N�,�
M���W�w���P�	�(/y@r��Bg��#�1fCy"�¶v�%��@q����+i�u������!.ꖴ�����(p_&�z�}b��4!�ZT-m �@��Mj��&�a��l���\�+`\f��FC��G	 ��"�d�D����C�}�G��?\��G��3	lB.LV7U9�����7���I }��Pv|H�.z߰�/�@'��2�e�f�W��C���l�AI�>��k��nu�w����V������B�3��d�(��2��j[��;�^�A����W�j�I�J&����{c=��_�v��:Q�T�[�^	 >���3@P�ʮR�T.��U�#����+��FAx�mY5X(��YͰF�j������'{��oh\S��p��aL�<����UhI��f�?Di�כq��T5�|w<z���� �L<�ߣ���tt}懑[$b]ˀR�U�z��9� ze��d����ׂ�M�HU�Ny���H��⟏�F^��bu>��u�s�����]<��0R�GQ����7%L�G�F���,��kN��,��"g��(��֘Hw�va����s�.��~X�u�*�Jl��)�x��3��?�X���R��I8�U�"��2ܸ�~Cq��Q��������lY�3�7]X���Z��s��� ��L�����	�kB�� :$�`�FE�u��{ ��*�	�	�eQKdS<t�޿�W�M9yD])q�"�mup�ur���ɷ�wˡ&��C�I=wiĭP����1@Y���H��u�R�ǈ�v�,3�r�:�^O�@pӽ�D��΢��(-\���8ߪ�SWx�3� I������z��;�C\�QE%&��+�������\6�źF���|D֒G;����1��2��"���pR�橣�:6'�i�/�ȗ��n�Ӎ�h\��8�sV��`O�UK�������B[�h��n�]5W�In�m�i��	�r@l�rɫ �)~s,��
���{�4Kv{ӂ�J==�a�+q䣠�`W�
��-��)�	�������3���,�((e���!��Uթ�|�l���R���H�k'�U�����6W?kf�/Y	�D��}����Ũ��F�x%��:[� .�
	8�"]��x��4溏���WM�a�n+gNd�wE3��9�o�S���~]a���ȍ��uY~�6�%�����Y��;R�K�`j����j�;�)�ї�0C���/�,y� ���CQ��5�6��L� O5Od���~	,*7���*5U�ܟ�[�1�-��R�����d��!
�
:x'+����{0�ɱ���J�Ƽ�l�G�=C,��~����߰�zŶ�q��X�K`>�Ŵg�汋�W��X��Pѽ7���G����EI0^ ��!eP��WGRe�醡�����%�*�O7�����[��VXf%���|�p�b ����(���13��9B���V��i`�m]zG�s�:��F��^,��y)�"�A4Г����a,�G�f��i}n�n5�NoL��b�pզL��0
��
͚�;�����2�n<��oQ��!�m��TQ��9"Ab���BW�2�UH�b��R^��>���#������O���h�H���wwv��	D�#R9��V�ÏP��V�an;���˦�Ǳ�WS�ȓ$�
�_RӁ���d485��1v�#=����7�7�w����]𐶫�jtn*����So�Hn�o]��U�+�{�����d�ј���!�@Ɣ��3��9Kc�?���)��w����.R�j�k��hⴛ!1TS�q*���9�b�lW�$.)6.tP ���Ǹ��3*Q	�N�k�
���v"M�c��ݓjg<�m�YO0цI���R�$v���ee�5vW)�Iԣ�X�?��N]~q|�B���_ʈ����5�[p���}5�R��O�>5���\����cմ�ޓ�b�=߅n���`���ч�m�׾^�I͒��R`�%S>��kZm�?�+�����8v����hW�����~�<��%��A�>.E��/h���֞?C�F	A=�*����[�����#�	��]k � �|�� ��`����cT������=��1�9?X�,��\�ꐵ8�5�4��l��_��m[a�|�5ml^�Ũ@a-��P�2� Ea�]~�ߐ.u���*�S�����gs�i������C��w�uj��$�C|&��LwU���pO�X��I��?��y��X� �^��M����9����������O�AothL�]ΙL����C������Kc�� |C��s�����I��M2�#�7���oM�Zb2�Ѝ����������i��ԕB�:������c�6�;I��r�=�"�YO��q͛N���������Y����]th+9`�~D8!�)頥���M��a3,[����0p6|���s0S+��,�+��,h�GU��N���<�X��ڃ���O(��
%��k1��N[[Z��wR�	h�[�*��I�ʹC�m�~X~�!�)6���`l�y:ѓNae	������ �񴳁�y��N�0A�P���bq(�E��ĀQ�X����6W�~�P�� !�͐c�&BI�l	S���?��������N��+�4���F����G�H��e��	�?����A����GX�G��\�cA��x3�3��%�)���*��q�<��M���ꀣpE�����ns����Wn��'Q!��@�.dZ��������ۤ�A��;]��U`&b��=,��a�5�
L���I]�AYc}D�H��|���]hR��~'װ�D}���W`?�������g ̜��a^�@
�Ǯ���G7(ݫ��A<�k+�Ⱥ;h��ǂ[�p�N�ofD)���c�1�։���%��4~��y�X����sZ�Ç�%Ȇ���$Qc\�!�k�%g�,��eVo��/���++����m�N�/��+��Z��j����-B�?K0Õ�;"
r�Oc�DҚ��ڧQn�b����C3{b�Y�5A�ЭX�._�SR,����>׬i%�1����dj,�Ke��*C���0@:���&'�fP�
��sp�䀱�����5턒��\>f��^�4�oB� ^�z���zc���
r�L���A�i�NA)�k��W�a=j�}�o���(�No��]�y����c��U�!H/q��Y�[� �5�`O-�D����rJ�>�3z^���E^w�����;nd֪d�JB��i,�ث�b�MMN��kK��s��w�~�7����B��ԍEry�C�T*W�Lc�"��g��/����f�I'e��]h؅�c�x�I�%�+�5�MQw����S���R��#*M���Ƥ��E�2Ynz!}�L���En���Zڏ]�~ǋ,�VL��e8K�'��nD�yҍ��?.��qd�
�  y>�;0�.&��yN��f����F�h��V�_ vk�Lt>H�3=,�/7d�i���^jz�b���52A��U�րN�h�,/��"�c��_����r��_�!OQb�	]�>|A�bf"�O�i�,Ջa��(��������P��	N���o���X��ED[���O:��%t<���*d�V�[�.΋��=�c�̌�%��i(io����>��ұ���p>8qϘ4�7n
!n	�'s[s�LaR��8zmv/ N��(��aQ�E�����P(R����2��������=
t��h4uŗ�V�ZҷD����d�a!}����u� 6h�q�ɗ������Ć4�������ߴ}�2$�V�^��r�n��C$�?c!�I�<Q}�Ya3e]�%2=�G�>�ӱD��~�p�!�9>I7,4���� L�B�牳�N^F|��5�
�
n~J�D!Ԣ���n�-���0OM1�"�ݘ"�8Y�Q���Ҟ����m+�g��ˢH?zܡ��i�b#�(�+���]4hTO�0|)=��mZݮ��|b�G�Kǈ�ܛ�H0��x��[����~G_���
�ڪ���s�a�xazȺ�/�$kY��9�0Bf�!6�P�s�q���N�Xgu������$?H�+��[��e5�%EI�|�\�b:�j9��]0��E�L��-BC�i��t��~m��t��~��W�-zk��9�T6BF@��giXU�4��H�X���7	O1�Z���:���Y��H��K�~*4�f�����VwYB�9�&T���H���=jIr�5�]�"]J`;�`�QCs&��t��)�M��W�C���G~tj�}����Ϭ>�ܾYcz��^K-�$�͠V�x�#��<n"�><�#�Q��kTؘA8� �����*��2�i�zh�G�ն�mO`?pP�35?��r�����*��C��RAP��rw��W��o�=�@���4�uҪ*cA8�]��>g���ru�g�G�����CO�"���6٩�@��m�#7C-"t!M$]j�W����0K�=���(�-���&�̈�*����cu���l�`d�e(Nf�����j�h�[�8��	�S$��#�_�����&�jE�r=��Q`qM)k�1B�ϲ`30�G�Y7X��!���n�w0�
̒cG8�u��~��5�I�evL�ps_�����A������)�1�Yl�O����Z�D�J�"&�T�.�����݉�(y�V�׎=G���>i(m��q�Nu�x��%�e��?[{��^�Æ����Й��\\���+\���1�oo���\�0�L������]���1�0�0�x����r*#c���Ĝ�#�W��B�9��ĺ��^��������.������1�z�	�E9��-0`�ѭ�5{_��`�ZLdS�����/�A=�,=�v�E,��"'�YNݨJ}+�nȷ\�4QD��Hj6&n��9$�ȋE���� �p�B<�,g���mWv���D��	�����n��p�l���h�;wTGg�U�	l�/ntk�E��%=Nq/No�'ZETH�U)��M�7���*�C1د3�Ȱ�6(@ТZ���A �R���N	��ƊI�7D�{���d��)(hR*$�rBÕ�a�a��%����͊�
���Fj]�8���v��}�Z�xI�h�M�?�3��Ad�����V�z�?�׳Sp��G�l�5�E���w����b�ّ&L��Ϝ_�{إ1�^<�]c,�TC��4����aٶCN�'�D���.�>w�vm�����u�m*��_G�~&�� a�»|��y�
v�)Ĺ�+v��2a'��N����y�G��N��Mx���������3����A��4��O���g����h�8��C��N\ҪTAJh6��$��w��[O��cֻ�'���<�T)�yx�y�y¹��{�eI��)<%j,� f�G=hi�� Gq��`�K�����<�����	���� s��:vKs��?���F@�j�@o[����������5Z�[)n �6�E�pT_~9Sp��k�,ܽ��}��;�?w�L��L&q���,�A�A��ԲV��jKyt[ˀ�'x�Zo
�Rzj��m��s(XNU�*�s����{{s�kr@iJ�R��޷�pyW�%��l�*�!��7���/��Ҽ����J!����p��z��R���,D��;�ԗ��+�A�ȶOfZx�t��LAGvk`�ǀ�6��>��7B#�>�"x���'(�.P�^�����ɱʊ'6�ԗRd�B�A.�1�HMr��GS�K�gk��k+G�ɺ�9�_��JLrV�B�v��-��p��#�5�={(0��&�(�
P�/�#?vy�BhU$Q����&R�VZ�p~�ZH�Mg����%?y���eFQ�ޑ��o�dÁ�u�_�[�QS\�N"/�{B�^X�s?̏�-��Uc��Ï��`_qL��&s� ʼ���V�RG��j�ŉb	
���Rb�g(�f�9P�XLSrF�l��xL�?+��mH��S��*B��ܵ>�O�Y-/�Ef����)@�����tF�@_�"��ƿ���Aǥg���/Vƍ����J��7�Δ++Z��wZ�&�O�S�q]��P|����K�2�'6��Z	��� �s ���T[����^��ꉪ�
�-3��;�<	�=�ܒp���v֋	D��'Q��m${����b{�R
�3�jݘ�*�Ӟ��8��[y� ]?%��0��'Z;�}��Ɏ�}q[�ӝgbu�8�<��z���levt�Xw1H�n�g;�al���
��4��>��n��
+X��l��rm�.�#�����>��u#��c'������H��˛s�[@�@X��b	k�Zr��U	)�� Qi��)L�s�CI���$՗SF��?�	�jfB�����`K�9�ج�QLT_Z�pO��\b �0��������ps��c�Ii3�v�Ô�)��H��p?��S��^Hß��"�'ڕ����Т�����u��%�R`�?���IG=ƺ<�xZ��bڅ'4P����������<��3��q�b��%��*.���*H^��4@�u�sA�'E0�怦ef�z���kx���J��s=%}'�{�7G-s/�o}��c�|�ۢ6�Q>�����G��McZ���s��;k�r�2w��9X%2\�O#�fPS�BJV+����u��Qx��C�V�:l���N}s�X�f���e��^�t���ĸ7<��ćô��K�5܈O�{J8�V��_=	UK��joi��h�A��КV�r">�����aM��T�WQ2�����rk�os�a��4�"�|�;�ݦ��򗦕��q�E�tz������KO[��^X�څ�e�#����'��L�w:�N�����Wk�]���32[%`>L["��<�������F�W�Np����\�9qE��[]��{� �v� �ӓaq��<i�Z�3U@�����RG���	}�|��}�#9P\gq��D��F_�<����ru�-nղ>:�{39W��g�G	���f%Z�OtAm9v�j[��|�\�;��R�c�_:��O��q&�ҸT�Oe�<ϏbX%+*�g�U��߻�-=h���r��# g�L��N���H_�p��Ed���ܮ��~d�<���˩�j�����t<�
d���6�����0�F����#m�fC��Ёl��
ި,��JE	����'N-�U����W�}���#���`c���J�ů��g�\B\��s�R/B.���8�v�OO|�.&4t�⟐�5HRن�/�=s%$D�	��T�Q�����	5��^���^YTt�� 
)Iy��}G�(*�8�>/�}ׯ�UŞ���9A�td0�ބmh1��uE��uK=��#�aIw�+��};�@�0~��� �+SB\�R�0��L9�W[
8|wTȂt$���x�^���v�F�6	�8�C���`����i���������U֝5����7n�Lx���U5\?�=�5���9�X*mScC�*�5X��G�S���Q��dC���ꪮ!$����'�T�[�w�iZ�o46!t����"��{���GX�#XZ�D�x۳���m�k�tǋ.����_+��[s�c���Pa���7�R�G�1���,��G�X����e(~���Ϳ�e���+���]-_����3�Lܙ)���-۠����'��*H����#�@���g?�X��L�Ő|����#.1%�A�w'�u�l��<����i)�|]f7v��	��q��.��COa�1Sď?�e�����|�"vN]��z��I,'���&��I݊�yXF?��|`��n�6W�taD�-�h�vK��V�܈:ǻ���D��Y霷�d�L�j�u�t2���7l1s�?�F#6
OZJ�u�v�f�`w��1���i�,I��š�GE�8F�c)u�{�Vɂ�[Ũ��c��1�L?DY/zx�U/ŧ� "�,���,!~�.�'���('�ecч?>�Z
�l�>}���g�2Ⱥ�·�������f���xNXpS`��$�ͥ���5n�)	�q�Tg���գ����n��ϰ^�T���_t��1���X�3��6��4��p�*��4S�n�zW���c��-��R��x��v�k��!�L�e�:W$��|�����X!e~�FEY9*���r��/�)䡛}R̯�s_y�[.˽�(���t��Ey�{��x��a^}��I������n=(�x,]?5���<�C��!�^_�>	�($���qy�M�f/��x���f��$P9���(�<�2��>t�+����v��	�>��<mMۖ�������W?0�|��ʛ���a�5�[����u��e���K��(�s&}U�wF�Oi���w�&y��I��h�Q�y�&�qC�TF�J�(��g��-�y�S]���T�NՑ3���,����e��,(��ȶLP��	d߮�a����Y5{-��l�h������K���Z�ߌ;fB�٬�-}R;��~ȿ���7�o���~�Gb���DE^3jrOߨ<������eyH��0a��:������1�G#��U*:����>�@�#��Y��J �q_a�w�QO�$�h-����i�}��d6�P�m�$�Gt�3?�����yaԸ	�>6�n�����p���`0ȍ��N"���=��K42�C�[u����3���i7B<�
^��]���������[���L=�A0B� ��UT�T�[`I��z}���N��қ������K{v���VG�; h�X���q�,	H�aU�[��}*�yg�a�qF�mD,��Gf͂4�ls뤹����rv��7�����(���gI״+�$�sГqO�2�0�gkM�{��J��~�=�w�?�^�' Ty)�_u�a�� n� =20T�V��0uZGb��_�V=�0��'��Mh�J�)X:�9�1HpMn�eKd� �V,!\����Ķ�G�|�d0�d�Ɨ�T�|��M��w�#�\̬u:.^�\,�[.A�t����0�q?!&a�����,�a[�b���2�q|�k���B�uҀ3��EV��5٥>�*$�m��Y����w��}���\<W4�<]�6h�B��>����BtѪ?е�����I� W��$�(l�Sak鸾��o����r$+�`�0�-s�̓�5���hˈ��:@���9�?�';��9Q�qT���6@C�f@f����s�"7�߆��mR�D_'yc�w��-�CT$�]�4S�U�w���}�w�&�4jN��	+t�;� ѧ�����U�e�C��9�я3~a�6�B�����2=N�י����f������͟��Ĺb�*2��S��z�.؛�'q4]���H��R^��v4���0D�Y�	���^���g��{��]����~7
���.~lK$��r�	�F*���Y�+����g`gF�C� �p.e����r��)}������E*+��xn�1���; �m������4[�J�Y �t����9��k}z���~�:�Σ:W2D��T��ֈ�����pI%#B"�'���TVa� ���2�� 6�[7i���A�ܼ��X;U���J+#Ƕ�Z��N�/�u�y�%�QO3wwM�Ai�j
9;"��v�!ӹ��<����j}���6���xy�+��z���9ɜ���"ﺢe�@)���	pjۦ���/��	̖��3�y�?���#rI�w�8�1��,���Չ�j�BXC��3W�f�v~^_;m�Lp��Aڎ�����s����cX��q��ڵ�HS۹
����&�Y]�;� �C=ʨ�aw�+~��#0S�Ya)���H0�֙C�}�$���$���	��sm7"?�!wܗv��m�:wEio�
n�|V�o���e��
0+��M���m=����D�G�	(����dM�ӕF�;�ӈ�~�y�9u��th�CRBEU1���MI;���.S���e��SY�{B��?epG�$-�9��8*0,�D-J0�T��xq9����!q,�:�{jBg�D3�ŋ�/���7_��(V,�yA����u��0����4��\g���|I�� # 
o!zq0��(�
zjm*ם��;�''���Iv*�0�F���ך�6U��1�@�H��#�E�P��H
�m���?E����,t�O)���Cۗ���uի�u���^��I��M����:|�0��v�����@�sك�Y��%Ap�̜�	IWY|n�{��F���/\Ԛ.�S����؍M���P��8��*��I�3_��ԓ�&�Ro�]ƎT<����Ho�Q�u���=ce�>7�+��8��#h�1ԙ#�+L:�<��E�aG����q������զTc�<!�[��u֍�l����	�,/P�a�*��	VeTf�0!�3[��z�L9��7�ٰ{8|n!�����'��9����X���k��K]��*O�^��Z�C@��V��,D	���n�PCQ*s����8H�&��5��oźq�r���8��~.<��j�\���̵֞1C?��\�kU�=��F�F1�V��t^���T6?Ns�%�$��N�<B[(��Փs�!�Epin#T�6�s�.�EU�qv%�m�pc���@O�״��Mc������Cb�D��߭}�vζ�H������k��2?D�2�P�6��?����
��~��j�K7i4��Np���$]�k��GM"�T^���݆�TNIzZ�7;��l15��zݳ�z�.��SXm��2����iH��?�У[�p	w��=t����Ʊ��D��y�1��eŀ�59��@Z"�DTQ��jK�C��TG�J�G��>���4����'��^�U�/�;���4���3:s��T��@�YD�8f3&X�#�y�j��V�p�7#lu���-(I��~� S�;|KϘϬ4A�E�f�T+�X���z�a`5&x(�cm�[���y{�A�������9�	E��S������J�*���P|��K�C�cK�+k*�g��΍tњe�j�����t�o-�;U��Ѵ^bj<8���&e!̍xA{�zӉD�m�-����EZ��{w}���$<�jIIn�O��
�}��6�%G���ɥUCCE55c
7��,��?���%�Dl͍�"å����i2�c-_���D��u��?=i���	�f	�L�-�׵r�H���m� ���>�����hʖ"U�����u���&�9 ����(譂0��M{X2�'
�F��U��ޛT�~�Q9;�s�6��TTT9e������N�Zu�8�ڛnaw�`�a�S���`�Av�`����Q|R0[t�l;*��)�
X���x�6��CB"��6D���Ӫ=u���@�A��#��7����	K��cvGu���R�ࢅ�>>b�O�J�D!	�2՛Ir��ӫqj~�w�:��(��qC�w�pe���K�|7U�/l����"	0_�3oI)c[�\��-d��YyF0L1�Dؿ�|����ʚ=���E���N��'�w�I~>�w���`�E�b��\���6&:&zY3ѻ/ۍn2��<�F!)`��H���%���>��C�K����㠾f���D�8I�5��"X����zc�B~zȁ�>�#�f�
	:&r�i�$���a �Gʩv�J�J$H�&2�(�'�e��g*Kf0l�yJ�J��!a�I�g�n��]#����`���ڒ��ɮ�IT��&ԡ�y �C��*���Ul�b|�ǳ|�	d^f����ߔ�!�r�%�Y�V�����>�;������A��*�"�^ۿ\�=�����G�y��6L>�xR�����JHQ�9�G4wϥk�jǶ�%8-���ƻ��6����r��HAdf�[ŁSW��-f����l���6�Ozʁ'��X�ך�IR��BWӹ�8��O<���x*��nc�?�|��ٲC��' x���^P��"_ֲe���1cG�W�Wj����v{�+��=��dh8ѩ�q�����أ��i��:o�ؙBC_�^�ZzR{t��'�����	�ΥQ����b�sS���F�:yl�}�S��7�D`�#ҭ�S@{uұ�x�|�iv��.��Z�I�r�G�3%��6�<"�$�x?�8�ߝ��ԇbX�')�U�t��g��5|�h�=L��q1( &3u�n�X½ե�m����O���M���[�m� -��չI;�7�@ X|3U!���&�}�M���n���,j��v�jю!X׃(���8$z�S�%3ޣ1q��&}П<+��B0�yo.��׬�����oZ"�����
�&�g-[)�=A���	��8Ȟ��/����\��F�+%��/�w8���=���W|j-0^��>2,]:[t[��:�(z*���&!��p`�v�4/��2C��yb���V���v���&f�a%L\v^�8Hٌl�bi����)%�}D�3)���������/t �Ԫ7`�~[X��(�s��:s=��l�G�V��`쌖�4B�kz�}�/��	�8�[�٣�P�Ȣ��j96�E�5v*�c�j&/��"_Z��M����#���\ԁ�B}{^'X�u,�	#Y�Q�Z�Ӧn/lޘp�-b��wC;+�f\�rZ�f���M����vy��᧛=��t�B�~��H/��i��l.1�A'L ��)��Ƭu/�� ��U��D�����oXF�7#���r�/bK�A�?���d�ڧ�-�N$���܏.���]�!}�Yr�_O�22'����Þ
���yO�²�_���2𪗇��2(�XDJ���s�?�V��:�4�K�i�qB+��ֻ@ZRe���}wB��&����.�o�Ƕ�J�'(B���T����>u��y���2��ʫe
͖"��t>��D!�_�Y�;��-<	
�YTyDc���=�\W<�J�Ig,J�nϮ��:n�`#EH�*gf 3F���D��e]R��>�k#���}t���Me��;�Fz������S��&��|�Kˢ+�Vu�ۚx���Ȇ���1���c1P�ްv>�	U��f-��t���  ��Lq��B֊+?�@{pջ�{*���~U�z\Y�a$�$��=7Y�x�k�7�6PP���QV��k�O��Cq)��
Bf^$6�h^Br�{�R3+h��;߹D�7����O��a$΢�	`����~t�b�p����m]nh�c`_������G�D�
�;���h�&��D���Β��U�FovY�0U�4�;��[fݸ�
���;X��� ���O��k�`e�%m;֯���*��_8Ɇx�$&Vtu�d)V~����s�ĭ��h�� &�	�k�N+I>������_I�E�N&W��|m>=NS����uU8�򐙎��-4��F�e.F;ѵM��;���Ae-r�[��q Mm��j�����V�'�����������ܙ�>A���>g�1)��GTL�j�&�3��a̍z�4�'w6���{�m�Ԛg{�^��@Y�$�� us��5c��������U�6�%��q�Q`�rh�:k�̅/���ۢz0�E�B�dnƬ��*݄T$�9�c�_�3��'9	W��A�kR���1�Eѷ�R<��3C+�ųI�V��0?P�G�b��4��z��	X��q�R��pF���
�j�Wmë��8�	 �(�?�ݻu����^�n��~ש��~���g߬B�.WmS΂'e��'8GQW���ȡj�]�x��&��;�߳��BR���� M��t�<�k#�?Du�'c�xR���W\M�o��}��hs�_�c-8=y�.�"�����bet[���J�U�J�i�55�c=fp��.�,�X��`����**��9ߑ-�g��_������io7M�sZq������+�[?ڵ���ҿd�ڤYF�6�^��`]`������$c�n���q<N����!�S�z�`2�"�Zr˗�����O�W���D�@��:x�[�^#Wm�r4�D \�H���$,�XpW�0¬�����n��:���+ g������A.��s��(��M�O~<���\k56��,rA6:�܄D.�U`i���	EE'9�M�pR��L�f��jE��2O��"�F�C8W((�x�\:��z�Y6��@����"�}���knb��{�n ;������T7�KG�y]N�Ѡ���V�Œ��ie�p�_"�,�B�h1����$������^�`���z`1��7�N:��!�v���D�Y�pL�<�4����v #F��3�d�J^7-Զ�����$T^��x��6-J�w6��)��C,7�B����eÂ�����ľ�R�'j�:��)!LW`��+ӣ������~���D��]��i� 1�q���Q9S��x�q�����vk��{ntaux�?O��H$���p{�򪆂S#ҕ�!B�Y�����)^�4C�W������4���"qJ9����iq�"&
��8,z�����r8 �n��y�^����]��,�s�%]O��m�x'Vx&�Ps��K�-�~�tM���x�:=1Y����<vݤA��t�qK��v櫆p��~��Wd({�
�wv16CM
+4����u3[�{3�`��U�.�ݶ�=wV�J2�6�m����>���xN�����#J����JIW��9�� ���R������T	`���#��g����J��H�J�#������>=���o�b�3�-�` q�>��U�������~�%G���_����h�Q���Z�������S�cע:4���NTއڇ?*��X��=���չ�~��]�����96�(���,��&��.�et��:����=�v����q�2���u�32r�n&�\|�f���LB%ܳc �$Ӫ�������qo�r� P�~��ǘ(ߌ���5��1g�!�X��D��!��r��˂�H I��>�\hV��$ 
����=�l܀n��,��b��-c}�C��l'����ua��H^��tb�������S�^Cf�	�e�B�*,�h����T�(p�,#qq�劷���Y<���Cv�<��ַ#�c$~��.�}x��-`�\�I�'��ȌQ����!y�?�_.:�A���&.��Ѻ܁�2tP|�m�b鶨�uHYך��U/��/�S���]w�%��aA���J)�r���C�M8��]KUh�q������9���9h����?>��:?��������bo�l�;��Ĥ��y��"}�Qf~�p���I��=���>mV8d=�5tE�Y4}Q}u���|]h���BO	���*��2>�/�5������^ۏ�%��	�S�%��'�q�9p�R\�!�,4�-�no�{ ��q���fh�)�zۻ_~�E��C�#��d�h�Ӑ֚y��6.��ƄRKm�n$Bp��(���~���ڑB�zw4��Z/��Qe��3g4���z�ׂ�������K�q��g&�0B<L$�L�gy$Ol@3`�6�H2�Pf�U��X�qc�:/�u�CNHl0u�w��|P�"���&)�c�����<|x$�W_�Հ#*��s�Տ1y�Q�x>}��֨8˕h
-+��db���_�Δ����;��d�=Ox����6Ť�tCa�R�j����&y��v�3�-�܏�CW|J����ᯀ^��lE%��J Ѣ��X���+'F11�qj�3����T�R�y/�N��Rl��z��z�)�b�� ��T6J]��x�-���;����j�F9+P�C���fb��	<�p%�7E��`��E���n3�@�(&8O*e�ا`C�N<�Y��N�\�B�J���5�b�5�H\�`��G|c!fa��*�Yʼ�s�6k����DCv���em���;���Q␿C0e{4�_w�9g[[��D�2.;��;)bۮ�o�������	b#�լ�W�X�A�~�A�����9��S��d����hj_0�a�m�kMz���q�*agp�r�'� ����<�
odypn��������;U`������k�ca9f�,�G�/붣�H.��B��6㋇�H׶��Y�`u�U�N��$��M@���Ok����H���_ؐ�}�nP���]����zޒC�D�H;v-�TF�w>:E"�(�����H%����4vE�b��y��PO
aK��s�?������h�-l�H"�2KT���ۈ~�EA!�w� �{B�"?_�6K��!L q���j��h�gV����D�?�n��m$�����PִfU�R�:��P �L�;+e8�h�4���2�{���(�P̶�Y���H�f��F��k���~g~��.�f;^�T`�Un�b��
����SiD�Ӕz�������6@	sM�5˭lC3�a:�'�-}R1�l�:��=�!'wi������xb�����n5J^ �\ �s2Kpl�i�W����	wgfĳ���?���&k0����һ���b������L���������d�/;ͯ�T�e�M��1
�kr��Y��A��"M߿:˯6��2�p��
��b��7B�0�5M�㕮�D�}ܜ�#��7�,�û/���2�Uٔq �}0�w/%gM)z=�r1K��_A
[�s ��¾&�F���9GS�3�@� �
1I�D�w�z���i�~�{
����h!��%�q��O6&/��,>��k��J?p������!-���T[(m?���p�Cz�2����=o�_4��ķU���S��3)�B��E�qL���]��R�����f~����H�`Z��)N�{b&x�4��9��'��fH���;n�6S��h-P"��h Ä�`�Q�A��V�J�n"wq: ����Q�t0*T�o���Rԝ3�#�}��;���׸7�i�P%/v��*��?#�����<�� ������Ca�aR��a\��{�N�I	�~c��GQ���Ը�:߀F�y}�Tw��^t��>EK����{��'��[��K�x��҉8l{��dM@�����[B���Lmgoq�ҭ��F��p;n�%DT����˘;�܇�[p�s���>��n��C����F��h��`x^Q-����5偁����G!Ѷ��a�Z�4��n���J�����J�] ;^M7/ȥ�<���,st�����flR��q���y7��ʎ�Oq�7^�@RUi��{�����f5Y�X�m��?���>��E�%���5�Ȁz�q�38�J]�����@e�(��7�~�<`���n�m��"��b���2T5K^H�,�0��U�)�ln%��3kd_�L�+{��CТ5/b.N-�*=jC),zy��������zD[���T��ǿ��u"3Fn
!b zn�=`y��yv��%�.�;r U�b��e.��H}�*{u�����t��L�j�VS�LPv��b�5Hv:3~.�<�r��aV/�5,�J���:�5�4: bdh\�H,L�\`30@���X}��p���G���@E���>����0�����x��:ܜ���8 �[�ּ�y@|���Ma!�(��3~��֋�@��vq/,�5�䈏mQ�����6n���[���y�ZԊF�!p�~���F;��K����v%�f�c¡S��z��7�p��;k	�W��;˪:�VK�0�[��-�G��V��S,�b�� �|�$���"�E�V�k\i���/'�G-�w��=��0��~��t��a��r��}�\P�t^{�̊� �D�"��U�c%P�q^��"�5���@uV'�vH'�� ����U~CpW��׼������I�Ȝ��!��ߘ���V5Յ`�([�e��Lw��6���B�3rEYx�tTFR�p�)Uo�X�7C���
��LQ�P3�^fj�0�V��^V�$O�D�]����'V��S�'I��a��:��<�A
��$��/��O�� ��>�KL��# \�/VK�\b'<���ﰃ{�5�,�l��g|z��Lp�Ҁ.(/�U~�����=mE��]��@�G�V3���	ֺ-W�}�#G�n�z��TPB��e������
����8Q�F�<�%y ;�ar���V��P�O�܉����N�D�z�����RN�]H�����Mѽ�'�e�����!��p��o��yޯٛ�����7���[
%�h��;��4d~�q@�kL=�1�B�-�0�����3��r{eb*ip�z�p���s���*H�非��1ZK��ӊ���~��Z�� ���\0�d2x��5���#���������?f� >UL:IA��e��Gm<V��b%W`�Ǘ���-7	u��f����R����� -��j{��1�A������\���dO��>�u��j���:hn4�V��������#0e�/��B3��͇�z�"����)�H0��S���9�>���Om�6�D#"�՝N�E+�ms�� ])���b���X|X��S$�q6 ���,�:LxA^�@͡n2��u�u�ṇ� Ȁ�� ��$��f#c�Q�Jz�0�^|Hc"5�_O-��B�\)N�Jj.sF]��i�hD�vq+7E�Gdƻцo
�tڑ�Bg5��w{tb�M߰G������I(�H�2@�����%Ϻ~����KM����%Y��I0|V���<��{��>nl��W��.�U"��.n�������5GX�������'�ڮ�����DB٥i��V�H���Co�{�n��9�\������S�(�mk�"�h튁�A�
����3�X��(x%�=Pd���Ld��	F�,52�_-likO�� ��R�_�"�~|B�T;$���=��`��N���a/��].N����Y��P����Ἕ�-���د}�2�����L�q�uA=|R�i��H�ז���@���.�
 k�(=��E4��Ks�(����������`�X�,�2}w��uq�bx��n���%��l�|���R��l���2���^�rq��!�C�E4��z����ꨝrf�s����k'�T]7�~�|�d��%z���D�|�|BҢ~�Қ��#�5�qj`��OoIb�*�e���̃��'�t�:P|S�� ?���P�ٚ�y���V�$;���`7��!4���s|8�:{��
�L�͐�l�(5�~��JD}L�G1�2Y7:���E.�x)ĵ�-��KQ�rib;$����_B�7fy--�>� mq�T�$O$3+s����bڭ#b����xZ��f�� �Q��ۘ@qVr�^����s, �Ł5̡�	������A:m��RA�����T�qf�8`�s=R5��iEo�u�����r��,�I��enೡ��N-�7ʣz�s�g>�](�bo�*
�h񩓹��ñ��b)�V>o�cn؏,̢Q�x�P���]SH�	�M\����f�||o�Wlf˔���IC[e�&HaN���}mٵDd5Bʘ!A���MQ؇��w*�L��	���g�$T�(���>Λ��%�b`�#���)5�;��*��p�5WK-�������Ϸ?��A�H���3s������C�: �3�-�������H/��ӻ� Ib�r�1��tʤ�w�!�����m
��L�Xa�U}|NAP(\��y4�6�g'��ڌ���>R
LRT�҆���O�qK��vČ���=��%�D�:jB�2kV��|��X/�I���G>�E3��]$�$�|;�o��������iB ���<+�֞w��
'ĝcb�us�V�B8��~�T|,��og};{S&��b�1T��H�L��['��*~LRyI�뒚�����Ɩ����sg�M�H�"�����F���+���Ί�����WE[.��sR��	=��p
�u�Ԣ<)�p U��SL��#��U�j����y�t�U��q �@ �#���	Sd֪���"��w�gJ��M)��"���O
�>m���璘�$���hH�G�l������*�J)M�]��WUPT���Ϭ�~opr�����*q�-�&��[R",k���";g~\s�Itd~���4<�e�"��*�{��8Rg������	*p5t[(h ���*`@���R��1��gP�����8���#�{��N��½�Ce��ȥmW������Ha̘"���1�j�]�4�3p��X2Ǘ"�m4�]+/�ٚN��6ЉLB���[է�n�<��M��Y@F�7�z�ȍ��H���B�F⇅<����J�Q8�y>O���M�.2r)TslL�t[r����P���y�|���;L35���S(���M���0�%��c��%�  ������|:y�e���B3*��L5p"����_�̮�+ֱ��eHU�AY��A��֞��>�(�4�
$��|���hg����ϐ��G�3í��bL�Z����)�d�WD5+1h��]�P9mN<�IT?��9j��i�{b�	�;G t�qg�N	j�t�zCOL�{�b05�	@����@,4��!�|tȢG~_2�YG���bvf�ZSӁ�1�P�iT*�h��+�:��[\���3�Cת\Y�\�=��g�v
&�C̡��A�&*g����%�1/�w�+�X~,�%ȓ�Q�����c�t+:��cx��Sb�@����FT���x������#;����61}����0�
�x���F�ry�˩K��Uq�|`^�_6��5u�����^�+tU� k�e@g:w���k�~ij:�U��x�S[�k����3���.� Ψ����M!���E�~��~����"+�`�M�?t�(m8�մ0��y�@xkc.3~�� .�����u� T(���<����ğe��=�����>����|;C-�KyA�*�3�&�̴͙ '�-��L9�Q�з�k`��c¦��&�삝x��C��=uy��l�h=�oa��Ed蟝�⹧K�/���D�u�=���h�w~g@�6���)�V���27�L¡��0l�����h�g�t�� ���=3g_���Ք���A�-\b/���+�ҹ������U}qH ���dZ�u��@A�vE�9֋+ЉL������6��l�h�D�cPV�<,����?5�wF�!ñ��"�� f4�ɑ ˨�Z���W�b8��+���N�&�iV4}�#�X�lC�2g���u�zt/܈��\�թ��b3_u_Vf�z���Zx�c��D-�z�TK������>!��<�K�㓼E�l�v;��ȇHV������	 Jg�;:^�� �|{��O��ﰾ� :�H+{�-�h��F��E�_,���/�Φ�FXI���87�^@�S~� �hv��i�ؔǞo#$��o܏5bXC$���@5%v?�k�Z躈D��sr)�_bX���� �u���j٭d�͐a��f�	d�U��
����$7[5���D��n��i�]�uƇ�� 4,R��G����<�c?,�^U@�!-`VXLx}˸�t�1O&���D��>�ÛI�������8�=�yIϢ��&F���K^*�1���dCVd�j�T|�tܾ8K�H���h`� ��Tދ6ϲե=Κ�=$7�?���+�[�O�Ձ7H%�N��J����
��3%O|p����8�2��%��-��xaL�a*��cn_�Z��j�ذ�� 6�����Z�no^`�^c�|��h����l@�q+�q$|�ė�ܥ�K�F���w��M\�a���,ž��cm��ݯ�a�6V2��f!��h|����X�3�+GN��sW��t��M�?%Z�tr'ۿuxثl��I��<��𽫡�hu<Q�0��ZL�:!+�8�s&L5W:���c��'���t6A�(��}��ǅ�)��زG������R����y�8ۖE@�p��k��m�R��p�MA@+��OҕM�m��Q7.eT_�ճr��S8��<���쏻&g$��ȣ[@�m�1�VKM��)�m��Hh�ʚj͜�DT�}恼 ������	�S�u��1O�*�)x3U��`�{���k��,�Ӈ&r���,1,�kn�O����O������,f[��;���-����@�$@{V��L�d��������m�b�R�������rr�Zy�W,hw=�?��M��p�
�{Sl�����H=�h�@�`�ݜ�6��aPU���,��%I+���v�x�x�ꕤ�7���F
"�y���?���x+�Iq)��s>Уp��_���!���&6XJ�ZV����N�m�Sr�0J�K-]�]�� �ܯ(g*�������L�*��O$�`ܐ�dO���s�?!/�<��:��Xtז0l��־]Y[ZP=#a�P���l�K����g �ݞ�%�7C."~�[N�">i��2A��m�q�?C2� Q�߂{�H`��Ⱦ�����tѨ�0��V�j��!���C�,���z)�ڙX�_ ��֘�H�-�s�\d�JR#�~+����@)�HC����W*S <���a�9T����3+-Ile���pÍcz<�4ߣ��Ϫ��;��ú< ��,�"�vt �3��Y	A�
&���n&];��
���>���&M��F�"~w�M;~�謎!aÏ��u��JU��z�!���x����0lf�3(� ��y�>
�ӎ�����g��)�MS;h�_�@�FM��H�d��!��^��Ὀ7�D���m����?5��ƨl;�t�owD�A�
о(g� �lρ�P+�u�T��2;먼&�ִ�p��h/S���a�%���￠�=&�1�Y���\�e����#	���(%�fjl�X%zX�~R�g�\��y�*.�{��}�l&GBsYW~x�hn�Y"Lv�Q	s�_���G�ԝ��c�ŭX�^x�S�f�>/6���m�(5'�97�ۏ9}�� ����҇N�dx�Z���U�6c��[���3\����Ǩ�%,��W�-?RU�hԾ��Y2�������_Y=06�"����b��$�<v���pGI�~x3�=��Q�Kgv,�x'	p��ޱ!^��9�WQ��r��r���T�H�95/�"�'*pB$bS�� �;��S%؝�pH���Ř����#�_4�(XyM��*X;ӏZm@G�&*�֕��ZF{��+���S�,����"��}A��[:v���G����Z�j7��f��_!���)���r�������B@(±�D�H�R�$����;0_�����4B�ə���syMm9��h���-R�:b�Wp��j@���-�&�Np-�9�1����7��g�4��t���@D�v��[��#�����dZлN^������#�,�O��Q����Q����ש�fH��6�+��%b�p��ft�f�+n�"��:��#GN��yg��a����P[���bD���&&�#!���.$�iN��w�]8>A�w��Q�wO��%�uլ��j���L����շ89���V�?�����'F�X�\[��S�e��m����������S��� �i)�{�h���
r�b#�ȷ{�J�Be�h�#�`�L�6NW16���.�Ɩƥ@j�4(����#;��@�Ƶi]N�5qSXv�:��7sV��x��Ŏ�/X�G�k�:�]�(�=A�C�iq�����ے7M"��窭���ф�R������+����o$C���\j�����e�֪�h�HM�b�aH�&����"/��5�SI	�>x^ޝ�ш	��! ܥo��LŔ&�V�O���H�T�`~J/�a�����N�9��0F����	�\�Է��;�ŵnJ/���!"��wz�Kb��k��.������>J�G�����2���f���l�Z$�ߓB$W�M觬˞��"Y��(�M/�E�3�W����H������ׁ1 }�[%zZ/��c�I���r��,vW��l�(w#�#�rC���Úԉ&5,d�)�^��Y�謘�Q�NO��gH 4���k�	u��������N�H�Vͫ�L�!eu�����*�F���o\�s-+�O~�H������Q\!�y�d_�{\}ʺQ�-��vk���,��L��M�_Jo٠��^�>��A��_A[ �t��dq3m��&Gԕ�ä����]����,6T�ޛv�Y�_�Љh�`m3��a�꬚����:��N��@؃�Ť�����0l�;�C]�]U��^�	_��Eg�L�b�$$i�x��O�t����_u���~���N"�	������ʓ�̯g��.,
Co��2�Ad����K;+����d�
i����Ϡ�-�ȼm��v+���&u�e�{�P�8��odë\jM>���Wzb�����es2������_3 ����ș�#3G"��4�_���nt�=��_^���G���=��6����R�������,x��:�4,�:���J�»6����M���tN����\Q���>/�.S�	�(����zGv΄���2��P5$A��$+�a�Ŭ�6�D, ����q%(Aó1�⑗p#�G<��Ԉ�Y	��>"�FL�+l�h�ੜ!d��~cP���}b��#h5�#s��)S<ZR�����q!����}�����՜�3 �L�����:�2;j+�y���������o=b8)�qʩ�L���϶ys3�	ഹ��v��A�� "
�,m�m]_&����w�{Ho�}l�b0��$6��n|?���i<*B����1�@���{��6mJ�������6:^�9}j�PLB�$�PA����]���5ǧy��z�^fo�w�Y�qS|/�Zlx�����y<�>�q��d���\�|(2��TXi�<n�۬���H7�T^���¢�-L,���wn$ǒ�`h�J�y���(҄w(��͡�������%���%�����i��#�p��Ǻ�s��S�~��.fE�a���7m(ddx2釉�}@]˝Ko�2Ա�j�ܰ7n:��y�b��E�=I��z�*L.[q�0�2�#9����i}	��ϔ~�F���;�xz������s{?
��E�������_���Zj��8Յ��H���/!�]� *gR�G!�Kb� �I�Y��Ⲵs��5D�s�����IŶ2ŁTyp�#��N$�L��O�>ok1z#�S�'V�PU<��*[�ZPYg��LkWnq�TXo�v��cm�u&4�[a:O�?��}�P�!$�b�z��!ܬ���U���cQ%���5�Uc�4�/Ѷ�oR��]��ey@ ��%���b��h$�[7D;_pJך�?����d	�?��S(�i��Chu�]���$�b��v*������s�t�e���yݍ��{��)��#�y�$���X��¾�)�%dJ���rU�H�U�5�f�L��"�V�zI0�d�FUK!��H�uޯ&O�E��h�K\�;�i�R@���ѫ�0��e�O:�����ЍGk�LozH-�Orl�A��Y������l��,x�DХ����0Qc=48�Z�&�G�g4H9B��|�Zs�$7�.i��}z_��T@��^l:)��. +��5��Q���	c�̕C�"7Ǒ�ؒa�7 ��z<�6�����yQV�7�.p�i�E�!���k-'��!	
���F`�]���Aj%6��Z�3�+��wq>�_h��IN����*�h8�=������.­z�G� ��r�w����s��@����(=�=K�E��"%jl�G�'��AV��+�Z���Xwn����$DP���_o��,�k��p~�B�/$_��#��a�����G���9�n>�7������%��(F#�
Q�jѺ$��؁89.���W��*{2�# ��<	���5%�拦�;���,<,��_�״Kt��c�|���#��'��R�]E�+F�k�ȋ>s|�J��`b�_���xl�tK�i|&h�w��1�f�*���B�S# k�bZ�!r�P?ڧ�ھn)ws���@aF�2
��!�`�!D'g�q*���z/���˱F�!���0Jk͛=�B0�^�[cϊ���P��v!n��9l��`3'2XM�����Jߡ�?;�ٹZ"��1o%�{�8��@�6<�Db5�|5F(�%|I(r}�l�<�6�-�:��H� �Ns>��.�B[��Q0�	��ֲ��>`���+��;&� ����3ɸoUG�v��]��N�Qv�ӗEّw����]�^27Q�$����F&ɲ͵-��u���]�g��r ��Dt������*��e���q�mZ,Dh1�%HM7_��\^���v��/{t~�~b�$�G�2X�MT�oX]Nr�5�O�-VK�΢�H�;��OtY�[�DY���-n��!q�? /���^m ��}�2 u���Q��7��
���n�M����8�9p�
I��ު��Qd�$͜�n�-���!��N	��Ƹ�7- &ކ����=C(����-c�t�4P,�Z��/K23eE���d���q�2U�.�)ĥ��E+)����C�x��z�_�D�RƆbl����s�U͋�C�bJ\~��m�m�9"\c�������`��:\���2Y;��]�7AY�p��Uz��V�I�ш��oor����k8D�##{�]��:���������:4w>asp��[����x`́4�����;�^���;t �����A��;����� cG����P^3���bi6_�]+X֕�ʠK�~�{���cR7Rb�[l(��\�Hk��`X$Ah���;����2_!�z5��a�Ye���(u���.�G��P��п����3$�`�H8�3ުcu�������#��o��`��3<Z�P��^S�B�|p��[n�iiRaU� �ǻR�?�\�?N�4������@)umqz��m�.ea��fW�&b/.��
�]1��>�2'֎Z�q�*��X����s�0 <��Y�Ni�s��h��}�ɻT?�n����3v���ɡ�W� ��	���6����lz�Eեtm�U�G�t���,�4�.�@�ti��A?�kd����U6E�����m�M$c��_-���{䡌�9^���2�4%2C}�Z����`Y:�����_[ R\h�U$�W�=(CG5>މ�r�^IX�q���ܘS�rx��YC�u���fy�����$wO�-_,��S��9,l-��~�|r����d ���NS�]si��4).����b>�(�0;f�$97�s����:�D�ZɄz?N�}r�� �T��xe=;��4Qb��7L㔛�뻌繿�[qx�a���K�i;����S��~2C�y� 	�W��`+��!�;
!����w�����xIk8�[��aK�l÷�L�#��6R�d���N�i���	M�N�Cy��!|ym���yw-���@�u��a;����_��A"d�{C~���'!��Qcx�"e�� '�U�}�������B�b��ܻ��Zw>w:�l�p��7�d{��z�h�*���ZC�m�qKIb=:y�Q2\łl�$�+��M�4����K#�%b��v�
�;�R:������Z6�Y��*3�4�Ci$%�TC`��F�uD	b�������@�2X&8��*�fO���'T�z���ǈ鹍vj�q���]1�n�􊼾�~���]���t�W-m���ڀ#���`�k�RW]�)���1�B�xU$��)ŭ�F}��*k��r���20L�J���^���������AR��Ir�h2q*��u��*a��૵K��IV-�;�gY��_w�~��P��i!�cj�|o'O:.�#�#A���Թo-��D�R�π@�؄�	�lq���/��\�=�ך��eit���lOAF��w;
��:���q�b�ଦ|���]K�}�g}��F�s�{l7���c�urΕg��w,��<�G1FdZjz��Z-?�2���I#�csf�K�H�#��p'1���,��� ��V�hP,�Mf�����E�?��Pz�,��p&��O1�#���V��.z�`�T=6?:�cq�ٴ��ڼ�͠05�r�
w99�w
Y�7�0�k��u�DNJf�p�'���q���R��z�Bo<�34")�v�Kk$M�+���˱�R(��ܙ�9!�aԊ���T���P�u����X���� ���:��2Y�ӴŮ<��*��);�ڑܹ7����>��7��Lk�Bn�d����6J���l�0������G)��.o�
��X��E��ٮl1�]�w~���{(�yMzk��@����/�I���)�-]��*�n��Z�bM8u�&�����4\��6//3��ʓ�}@c;�Y�����zZ*-FR[l�#(�T�������ݓp� ��{��W������Y��KV��J|�b��$(�u#ͱ8�U2p][�D�e#�D%F�L����ݺ8�n��W������P����	��[-�eO6$�#�
E��qO�:�yC��T_�k�p�r�^#��QH抝���`5�d5����.�i[V��M>�+=F7o�V�<-�%�����3$d. Z?M�O�P��*y��.�1�UW:kE�[g������=�?_
�39���T;��[��ɷ�e�-�d��E�ED�9�Шm
�E�!GU�`�S�)pJ�咜s)��=`��	��w��a9Ч��{�?#��ȔhzE[a���s����tlE�'���$���+�U��/S���KP��Ct��)�'��ݾK��@T�&�
&W���'�!�''~R})��wN�`�U��>Thh��g�lZ��;��(���+�њ ��r����S����D��I�پ=�'G:��\����2 0�O�BI+XD� �o�o�2�"&�ߞ�[L|��]:�[h���������Zw���l� FEX~�h�Ț��[jͻ�I�l�k����J/�k���E�|���Iܸ��J˱��z��i�D����3i�6.L�G.;;��®����E�ܢ;Dfv{�\��v�~��E���{��9%\L�Ȫ�TSS, ��l��?-w�u&�29��%F�n�O>]��@���t�Ү�y��Ѧ�����g=;ۦܷݵ��{�c)�!�Z�h��c�M!�`Dm���K���^z|�?2~X~��v��'�����x��<�ΓK�H���~�庵����6Y�q�܋�q����>:���<w��j�4q�ky���?K���$S��**o�hR�i� [v���e��x�L;�*�$�IC��j���_�[� ���9Vbڵ�����W~���>����3yDkS���#E���Q4�����|V�����"�9�ʴ%�"�y]Ճ�a1nI{?��3W}˸ �M�oU�W�,������JP��u	~�zk;I��2HF*Ϗ��ч�L��k����bA����y\܉���?���Mv"�-M���~��%�VXN�>����E)hO砿�m�Ӽt
x�8m=g��:�����\� �M"�^����d�)�S����}*�ۆ[�?�ø�����}˪MqRD|���|QrH�t���FJk�o3W��0-9�k��!̷�H\{UG�C�A��{��g��N>1|��,:�#g�4�M_g^}�5g�X�F\o�Pf�2�F�>��{p4B�됑Y���	����{����1_�w���B��~D���8]0����ʱ<�1T@���ꂼl�ĠHB�@q�#yE�Ǯ���m�.��>mo}��uJ���kj�۱D��Tg��Þ�r���H|��y�p,�Ubw�7���3%I1�Ղ�y-�)E��#/ ��$��1�/����{�-K��1����` Ǐ��ޘz�S��M͗U83��6+����.�`5_}GR�!+Ռ��v�N�����]���c!��x���L��I��<l��#[恾����l��FJ�Cğ�y��xVFgfk5���ʌ��P��z�B�)�Qy��=D�+��a��̦c��
�P���n���Wz��Ө	X�4워l`^�ǻ`Zm��Ž>�����a��~|$�`Li{��U4�uV�7���e��>A
�/>�%��Iwu����ג���3nV�����xjF�2�:�][C�ytl���x���l�P�^�JN�t�4 �,��U"��xЯ(g���&�� �G�zmҸ�x��8/�υ|�Z�6��1�o�V�_]{���4�ܳ�,�CY�Yh�؂�+�M#l���|�bv��6Be�|1��Vnz�*�lZ����G�[6Z�,�������>���*`��u׈�m��|i?�/�FYP;�(��H8�U�X�=&���S[WF�3k��z��-�M������� M?�E��m�7�8�'���!*epS��AK�?�Aw_5$��F��9��)ːg֏� c��U��ˑ!S9Ґ�G�M�Ta�F<�V���f�^[�~�j� /�s����+D�lƊ��
��[�\�����~��VdB�!_B��� 2]�x��ܘ�zKc�2N�Vd� � x���7��kGhy�R��Z���x"�X��<���z������ύ�06��"5S�c��$�G1<�ݶ���m�Ǥ�纼�ێ�zn�r*l1���@�/mu��`3]�r��Upn�����c����$H}��1\b>/�� 0�r�r�z����h��#�o��N�е:	�w�u�2����|���V��P-��hF�)2�9*�^*�����цXx.f-�Qr�2����f{y�@e:y#���p4�[��n�O.fl� �Kມ��Ђ�c�F��.耋P�e?�=�0��V�o��'j��3���.�٢�����J+YtKŷ4RbVD����+@е�1�ă?^����-�HIx(�(�hLj���������ұ{w.;���O�&Pp�ۖ�� wq�
�����Ä@���$���)B����A>/�e�sI�8��:��T��:�Q��W�t^t@H++��|+��!�=G���P�@��NZ%�
4���ԗ���F5q�C-ٺQ��w�����5���{�X�y?U�Ǳ�z��.ٮX����`�&�qc'�P�b���1?�7v5��n.�����q�'/yے�t��zA��B��Ni����x�M����xMv?)�S;�Յ�9���w��{�u=ej%=��G���R.��l4���~��D	�xh�ڧ3p0ϱ�~�"b/�5���X�P5B��$,�e5��1�ϳmG���~�0������[��%�_�r��"���Ȁ"vD'W�5(,{L=���G�Ƞ`-���&�_H�5��9]�}�Of,	�XWe������p�?8qw����@��~T;F�S��/E���E�a0N.IHă7��b6垑U���#C�H��[����Z��(w����m�p����[B�vw\��y���F���7_8�:+�zx��������@�ʧ\�ҽ5��VF)|�@��+�k�)~�q�=%ދMw���������}�P�<s�Ȼ�v��l^	�Z���2^S,�2D��V>�6�[<�u�#\�k�৑@]Xo�"��n|�.D�ia:��D'�B����]��Y��ڵ�7�<a�Jn���H�u�h��9���k�����z_Z-D���U�V,���#S	�D��`W�� `�WGg)k�ȉ
b�W�!�w��&D�zs���g�9	y���d�Ӳ�	:2�K�㖘�!���q��}N���D���-zIq�/?�8�A�R�������$�
���	�V�V0s�B��4<�oh���{�-��r�������&Mq��Zo'�:�B�D⹋�e	�vS��Ţ����O��/?�>Ծ4�&yat����3pt�4���sU�HO�U����v˿��91���z�����Z�Uy�%���A(������m>e#�IA��o<>�'�-j�;�Ԇ1.�!��V�:�+�j�	��}lF�A0@��s<O,���t��4~d�p�6�92&NX�m����
N�R�
��N)$W6E���b�-�}깫ڥ��B}��+��<�'�%I����zT�e�i�4����<�fL@�77�V�)z��DAD�-.�"Y@7m�V�9�e�#�Wq%�"��͋�n'l��	mJ.�	C%���K��{�M�W�T��}�ŤQ??��󮛄��>�:���xU�Gs�տ� �c�,$jO�a��tu�7�l8@z�qtBң��c�ϊ���#rp�ǁ
{p,>�68.��kN���!e��n�V�Y[Z' ݓ����^S�=�ji~���z�c�L� �o�8����>z���T#��@��Dvp�v7�,��A3L(
a���Ӯ��H�{[��t�T|�Fã�shn�e�9E��D {r�m9� �:Nl��!����V�j�h��8�����-e�q��#m�j�W�\G�)�nj
��G?n֓�po�1�灩��R�{�1:K���U/��~-��*&��NU+��5u�.�4���+�%���N����Ӊ�l�}���i/R��5��PHz�i$2|�?81�F��w�d�f��;�$�n���� �j�����$K*I�T��̆�k4+a�����S�A���p<.��`�i�����u����&��Qz�F�B-V�C8n	`2�+�C�$�B�ǅ����q��&�7uO�~-�

d�?t\���Π@Uך�% :.����C�R���oVcK�z�����W�?�a�(�m�<���~�s{mv�יG)z�@�(J)��X	<@�z7נG=�b��O��c1y#�v ��r�lUR�Q�<�תF�%��(+#H��! ���d|{4�"3���L�����q�������"bb��Lb}Wn-X�#�\��F��󎑎s��Gx?Z2�P]�pn���d�2�\hO�1~��SÑ�vN��ň��\2ܷC��)��94{��ʨ�a��Y��D^cg�l������H.7(0��(�]���^J�[TO�����t(���PM�el�B6��F����:0A����UX��B_���Dw��m�B���|x�&Ա �y�@j�쩜�,t�Uw�dS�����e!P��O�.���Ǔ��b��Ì�#?�xD��}�&j��a���&�u�+��Z��Y}��r������u�v�8ض�t	���<���A����w�\���RQ!wi־��'��-�:Q$gx�T��Xv{���<ly(Rј��ր�����6��"�Ǩ��L=�b�����}e��{$DP���f�(�5���5��&5r���V6�a��u`��d�ĵ���}��G�rr��c�Hi/�=�8~��ɳaIUE��� '�����̼�N���ׯCgl�L��b�	9�B �شj���|��˝	2/EH�q/8��ᶮc�kl�T����).�eQ7��4������熞��2p"��"5�lZ�c5�0��6g�]��2d��"������J���pÒX5FTJ^u�8����d��A�����w9�lnTE��e�,�JmX���J��F	�) �͂&=� O�M\�P/4�{mi	3�����zZ�}��׫��`�s���O�P�Cմ�s쮁GuV��d��:��'E��M����l}o�`[QMCݛ@ ��}q� �.�N�,�1�����y��>�/��e߰��$`�0���`;�S��|��I��Ǜ&h���7�ͽV^�+�H-q����&�9\��JB��w��v{�#%��C��_�d���u��:ѷ
�Y������n��`p�~skb���T�q��Wt���y��ԷinXI	�%b��>C:�&�/�)	�.S9�6e� �����=l�������ZO���N��0#�}�#���2 �,gN �"5��B,S��5�OmY�3-A��$,�Fi�o6�d�9u��tQ�/M���k���	�4���\}��;ŇwG?)��%nF�0��I�P���3�����{ �ч��X��XW�1sr�IW�Q���<��/�<l���QY0����-��ܹ� �Α�B�B�F��ޘ������Ϫw�M�q7���Tb��m����t���X�ۀM ~��q*�r�t���z�=c3��b�� ���=��T�t�0�0� JKv��ekV�mա��yi�º/A��"1i 3���S����*j��d`����pp=��HT�K�Ǉ�ÕT9�nn��f�_ӥ�EV���1�o�3�G���pZD��ʆq��\�p�0�RDA��D���/�aZ��* ��Z��H0\~xu��k��,`��Q�
��|>��|���`1�A�*��D_����P�4�P�?q���3�bs�AAj�M�؟��,��&*�������L�.��WP1n?�}�!��6���i1;�=���RЋL�]�4��>��R��0��m�,>s�.O��\��[\�����2�>���w���G�A���T���<rڴ�POV�=�V��"�K�~ު�bj�6l�\�bt�l��v��a��Tz�̖P�a��T:�]�w|���:�*U�ߩ'(uJ�s��h�1C2w���%3��/��b�lm����0�&N��tȱ��Uǹuj�,����D�o����14l|��S��2��K1�I6�0�Yn��a���y&d��5�!D͈R�k���p;�$�H�������4ЂU �����[a��#��N�t��5vw��	�����:�p	��Y��ʴ��~�v�*z�G5ɘ]��y��>���
�J���<�C�q(�x��t��3\ɝ��Ju�*��8V�᷉�pkV�YM;O�w���|ޔ���+f��h?�u�jc��+)���G"���N/��MKY����=eT�|��s���uϚĽR�fOv���Q8SIE�W]W��S�:W�"�/F�Vx���{@��,m3|�$�}�����5~,�U%C\4d�E�H��|!�.�:�q|�q?�ϻkφa���� ��D4��?b��
���U�]Y)D�]+�ս{�,Q{(�����ނMP�u|�d�l��`@��3�AF�/  �/���8�9��IA�l����o'dY@�kA�{���iSM�t̿
��A���a�z�.��NV����G�P�����7ڞb����~��ż����n�]z�-�ad��ʕ�ٹHM��$i(<��#�)|saiJ�v�˧��+q8�C���
H�)�����G���'!��+E{M�eZ�"OG
'����XO-�C�CUN9/���[�J]d �<�4��kI�=��|zG6�E��A�)����5I�갼��4@�7�O:nAK~���x��oZrb_CL��Oܙ[�kcB����H����P�ߴ>�6�.�f�ʣ�l��@&�)iy��a-s�ͨ�
O���]��3@�kO��8(����j{�Ȱ�!�ǻ�ϒ��U|��\�,�������ޖ�ߵP�]t��^c�H�\����O��'g4�F�;�Y�sR�b+�x�ߤ.��`���LYb7�?1:�¼reu��Y�_[�:<Ý���b �M6,��=�^�E�"n�К�s��Σ�,�9�e��X�SY`BCS�K��#;�p�b��+�=si,���ןc�r'b�0�b
�����! ��̱� t	��+�����)k�ݩ��i��Җվr��hp�N���nh,O�t�j�_���w��+H�������Y��a�h+�in�+nե[���F8U�8�M��Ks�Na`*��N�޾n�v��<Qʹ��OwC�XT��#7����*B�;
#��M����d�L�IJ���~wO;{�HT�n�Zik���(,���I[�,��$VԞ���K;A�� h�亳QD��	LGc�^&�e9�x��ߔDp���[k�*T�@�Ѫ�W%�ʛp��M�6� Cj6�r�*ӿ=�E�n<�\�(W���"{�������c~�AW�8LW*4X�$�R	��K�Da�F�����������Jqw�o�Cc��o�n�^"Ws��4�1�͘�h�����u�����J�_�ⲝ��B�q(��k�~���9��4s2��u
�<�q��#��E�/��-J��3�v����2�=k���&�T���On�p���^��J;\��>�wh��]��ҝ�_;ƅ����O��X���֟����S�;$�
	LS�ڸZZs��/��K4X�������D{�D�e5>ڼ�PbW��E#��O�4��xXv����O�4�u�D�8+|��T>٬��j�A}�P뚉�`��~�>�k�b]����@�~����}�;�-Vۛ��ZN���$�n&��Nj�ԯ �Z�K�T��w��nD�2$�B��D�C���0nPg~
�d6�"ouF���%c�U�L�Ed�L����fj�Ɗ�L��(�,��q��SY!�j�w��F��<��1�j�q�О5áH	�ՍLWg�v[])�޳�:�[8_�}�?U�i��|H3cN0vm�(f 2Iie�N��݌��ׯ̽��_���������"'E;�E�Z��K�^�+�SE]�9lŎ"�|T,���AK���!������>�uX0�"j���+�ఎ�Ok#-x�l2�:-)�{