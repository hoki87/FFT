��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ���������)�dqd߻��>߆c������)-�)���q�����������Fvw-��xa��D��=S�3n�M��qb��Fxc�\a�b����,����Ly�,��s�8��O7�Q�����)j�cQ�p+��z����Q h	��e�	dn.�f���¶a�A=^�}��]�~䨇Bܔ�Z�*��<��EVY#������3j7�/� J��'O���\�W�4��n�;��ߦ�;��Þ���B�������+UJ�Hq'�_�W׈�6��S=�^�֡>��.a�K*��;�V7�KM�5�=��Jv�J��*:rUv�Ɠ�� ���U<�3��Yއ���[v�&�,y5Q��&��0���҂g:g Suq<��g\���ŗ?a�5�¡@������LS���.�l�[L�;5�q1lg�fS��F3�d��>0B�o%Tv��d�	�\�C\HG�C��j�mmɁ�
9@?�����7+���wZ�Âg֟-?�9������d��D�Hw�����du6:��q�=j��Wf\忊 h`ѝ��gV/KKmk��N-F��g~�����|��/��W&��C�	�n�K�~}��n�������
���-
idW�Fʕ��-5��
�x��#�©��®G[�[�+vy���P����0�]���^?��!����)�q�۵��<�O���~]%��f���_	���Z ���*L�^,��v�{Y��!;����nD�`�O���!�
k�B�cq"�^�4��G�ɽ��Z.i�@Q)����8h�{{�rZ��|���Aw������T����<Ţ�z+��=8���}�I�%h��SEX�<�2���G�4��1��G5>��a

�)v�vg�(�1fҒL$�cȫ�.-z,Ns9*�G�l��y��(-�Y���\�>K���sv�V�{$���1ŝ������Ͳ�꼀`j��v��oa���폷��M
6dQ���b#��m�/�h(��:�IϮ��Q�|:u޽�'����d�q朁���!�@�*E�fMd���p,�Q%27|pMLg��R�`GGw���{֕�L��y�wN�]U���C���&vz.�ng���h��%>Y9�Kh�cڠ��
�t:��rq-�W:��i�%Ҵ�u���7���%�-���Y�I�͌벵L�р`�x�D+B����~�Q��ޮɷd2�āRњ���`��|��'�{����(��1�[�M� :(�EXZ�f��k*9����A��<�V�y�z^�����|^H�|�Ĺ��9��3½�?`���0����~�5�
�f��7M��<S����_G ���0
A����#�����Ɂ%���^����ƧK[@�H��"YҰ��#�%0t�'�~�>��'f��?��k��&(�����%ڕ�y��E������i?�,��ؤe�W�HM�Ӹ�:d��{�]E���'tmx��0���D�U)��<ϲ�fO�AP���Ƿ�~�߂���c.���닛<i�����:;����8�QC'�.<`L�Y�A�l���Ѳ�Ǹ�([)���=��?b��?����!Zչ����_�+_���C��������N-f}w��MV�X�KQ8K�P���g.$�������"�i���<4^�2���?�:eq�pYO�&j���i�5bE#��+E���1R&���ƶ�n�9�y>?�F���QV�k۞�u�2�J�7�4R8N<�?w�~e�!k�1�b{}�o������8?���nu���(�=�1�^���:O_��]Xl���)Qgaըds�+��8�*�g֢ ��b{|�[��bTRK��˞���V �����:#����j�Ow���������Dg KDT�0�����HX`O��&��>ɖ����$zŎ��6d����i�d3�����(�(����WM8)���EM��D]����;�nS�ڎ��g�W�� �^��[��A�{����k��G-�;�*�і��Kj� �6AA^�&푃!S1��� Ӊ���R���D��Ro<R/JJVZ��B߱4%�/w�|It��s�l��\y-g|�ӫ��y�p\�5e��Vs
���0*n���w��K���^����'�����ޢw\����;�q�u�F�L��]����C������1�ĴA�&�]:�v�[0d^����XDױ�f����{�GP����	_�� ��B�V*��<S�l)��I�d4��|7��Z��T⣣�!Ê03ʩ7p-O[Y�e�L(����������B�ǝ�`ܿ^��Ğ�>|����-�P8�J�_��a3R<�ܯ+T�š:�r7U�C���꼒���+��0�$Fj��/��ѼU������s�t�I�˝N�\l��G����8�9�F8y%���H ��2k漊����1�^��kE`���Gɻ���K��y>7ǉpX�ǙFj� �-�v^^�ZNѦ���A�+��5
.�j
�,��®+/�$��^�����t'B`��)j��*��\N�w��C��H��RWN69���5e�.�H>{)^�<+Y���r����R�*��p�����į�m���d��l����*-�=:r�e�٩a���CYMmgU�k�7�*G���Tz�'ɢ�Yɠ	B��O�8h�+LU+U��{�)̢�SL�2L����7��F��UT�7i9���wM*纗������YFA��dɧbE�቉;��r��|���۽�~��Mi~������+,��փ�-:�2��3v�^
*Bh�U��mϞ�-���?���HJ�)�;r����g0� �m
��X3{��#�DچQ��D���lHmL�����_H����O�w��u	C����C�� �������BK9U��\��d04ɞc�!���B�M���Ę�)~fX��q|1��16!���;?�ڸ���=�I.G�C����O\:�Q�ⶍWQ1��4xlY5�[��Z-l�=!�qB�����/;�Ҁ:�L�|�ȢP�8�K�̛�F���ڕ�։E!��X�t�����ku����7�2b�i}~�g�QG��w��ÄN�����a��@����n��G�����~�z0���}ou�5S�u	�]Co��.�y�y�����+$8�k6�}�n+��S�p�e�ɩ�?�E?Q�Q�K��Os�ai�� �'1{Å�x>x*�)��H�M�Ӽ�K'�������H�&��S��6��b�(C����).-��c�h]l!þ>�
}܊��߉��_]&t�y��w�a�A�?���	@��g�,�o8y�h��+�,h{OM!g��?����T�i�6[tZ��{@o/l��Tr�[���Ô �+DV)�<�� �Z��xO,�)$�w�As�#(�'��hs��s�^#F�8.o�]�8��B���%5ΒM5_ѳ���=A�WF�2$&�F3��	�y���ҽ��hBu�Y�XD(x�hrEf�Z�.�oR� �uHN�(�\���е��>�~>�}�Yqق��"L�9U-�	�r�u����W�wTS���Ԧ��\�I�E8�F��7upl�y��Xڗ"��� m���v@I�=E:�<���jk(�aѝ�Y+���B��smM/��ᡸ!�E=�c"�)ސ$^Z�4���>'V�E���!��o(��6�L5��̀��l��)�Di�eæ�AJ�??��"]��kz�>�h8^��ߥ՛DK�M~�{et<R|��|��i�C}�������<{��]ｈ���0�J�LK|�p���,Z�TV|�a@��	�S6 ���=���}U��.E��z2��R���h~`d���{�ģ��u?��?_[���}~E���pW�*[�r�=N�c�(�,>frќ�A!O��/��s�I��ϔeb�l�#$y�����atb΀��B�`6�z5(�]E�o�\A�8�}2��o����<#���Ƞ����@|1+��1Z�){������g/�e�y	�mܑ�<:��jJ�]�S��Ť��>�ۓS&�c��f�#W*��S*����^z����:�?�k�SMa�(���\�<�Ŏl❕���`�J�]��lKJiN�~���d���Q�["K�k#�>�5M�w�H�/qY�Tz��U�o���
ؽ��Fe�`��w�i]�2$R��<T����C�pw(�i��C�.1}���%M��P& {���B	(u+���{M�c��	8	����\�M�Kho�C���pǃ�	�|�� N��'R��a<f}~�6�P�;�-��~��bnjÉ:���'i2)��ַ,^�����J�sb����s�^;��!@D��ۿ�@/���h*/|���A+45�_K �5�ppv� c��Ԟ�5[V<6#m;^��,�@?���n~�( ��2&� i$�qf~	R~~_��bt{_��<�
P�B��@"C�-@GUB±m֐k_:
���å�����*esL�p���*aR����d"4x�3�ޢ����z�_|�yѩ��;���u�y����w��3a�~z��eZ���y�G����߼���.m����C��<MK�L��iL��T�z����b��R���B��֏�u�|AFf2���s��Q*����0Yru*�����a�,����_�+N�r�%��u1��������q�|��Y") 
�ܝC�q�a��"y~.n���d�� �傭]-E0B]![M����7f'��b�.�����;<n��ÿ�y�
h�$[�Սΐ	l��E���d���4��:�m7+nt�f��V�_U���b+d1*���@���i�ɡٔM7H��u�B�D�͔��9g�5"ң��%�����;=糓'�����Ǚ����A�י�k�O �o���/q9%��v�/��Uzxy5K(�]�����2qڃ����[�i��
%w{Yw�Ji� sw�O�#=�������Ql�Ge�rv�4�8$0l����O�+�8S���J2���o5cÝ��2֋�גr���]A�]��.U���dwU�Gxo&�#��8`σ�b(��J������a�~�F��Ǟ�O�$��7܌Ǝ��|�^����t����"�Da7>rc����+ר��:WBA�Ժ,j���7���ؕE�q��|_�~;��׿�pq8��D�_3�6�2��x�k#���b��X�[�~hHl�" W����K��P�Ep�Q�W#t����ϗ�����<aJsPe�|�jJ��,	�&�n������^;R./O�_�4����o���ųhW8��7'���0U=��H�X�{�8^P�m$<�7��Y�md��/�Y`w��m�J\٪c�C����"C%*P���ī���B���݅�B���4�Cw��z��o���W�i�݇�ںp�@��F��>��7EBx�`~щ�/��>�T����3���s�r��{��N�'md��t^V�2��`��f�ĠĀ������&���"��^��yHǕ��O@{�yLS�Ց�h{lX>E"��G�*o�4l/��GA��_J����lE��1��*��Bs ꪭ�K�(���[Y1&$CI��d���9����h�w�O
||<5xj�|�;�a����֜ś\��^6�%�>�v�XD�^1������Ӝ(�Ti]�<�#k#y�6����o����1ڼh?�ōV�U/�(��l�����6GK&b鴮�"�O��/�#��;����}���v��W��8��m��\B3���/뒊m[+~F̬2kZFJ�݃]F�����n� �4a���\���~�����Y:G��z~+<V��NI�6�v��Q��\yG���J���y�W������<۩��)݃�Lv���_ע1�*1l�N!]�'GBwG]���}~��¦a���_�QGh��I��+�"�t���M���8����KM3Yc#���Ii�v��T~z�4&�R��8�f/���`#�B�"�6�B+�̣�nҷ��Q�Ld��3��[m��������4�3�j���v��<*����4!�I<;�} ��fܳ��}�a��f��1�3���8]�a��;pE/���1yB�JY�x��t�Ÿ�{�cRa��[t/@�%��#����`�z���¿��	d�&{Fw���V���Yr�����"(��us�'B;h�}���EF���H���p'�U�����!���80]\�y�7�ਨQ/> �AM��[� �&�Kiyp0}[��θ�2�� D��\NP>A����}\lŻ/�C�$S����%��Vc�~���jɬ{����8��.��ao8	b@ާ��AOZt�Ńg��ʿާ�U<1�A.�5�aq��c@Ç�k[���9#�� ��r&���m�A��y�$���x_8K�G��h�ܨ�^����Y��]~��!-z�Vc�oe���'q�,o��f��4�G���T��F�,��n�p-��z�k~��T�ɳ 5�k��ز�sp�g�s�-Is�6��N����3���~���׍�L(ֽ�E��m�w����]T�TW-|�߼��td�ԧV��;�@g=���fْ��o�`�����Ѐ�\��1��-xB���șĮ�P�D#�Z����;
z�>79��(ޡk[�����{���m�P���q21h_���٦sz��C5g�)^X������}��C�D@�'��4��V�Җn��XqXX��2��5�N����XgzTƑ�$yht�E�_�4�Y5�<��b���4���c?4q��ޚпZ�+�P6�ЍO��^�d-F^��)��I�(ؒ�2�b��Ed+��2m?�R���<�%��E%�t��+��FͦvVh��A�Lz��|7��!3U���޲{ސ��-��W�|5^p6�߅�o(X�"����MW�{�,[D�#oN���B�4I�ǨQ���LP�L�7/I����%�?�j�ض��s	Ks�C��];�w�NN-�&y��^�<�;� ���^b�Ć�C�yHX?�����y�����SU�8�$Eӣ�6�Ajn����	ڬ�ƒ�ͅ���q�Ȏ&�+��w;%�_�l�3�-]�1�aS�n��`5�-4C^�ԫ�ص��P�i�{js(c ��9�	&T%�m���"}�M�^UBChŁ��A�wh�FS���������GS\q�Ծt%n��/|�]��ʾ�f=U��y�U�i^����`ݶF�X�^L��c,3J�[Jr�F��u%	!%�80S=B��MX���?����y\F�f�b���]�r������o�uV�'ĿYr2��k�~�=r�|��v2��z��p��G��P���B�-,�ig�m�K�e�0��?�oM��=|�:�@0���*���ֵ��Pwt�O�����Of�����R��,"EȜ���
��`�/��g�'��7�xCX�J�2���{0|�g�i��KFJw��vl��\RW�����kW2db)#=��P����	��d�]ǫ0����r\׻�r��ם^tѱR����zNi�.dk�s�F����g�O�:F@8kHi�ś�ߌ���b����B��//o�R�
'^���3�����=�,�2�%�G�m�_0�z^g�Q�dx)x��tӛ�g7�'�QvG�=�����<Jó���Vh�<T�<��׵�������y����s+�Zŵ0|�$�he�>�F��y�y�P��I-c�q\Ue�n����H����9>`�j?�P�\���uݏ� hX��+�Y|B�0!����8��.mCZ��
'��0�d����̄��Ɣ�B�Y<G�(z�+P��&�#�) ���b����D�:#�M�*R�vhrU>u̐�q7*�88L��ŷSu!1�5f��"u�� /b�U.��(
��f�� �[�����!�H4���"� G��;����/`��A�?���Z��)�܉kے>{��u��O�k�[f�wW� �3� 
�~�2�%(2[m�y��Y���U1�8��H�XRP@7)-� g4�>�\m�,�Nx�oF�D>Z��S���1��d@� ���c6?+~���K��g�I�����\��ξ���JD�/m�UH{�s�N=6���P3�D;\�A��d8��X�Щf��8ԩ�~@���k��Fsdh^mD��϶욃e�ؾu��ǅ@�mC�
�N�ʩ��N��V���\�$��D`�3�WV��RIy�C�4�i��Vy"%�?�͓JU`{�Dx0u��Yu�ݭ䷳�7R�����xЋB�M(�`<��Y�5ɂ,{i��讠:y�bt�7��Bac
ퟩ��OB��pdy��A��u7��&�,l���Sn[PѼ7���5@�=Ɏ��d�\���)����:H���:�쌊}�8�:����H+z�Cm��;�@*���lq�<��G�� 5��_Zd����'xz�s�ׄ�䌸�1���$�3��׮�.>��k�^g��9�o�M!�Tu���M���m[�Ie����BNZ�$��0λ�������O�ތ86��:5ɗ�o��At���`�c*�տ>�H����U8�9�A�K�"�c�Q$_e�\Q�	�xb&Pl���Iy5���������Mw�㞬�9�q_�0m��q�h.M����#��H��^����iA)~{�M�-p���j"!:���EW�)��'�Nv������1��AL?y�8�'�#�V5�8b�T�%�����E�j�&�x�>sН��ۨ�1,�,�����A�;V�+2��Ĉ����[p�-#�2� �%Ş�\�V4���q���˞�Wn8�"��$���Iwy�\���?�=�܏�Ƿ"��	ӑxp�ie�t�0/��9Y�˄<����넅X��i=9���bU�k�*���kc
^:�F�:_�:�?����P�@h��y$�t���$�-��+��cvA�.��KJ���uR�l�gP�
88*�o�_��Oy�i ���w�̦���%��=�<P��KD����\_��6JU[�_��]=g>���~G =t��`i�ôA�T�3�@�����p���~�������;�Z��h?q�g�����������Y��:�U��1�Uo#�F�5V=XY��̃:4���7�w�ꑗp�Aߍ�z�o)1�C��B���Im��7/����WX5}� o��u���X�2�Y�4�#�Ig4��>K�?<���t=�[��6�79E�er_m`7t���,�4G�l7d8�����[S!�XtH�/�Dq�@Y|��b����Z3�G�hNj>:�/q,þ���V-C�s�V���?�u�U)P��f�=�4T{�|	B26��n�٨�K�Zt����*+�;�
����煶��z��}�Q%��'�tQ�S/2���\}��a`����>WZ�zQ�B�`���ύ����_:ܞ�}'Ü!L8���L�P�*��*�+����%c�*���P��尵�1+����?�5sb�U|^�8�<U�a�'��E��-SM���w���}�cL��˅�~G
ٖu��*N�b�y��!y:�+�ɗ��VC��G��>�ep��@���ā����'�������E���ϙ�멄�s#h\���� �I��;Y~`a)�6����-�9
,�R)p*l�}kl�ö�D1 5}J�QB&U�`
��@���Zl���Sz�@���J�Iܮx�_�P��<�ʎ�<4��P;Sjy����?�&��7n�4�3S�\������C�C3�\���\荾Yr���Jl���7z�[:�S!���٦���9�oD������ P};�s�A/��ԞJ���OV�T�T�!�/��\=Oٖ�H܎0�\۶Ϫ��5���|��5�
l����;��{�U���*�R �q�T0�0-0"Qm�f�%q�ژ���+e�6{5��k�w�ơY9},���| �ѷ�c�"MV鉗㏊l��pЄ������S4�c2^��)u�E�vՓp��Cx'u{-�V�uK�������� �I��},rE��0�i�>��c�������B,�6j��W#Y�b\C����:������ڮ�i������7ޤؤ�9Oő����tU�T��KϿܗ�����5�"+>��f�1Ty���\q��|Ǘ�R5��8)�Q;�G�~9|�ؒ�m�!4�䥅�*�ЅϮ�U�8�cd��e�E���� ֤��pQ���e�n�����6���S�.~���b��I�l�'�:��=�\�A�#�u8[�Qv�p��zaH��ʻ�y"��!8G������,9��zzp3�c��~.8DwڅF��i�au5�H���}�;*�"�О����Jt����n�,?�%��:�jce:.٠jюu�K�2�r	��	q��e���H�)ģ�ꊡp�
�����G��Z:-Ӱl��Qs{��YD��y�|G��o��c��+�ݲ~�������!��w��jda���з4���F:帻i�yv.���6%�'�V*Rtm�;�B�2&b�2.	�?ǡ?�t=<�E���"�\ʾ���P0 -��_!	�*U݀���<~�����Y�Yl<�#�3 ���~e���^ِ�˭E��crܖQ;/E�+l�1�<�ExnV=�W���lR��&b��8zץt��#��9����ÓM�0HB�]�q~����L^�=(�-J&!���{�?G@�%<t�=���!h���b�餬0Д��a�������|=���Ǳa��d� ��U�iæ����&R:k��� 1{JAC�Z��R� US��7����jB���gXw7��u��;+���F��#̡I��g���G��"�F9ݗ|X"�c՞$��Y�����\�SxC���,o����]�>�k#�����Qى��)1��5Qb(����ID0��N�9���*q�aA�o�WQi��G%���N�9�=]EY����j-�rǍ��|��<2�8ܢf�m��ZiL��護�!!�aIcW	���ʋҲ� �؇�s� 7��2���d�<�9���)8.F::�Э� ���u�p��1��������]�%�rt��hU��ޤe�>d�g�3��.�!}�%������}�ߊ�� �%�n{���L%;܂���hx�ԋ�9#{=L�$G��V�w�Y̨�>N.��L�5(9���+�H$ɀ$i�t� 2��"��X��>w�2�RW�l̹����T��>n�go�ק�u��u�_��}d$�3�hs?�U��:����x/�u��@�_K�����[����W�[V�̫8�"��b~�w(�}��~,�h|�.�/��G����+?���54�>DV1h��2�q�Me�J�ӥ���1�Ss�R=,�:A��h���-�h�
�c�]��Ǿ��}D�C�w�2��w�<���є�~ㅦ��
3���#�v�D���%�)�&ԧ>Ɩwz���0?�s�0��{=���G"㙤�h��C�u���3�bv螂��y=�j]��Aq]��I:�$�u�E4���3���C�&h����"��, ��a^��*QqUܻռP�L�1j��ga��-	ŅGb[�p�xH�;��+>�|K����w��n��0�i��yu�`97zv��/~��g�0yh~Dd#
���nԡo�Ygw.���$��_"b��"�!�\_H
D֌j�_% c�X<l͉څy�{V���~t:e�,�p�O2
e�ȦT�p��{��Ul1`U\� )�&�r��2��{��K�e�K�u̺K���
%��~�vr-U��@Ps��*�l�[�!���4��&���R�-�2cY�`:튮b�ی��Xf��n ��yɉ�]�oJ�?�1!q�c��/���A)ɜu���+�W�'K�<��@y���$&�s�<O�.o�U�@%��|�����u�ܔ&8EW�pVחMO�K��RG��
D-�<�䀃�Q�,���Ҋ��
�:�FJ��Y�y7u3�:Β7$�,[O������ic���[B��Z`=���S~~Jު[*c8 A�i(��5�ӁS9�F~~j���*.���CƁcn�
��
��{�W�o�pڊ�h�1��AP�ݟ��GKi�)+�����>0�Ɯ�. m� @��+���uF|���?C~���M1��~P�{gX��e	�a�cF3�n2x��ѝ��D�P�����"��6>�t�%��H�E�/�[�7$K���yޜL�L�ǎ�#���7����Y��B���6e��V�S��j�;P2�$�$����z����9|Cr��PPhY��&i�|eڳ���R/�������@�t3��.A��'�>���!_�������"��hb�˾ۗ> V����q~<�)CRU�W�"�˾4re8p�v;�k����Ka��
ZR�O@ƈ{�ܿ@L�����g�KrwK�&Q�>;���\����IQF���p��<dD\� 	���O�8���q_l�Q�X6���ؖ�eL^డ5�G�wlh����b���?k+ zƔ*&�����KN����X@�o��D��jЫ��A~;gP���-�P�a~��� Q�F{����;��Vd&L�:��G�&SUbJ"����+�Y�� 9�8S}9|ء�p~����0���
��$�ɽGL��V����'BL�9��D���3�"K^��s]�`�w�E�*f��DO��d�3,e����~�;ǩ�Ku�z��V�l������P��4�����x���m&3�l��6�#�Y�D�u��Ѓgĳ3p+�8��@�4R��`:տ��xOi"l��U�����:�UB�l{K�e�3���7�5�
�tZg�����yc���K�*S�<�\��ٔ�53��R �)�?p|l.
|��5��eȟ;�<)䩲(�f�ViD�i�-pl|� ��0[�zB�ۆ�#���o�
ƶ���̠�E�䲉��˹����:����Q��>�z̔{V�*�|7]���N�"=�}�y�ʹ,Qְ%�I�c-���Nk��@�hp�	޵���e0]�I�!�&��~`�
7�6�����)a��Toe�\:K�ֹ���?c�Oi�Vf�;�;��g�S��3T�LWz菍��gd<�y�8Rd�{q[�~IĒ�ź��k�g���ں-ce��s��-��;3�O�Mf�\�n;�(���+��j����^{u�7��h�K��T�*P5��P:!�
�b����%��",e�����Ľ��c������l\�f�Ŭ5#�6�`�ܿ|L�\L���$'�m����qGv%��n���g�{�螻uof�������Vf)b������*~O�iS�G@l��PI���GJ�0�Av��P��=�=��:]�gH��,u}���5Ap^v@���}  gQ޽Qrx/.K �T����AyUEW&y��鍹~-/~�FD�ϸ@��:�\�
�I�F*��
�~]�Z2En^/_����+ɏ�kL�^bs+3�n�*W2T8�-�;���'�l	��ur�*��G�i��H��`,M�s޶vkcіt���^[D�A���zݵ^k��*�. 1A��K�#ol�xV�rt#v���æ�UH��/�$�s e���Q�dHtW�z�#:v���F����{7����}�����&O)��9��e%4v&Z�d)�`MY"��:L#z����8����c����Ds>k�Fyk^d�O�}��B̸��N ����Z�6���F4�U��A�u�����RŧԗP�ɕ_qt�--�6�@X�.�;�����E��!n���ZwOg�r�u&N],���� H����0#��!܁�]iz�b�d����@��𐫿_{��y�M�
�L[R�,���n�B���d������l#��q3��Эa��v���i������UU
̌W��.�q�E|�}�]�����l�2��!"������IU�T�1���@�io�w�d�z�t��/�f�Z�ϭ����a�Ww��jB9��m�R����V�֥)_V��ޓz[I�x	�X��Q�/���C������U�\b�O�׼-�
t��?��Uʢ�����A�_�6�@�
r��(� U�0/[`��!x�$L�-�N*����+������ы잢��Aw�3��m�.׋S�G�x���oh|ԫo�ʩ��iKl�L�L�Y���<��[XI���fر�)�aK�<��`u\!0/�E^{4�4����(��`��f� ��'?ȥ�����XM�n<�l�̵�@�����Q����6ؕX(�G.��>Hp���R)&���X>W������p�ѧ���(YՆ��}S�O[�*9^�v�<��3�Wʚ 0�i�x�[�)��,`��O���j�Vk���#�06.�ˀ�%p����~,b����@�k����d(Ѻ�ዓ:�0�Iwv4��`��H�s@!�+Vj���O����[#�eh���l�n�^� Yi*3Y��U;E�l�-��	Y�GpG�	

�c�%
+�u��x�AŹa#��e0���,d�����/���I�S��<�:�b�)��Iy��/�Hn>Ar������}���(*��s��Fx^h4I��f�MUb�<�8�e���m낿��	�Þ'�F�!�sa���^)��,6�=Ÿxoʜ�j��W���U� �$�o1�p�J&�e^�h���`��}�!���61�j��:���le,w5ڜ�:و��^ܱ���Em_^�^�x垭��dg��]8N����ĥ�.	�=���[f�F�H���Pf�Ǫ������%��< 
�_�T��������YսAƂ��a����So��K�Rq��J��G�����_ԟ���9~�y���#`�j]��.��:Y�h�l�d�k�Ml2J�Z��Eۭ>�m�7-���R�m���n �1)��o��?3@�VI)'�u{Ez���2th��^��M��S�PdMiT�1[dJ��Gg-���[����lm��d�=̀dCA>̙�.�����H�ai��&>��q�X��h�՞�����7{�4!�x[�밃Tm��>*��a�<|�L�9W��@5j+�YJ�E�X��7$�l�������1m�r�J���OҢ"��&��\_���S䂢W	����1�_���e�[r
w��(���g<.쩪�������6'b;�Ů�s���S�d�^I<W���j��e�y�dZ����,��f�`�Z�IL�͊��Z��0	����8����פt����y��G�,�H���z�W�Q��U?��Z�b,x��d��̒_&Y{*�/��,i�a�.-�o�Ӏ��^}�]H����
�3m�����q�{���*a��r��0�5����Ⱦ���W+���)S��MY�G��<��u�?!P����.��+��r���p�Tb�Jc�.�-re�@u.�������1�]�����HC�9̉�`�J(X�a)6"�f`��flߛ�Z{�p-�@�Y��a������
�(��*�.��tD��AUtSO�o懓H2����Iu*~|����!!g�Y�e�,��p���X ���n�Č�3���|0[~��*apN{ɤ�j�Q�3���4KO���O�&<�nYN_8e�)��;(P�$x\���#�d�G�B��o��:a�u��c��6hc�r�=l�9���d��׫�5 $�X�P��8�3��!�1?��W��o����+�naT�Z��k'nP!��?ے�b �?7ӄP�u�0w_��~�h���i��3l�_�m���M�0M�_cƬ�f�"���Nl�o����b�:���ÂF�w����L\��sGR�"�� ᙠ�'�gQ_��d���ګ,��J	��k�t^i#��Jx�JgWFQ�=;[���(��,�41�����|׀m������B���Ǩ�����iZ��?��n�s>�I�W�M|$p��Uz3 |�.�/M��SQEl����i����ι9>q���������Kk� ���+���C����b�0\���d�/A�ݫ�y�d$��B��� �T;-��o�W��fhynX���q��������U��*�''���al3�@��e�.�=�n�Cc�t#
RFz�h���i>���0=�u��~ "�y��D�K�})�Bg��%3�b��/�4%w։{�L��'w
�oVS1�]̏{���z5\U_d�;���gy+U�7+���;{�=��U��a���д�C:��Pʳ�L񨼞[F��5�"rwi$lS�����Ϡ�G}8��1C�AlɗJ��w�j�ml�IƬ�m�!�4�S���?2B\���x�p}�ʋ`{g�La�"ò����$�
Fj����iY��8�[&���L�U3�	�����Vd˙�[��O�2`�S��=c�����9����[� 0@�*�zA����i�Ѫǭ���rPy��M�T�����Xٱ�r���
�R�s'��#f����q��NY�����]�갸�=����Z����7)�{ݴ'?Y��������ى����o0�3ցR�z���8��*0�S�DbMpp��e�����F�������ˣM�m���m�1O>P�9C�h`6+�JgF�,_���߄�	Z}0�4ܒ�������d�ϕ�!Ab'�l����q�ю<*��<�'ea�n��(~��Ff���� ��nӢ�C��s�eh"�7nN����~ �s�LD�yy���4�j
�_��ϒ��=�L!�4��� �vI��^ˊ��y@��!ﱔ�6�N$˘��.Ħ�?���61T��
�Yq ��s�if��Ħu�*=�do�AX�+�K�ͩt���{Vnܼ۟���I�����f��y����a.��b�����1bR��Ye��!�8p:[�$����:5�.b�����Qr²lu���x�-#�����~����~�k�[����˭��8�2�*%T]�k$��D0|�]m�:Q���\���e:�-��hA`�={����!���k�<���s�� �����r;�60���4��[�^��fw���1�ɿH6�}�k`_��w��&3���6���0�ɽ�*��o�,��۱�c�D�
���Bb��M���դj���u��������?���YE����ҙ%�Sx�-ᶖO��);f�������^)t#�[��9`=�Ej�}�c2���5{�0����V�	$�K��B
�x���G�a@�]w�W�I�k`,7*3S���`���o/���3ПXF���NL�:B*�8��Wo���� �$�4�XKrقsn�R�o��W�:��S����GUF�}���o��i��O,�tyc��(����3Ih�zx�����{��A�Sz݈�������ސ����B�#���U#=3��-�	1�������� �#����u:��H"!ǉ��j��tH�?�}����֌���2�B3N�T�W���P~2�͡����ǖQJ��S$6�����#��Rr�~�֪�(����O3��@(�ɲ�@61��9^@�z���f��y8�����k�����d9�V�$����x� ��ɓ[�W��[ ��	_��M���X��(`!�Ms��y����b'��ݏ5݁�g�)
�%uS`W�=҂�|�CB�����D%-\ߩ
D�q�R�~s-�t�p1�Z��/�?�װh+Ar�3��AA"$�[���D�ЪΝ���s%4���-g�TF,��279V�|�J��W:��gb(��eh�u(���X0_�4಩�I58�%��t�ȿ�vmJU�i���֕�M��`��LZ4��������n��c.���.p�.��}��u�ck*k�M+��`��X��"I�e�+n���m���V�}k�!�ƥa�t���MKz�Y8��SO��(nj��h�<��yz�#Ǫ���_~�[8�V8�}�i n�
eZ�K9�C��5X�3H����� �?DPn_��d�3�=<;}�+��TT�^��Z�B��5�E�:�������c�DU�i_�iy��=��M=��c�fn�:�^���~5a��.Y�$'�|v�z��7C$�����#���7��(nkF�sT"�(PF���U�FyTj���E��e@R�AH��2a��Bo�����N:�Lh]w#���?B@#&gЈ��|��%�G��`ݕו�)C���*9��{P������q��&7L��<I5sOiC�wk>��>��f��;�*˶ l�:���f�RLcʻ���R��\ 2$*lv3|�nY:
<I���� ���͞t���g����e�����#� b�(�XSʳ�#C�?N��$	�n�s:ma�w%��H�{{X���6���I��n* 㺥FT�q웘Fc�|�q�%A����|�{�i5��#�k����a%T�ҥ`�2W�'���x��"G��,;l#��S
�Қ�jL�(�8@R��8� �WzP�Z��Hnd�fÈٰ-�rf�*�@6�ϟ��]X��k+�'��M7<�pe=
��i�nW�.Of"��<���)���&�6�ҋ9����������;Հ�sf���?!a'�P�����d`�C��Z}@��c1ŜGT���x��r��Ѳ�L�hk��,l���a�R٢ILU����ukI��)5!�Rbj��	J�8��O�����_�X\[�C^���g�)ސ�w���<0L�՟?y-
�sM>�1���-)���` tBAQLU�`��X��O�e*�g$ ��y!�ybK�q���:c|-�����G ����a�����W��PBۀ�!�/5�?s�Gk�.1e1��:��U3��Q~T0�ty��a��\Uj©f��S1����������
�����D<������t��>�]\��D�"���󠗠���hjCN�{��͵?�p#�":�K,B�C|����kJ8D�,ґ_�=���PX�$�9��o[F����xuU��w��͹.c[8c7���T�̠�����ǝD�-è�8��L������
A�i�Tp�9�`��nN�=�
�%��¦⏱������1���	Pw6��ܤy,^GN��Ju�]����n���ky�,J�}����bfɰ3�[�����%��L� �����j/������a��i�ֳ��4�p7Mjɿ}5J{.���V�2�zP���"C�&&���������xWDN�8���~�{���d��h�Px��hK��w��[��Q4���8,�m�Ꙛ�k�"N/?9�OK�B����y�~4�-L�/�>g�� R�0>�o���"d��(uτ�Z�,�kg5���?,��������7�	�4Ȗ@)����X��ή}�5n��N��p[��-1]:�p�rJ�{��:��"�=#oRT71��q��WM�5��	�l�$J34_�@f9�X^�%L!��%��U��;AZO��퀉��"�{��*�Wt,uA!��Iv����G�o�7��x:*��ݻ$2-�q��J.EhYVT�P����D��"ـ H-Z<4���<��GM��h��J�+���lFx�:���ix/��8�G��4��&ÒAx�]?CF�?\Js �j!�ک�Z�E��9��@^�ѓ��r+]Ҽfq%a$�.}̐�]\j��P����[�9?�^ȑNT_�eo3��}"���Y�\ �.�N���s @����fV�6�Zb2[�s�f��ˡ�P`9W9M���~���xk�[λ$]���C>�`9/�QK9�s��������&cC��!�@�Vu�ZG��)���]5�K:vo��Kُ��A���-�̎���q�#xn�B(\��� -�{�"�"���B��QF@�4bʬ)�2 ։�Q��B\��W�d�$GLA���<�lW�}�c��x�z�?���D�� V�)������\���V��yZ^Jk$�&	c��#2"�WL���݌��X�_�xe�o!2��7�P���h���YkŞk+����������ދ���s�p�Fӡ��b(�Ǽ(})�p�"X��f*��V���ұ���B7�v5]Nn�������7���<�#�"ΔÓ9W;.C̾�$�z����M#wZg	��ι�8Hs{�	x��"p���=BxT��c��j�.�H�"�w�Vg��,CF&T5�&�2��1��<�D��A2ڛ��8�N��SĴɔ��OpM�(���r���
�
����7!�v�!��W�P��U�\�O�B��mt�g���p�Ŋ���C�!E{�Z�\��bJQ�_�:�<0��>��qq�;2n�A��eT(X��)�=�[�Bp�B*&��i�>��¾��`Ihcqs~r} ��$�t��UE>�nn��-����n&H���7��&���=H|�A�3�آ�
͋�� N���
 �8��x�-�6!/[�9���2�۲m��ۖ������W3^�>�]�4q�eR�hǩjf�i<hӤ�F�Ek�Ena�i�u�]Q�2��jQ���:$�X�ml��0�]+�b�
���S�5fwL��HGc�ջ ���ֿ��Y�{�>��B'��`5��/��B��e��!��`�]�+L%�?(=��?�%z�0/��`�ē�Q7�`��2��Ğ	A�M	���V�n�����%�ԍg��q*�;[�b�:c�M���>�����BN�9��Z���"]��D��a÷����V�4YV��ƃ�'���>��6$��B-��O�]�� �i� *�&%��ߣ�@��MAIӚvzTF� /�<h!��W��V�E8��Ȣ_�2J���*�8�c@��U���v�x��:�+��{*�K4��~�"7�c�� �wK���<�����we�*�@�Ğu�/ͦ�Լ]MQ�2�0 �Ho{�%��K�-���%6�5������u�,�,�2�M����3*)��*q$�}��n�p����~D&k�´�Yj{�����GP��`��^*�C�/�xb���eM(��t��n|���uw��R�~}<�f�&�]�ފx~5�g�T���gd�%�)Ͻt�V��9t�u��j�L��]���k�c!� `ʞ"�-s l�V���^��ꠏH/�#�;�lp��?^�F.����Z�	�@ҍ�"��
=w>]�	�-ŀسϜ��qf�f�鍠���cՖƱ��m��������b�H���t(5����cA�1���'�.�'�Kj�qd�bY�r��V����b)n-��96�J��B��yɭ0NU����]*a���}�ר�ߌ�_�Q�;����ѓ���^�T;�-l�ԛf�� ɽ�6ͩ��Zez��E�Lx�O]N�[��tM�4�=T�f�*9��?�޼�~�]N�$�Nm�����|�^�osC�5x��J�F��m��Ȱ�h�K�I$A����h��,r�d�0;�^�4� �U��xc�l1ը(t���[ˏ2�-%YC	l��\j2�]]� nb<��ڄѢ>���;�.^�7�n��ok�9 n*���8��L{��t:?��9i׵��jӘ����@!������q�p8���r�KS��f�u*�/2 �-{}�B
�Vj_O��o����K�����Ӷ�_ڗ&P��.��!�6F'�A��1*����*�~�	V:[�|��Ү��,Z�t�1���+Ul$|j��`	�3��[�ņ������]���bi	��:v�/����btK0+QNX�Z1�q'hU5���2��g�&��?��������P��Ә꿀�cB�'��� y��<�B�_H�\��]�M���yLujǵV�ӊ(�'q�I�nd-i��K�u��g�?V~�'E<^���,M9���pke�GI%D�N�����5�{���!���r�9qC���يEj�M��a��o��F+�KUY����y3�L�Yyh+��z�-�Ҋ�����ek���4��>�L���
�l}�(q��A�
�$�a����W�|�%�A	�@XK�*�ԥBY��UZ�Tu��s�w�����3�b�8�N&�����2�7eq�[6���D�����{��b���ݹ�%y�n�'=�ssV�����ʈE�
94�<��������$�����L>�c2~ɍ]H�*�9�V���JG,�T���d�̃	Q�mj�?�Ѫ��5I9��=��db��	�i#<�Qԣ��I)~���k[l�T��>��$wUޕȭ�˻V&�&0���6}q�=���;�b��b7'����q|�\�C�������Y�79�}��-���,��j�]i��;To��ƭ7m�\<����{/zP@z�@w���������w4�OX�@>t���� ������r.����}���f���mէH��լ�����e";�D�J�݂@�E��ƿ��^;��m�lN�V״fUy�<;e����D���k���㌣5�K��!.���ٲ��*�ۍ2w�4 �ƮQ� �U�j�K�_]~N#��a֘HV�nJ$ɑ@Y���g|ę��FP�8W��UgAy�x$����y�DCFi!�A��2����q���M֬�V����w�o�kr�~Ԥ���,Ȝ�e@/s�����((Bfbݵ��V�F&n��qU
�Z �U�>Ԩ�(oC8�}(�����&�)����+�Cn=O4%\4���6ȼM쯧����do[�������Ȼ��Ɩ�>J�&g���eq�'������t�8��m%�{%6������+�{�Fz��GYb�dM���=�B������9~�����5ǉ��� ������m��r������_Rc����ū'H�1#��g���k�����*g�r��O�RX���o����Y�I��Cm��Zk��`Xu�%�]�E>�jn#T�����$�ab'wt�j�����=�X	{�d^Ű�*Y�����T���*�Nn��U��W"��Š��^�O	A���@k�w�`�{���!��C��m? � ŖQŔu���0�V{�-1�7b������{�����jhx�iD��V?0��9��*���Czg���n%�������"�W�N����G��c��._"^g�)�|]+����hH�2l�"a���7��p��6��|�ϻn�7�{��++%Ë�ެ�. �	�R=�P#Ȃ�G��$eO�V�د�TN��鷁�������@)i�|���9��r�X�?'3�0�����%T��F���Z~��)s�|P��w7����:��c@���7��Ztu���zQ���g %Z/��X�(P��њ��P��Ͷ6I�3����6����l*hlV�v��*�x�� �a�GH�r�q�&�W��{�󤥑G42�L�
 dO�MG_Й�OX�,lu�o�Ob�c��s�r^�>{�+" ���`�o�r����q�; ��q�<lb���QTu����$��?k狓���X��?"~SC����v�i�/&�_ꁱQ���Vg֛%��i@�:�I���i�Hv�%mn0���(��~����k���ޘ���b��}ַ�[��h`���bZK����#۰v�ZƤx�^�A7�#P��0�Xm1����s���QxX�/�b1��ڨ�|�u>��]=�Ѡ6������n=������|���
	��8g�������̓nW:��FNxp�\ڗ:�q�$a{fg})RQ/��G�|^��;[T;I��˘f6b��d@k����ֶ��ǁ�!k��.���΅�ꭤ�G���'S��H�Y4��m������͍��N�Q�R�
�J�6(�p�f���Z���a[���m�	@�,K�����X�D8�c:[�7zq�eL��7
��o�b�ތ��O��4�n,�I✽MG8YBI	,��ux��<�lZ�w�g���!H�p�2UP��,�(����B�k��₉���.<��j��i����;� �$S]�tl0����R�~%>�83�@M�����4�)(��3eVV�j �(�-��ב�C5f|�R1�i4�I��~Q�	ӥ�I2�amh�Q����}�ғͯjw+��+�z�����-�$p�pIC/mM��D	�ԡ�f��h&�1�cT1aR�`�l6̣�����	�V�r���AiƬk�����[��w�}`g���R��S����me6�A@>�(�����/�|:������&�����3�G"t����gd���'�M+N�����*MSw��H�K)�+@�\5=ti5�(����v;x�����n����|��@P��A\�����5���5����ʦ��53?�T��{�[vo`�Ӳ�`��	�H��K�sK�{%��'S�`��c�����Lyc�AG_v/��u'�^Q��oQ������7 ��St���H�T�̭J��O��A�x�"#�e����UY��48��N��Ͽf��*ٳ� �K�Jˁ�������U4a,��:��Ա�=!��9�!��<5��86��dJ٦�KK�L�_w2r+.����L.��L0	Z��骧�u�0��h\7��E3��BO�hܘl�rJ�?����1�oգ�*��z�����D�_�W��m�����B��nRn�)kŋ�w�~�/i[O�9�f2�?�=)k�ct�*T֚�,�;6�������`Vrxٕ����_Q��!!
Bov��LC�c��-����x�7��fu��b�R3�jRΑ O�(�O H�3:�1������K0U���d�y�$���!U��Ɖ ��P��ʳL�0�fb�> M\�ѷ��P�
9�V�+P-���#�(=2]�X���6ױ�ix���a�	J������\�O���w��rN�Z�	R��P��%!J�i�\~�*������>�Q��>�oqM��~��i��ѽ�U��yÖ@6�d5 �_�5�u�\��e]KX=��i�[N!x7�(�U��4Oʓ�3q1ZR��p���X�R���,��>Cߦ�Tܙ�uF 2��Il�Q'-ӕ�:��E	�`�+U�Y�3�������`j�r�vfX�����Oأ�!�ȯ���,�F�葆�ޥ�T��J�KJ�?��+�_ͦ	3�L�e.wN�g�o�0%iEZ��ף�{��x�\��&�p��*p�-xN���G{�� �6���o���w��6�0G�쉋��5��Q����P��r�0*�\�vI�J��ؚ�<�\�a�����)��z��{�;�|����w�-�\�^w���km�\Ƴ�ı���(�b��J>���G��I� Sw(�P��2�\�ն�n�1����KfJ�b�0�y��a��2��
0]�l�2�lu�yh,.�k&0�c%Y$��;��az�p!���`��!L��8_�������t���+�y�JY�y��M�Nϥ��
�x�VZ�jس�Qt�+MXsx0���������,0���(q
���z��������N��M�/���+}('2^�A�x����ƚ��y8Bo��E�����ڋ)��:���T�(��Q�X5�fi�I^�V�l�_�%!a���d)�3�0���h���ˤ�W�A�(��
2���~xe���/N��CF��J�OT/^:ح7����6m���}%���DB��teՄ�lew����؋������lu�:��-�.�޾����l�܅�W����cwA��k���̖�sV�
z�j#�OXC:hhT�)f��e6ED�T׿�
�'d�Ot!V�]�Wm�O�vĐ��BN?���˸}�����A"�_�ѣVv���M�y.y�;�i�t4��?�e&��,������r�v�~�e���I&��#1�#Z�<���$�0"flS�ϗ�n����.�P���Z0����	L������P�GN~�)�RXt{�;��q�pj��Vrà�9!Nf���f���A����Q��P7Ufِ��Z2-\�|\8�n��hhY۹K��;o�������ub5��=pKLG/�*@+�IO�f�%ܖ�5�|b����F�d���b}ߓ3���g�U��P�~�8,ؼC�Wq\���FC�W���#�Qs~�8��1m�B��y�@�[C�1�,>Ha���J�#m��P6v��	(�k+i)��6�8@����B;�g�co�	�����*ל�h���|I��ȥ1�:=��
���w��*���������W���݄����흱
��E留FY�L�B��CS��;T����j���v��e�K�c|D9���Ƙ"d7�X|^��RPۆ�D�hg�l-J/B�[W���OYd��jŢ�L:�B/Y���h���22~��,��g��Z�ID?�ƵŰ��O*�0$%�+Z�xgL�kH��5K�M\�^M�փ� !�Zq�j�XA��53s�83j �������E�N����-�[�Q�Hj�_���tӸɤ�x�w@U�!s;/�uc�έ����`��������_i�*�Z�����̈tt�ɉ����|9�,�6l��1�r|��6_m&���;����T����-Ī��K�RF�fd��H�۬"��	��_���DW�-}U���B�F�5�rh�N<�I�������ɨL����'�G�N���8`�Q���Fp���o<uU���*A��S�>�#^�Y!���K�M�+%X=�$�:�~uHR��e4l��{'ꕯ�n��Zs\�VQ��)����y�e�_m���
�*�p3[x"mT6��AhF�l�V�٧�J�Gnܹ��k�a��!�%�l�{!�������?���;��Ҥ�"v�*�
��u*�(�!����ɩ�9u����g��)8D���f�4���@��>=��U��׬mF	~Ub����">�:�;
ᙗ˳�����%Z��]f�"<~3�5BNk��H�����	�I�3U|���@�����MG��Q� }q�o�l�}A��|�&�v��@m�-�4J��U8j���ygiw�0R����ݧ����2o��l�Z풫2rx92ھ��	����<l��X��<�,�[)���ߤC��7��b��L�,:��pA��ê����$Vf����/:�L����8m�M��gՍ�t��3���_[bQ���
��������ce��1�/�L�ܘ�8q�k��/K�ߐ��6:��z�f�M�r���Ml�vH�~�VQ��(���F�)׈T�XH���BC����<#LH��C�6���H�Pн(���
�="72�)�(5@BBz���P.q�
@�<;�R�q�, �*>�~���!��*#��]qYB����t ��4�8x֎���/���w��x{�gU��١�~ۉ���y�#�.�������&^�t72h�b���M���XA92J�UrYFQ�[�5�t����ģ�CZ�]S�퐔Ե.���ax�|p�F7��p�P:�q|?$�?}&��H@1B�����Z����4���֦�͎�#�1��͑�Pn�U���8�<��2�u^N���[����q�5�3��_��Ts\���}z�֌�T/$��^ƾ����<�2�:h%o�^�4�c\�"b�l|�l�$��_��1�ƃ�NlC��[li=V:O(��(`�P#D��D� ���(J�/�%����鮞��s|�C6a0��%���2�j��o�%I�pPL" &]ʋ�7�٢Hm�����t�n	(�8s��TчC E�X�+��n�<y��B�1c�q]�^�11&��+6�[��1�K����J�]Q���T��mucL�V�a��hU�9���[A�`lB�E���C�Z@�'�d�j�"�|��P�h�!5<>Vv��>��(-\@\!����}CB DR���+�K^�x�;�(�b��eK��8����`e������˛��AS	�,U�z6�ԥ�uL�� YPʵZ2E�,��\�Cf�[����B%<w%ʆKG�~9�Z�O��z�&�-%<�'�>SZ�)��o3ye�j��ܴ�e�,?Z��؝.`������k\]V�<��h^�¤� �����X�ʚg�2�ųi�e�xiJ�mZ�6G)�`����)m�(�Mpɨ�@��q:BE�� �{>�zB㩽*��
O��k�v<�k	&J����&�%�tژP��	 zYv9E:�(�U���C�����^`4A8�&��[J��C�&/fѷ�l��z�FE��UM La�x�q�6�W��4sHN�����r�R?X�ʣ�zR�FD��7���w�Ao�I����,����"�h6wW�����5$�7���b_'ܶʋ���uG��so2��<��ew"e3|`�&�ņ	S>�;UK��ڑ�.J�����ės؇�Ԃ�,�Q��yv�`��]K��|��66�H���C��>3��1d�#V���MRr�uny�/�����"~b�FRtqt2S&6�N8��8�>���R��.R���Y�u&/8B{w�!B�x�{�p 	��	�L0�N�v�AyXf����Y]v�/���K��ed*�*���Q�WvG[��Ao��[?�M1_�IW��O��ܝ�*´���}TdY�����0�e�	�~�I���D�<Wx�)a��mEr��$vR�\qO���{7��~r^
J����*���D�<^R��|w3f��o�sJx����g�M"�(n�K/}Uܽ�������K-P܈�*d#�P�e�*]t~�D"H�@g�X\��ѫ);$z[��$�%G�05:�0����Rh?�<�yY,	��}�&��y�/��j6���v��q�#����|/w��wD�4+�6�v� W��0i����--�%�;.i5�:8yuO�uL��@T���G�!Y� t[�� T,T*8f��$�_l�Z��
��<9����p�(rs�u�N��=/���k\��1�ם�n�Ҳ��V3�G3�G$+/{�ѼC����A�&w(��0t�,!,�����<%s�����Mz[����`Ft;jB�Yt�Hܓ�6mX.��'�k�K�	SN�c��J�k̳�$�B��9K�_/+�\�VP��D=n��b�J�����ҋ����"���'��P�,��PV�o�n�fF4=K��[��4����G�Q�w���|��>pOZ<�cM��A����t	�X�GPk9�H��}��GB8FŘ������h� N��K�δ#Axw�MeK[�_���C�2�F���l?�b�9� Edu^Q_�0� �0�
/�j�T;��T1[�j�b�`���]�T����tZ�-���EuN�x�+) �h��	�I$��N�\>-7)y!8EN<�25��<�آ��]��LUV`L^�&~���u��ң�I\>���N;ow'���?�(B�o����`�y�IPہ��1Ԉ�nqa��=!��[��ѫ�9x�����?�O��+�>a��k��+���1���rUO���ڛ�g�͆���������^So��/�����(�TX�+�l��䐾"��Py��f�"�B��=r���hS�WC;u�N�090`_.�8h<C�z���;D&&m���
�L�֯��]q�3���S�s��h_'�Z��Ki�C��~oر�x�4��7һ9�a-'?4Ǔc@f�;�/��E'��V�K^st����b3gzMe F'���Cs�x]K�˥����2xb���U�t�~OZà�·)=�?4V]��]&�0�U��D�9�#J\�W���ی�I�D� �cU�x,9f̈��zH��ju֯%��m�� ��p,�G�3����
B�67�BR��*5N��@�=<�W$J�e��9e�s�[��L�>�c�>?خ�(/�Z��"(����Cw6���㓴�;�DO�Tx���^�gJH1:����	�^�!"_s`ֈK~����O!~o�k54�]g�����:p�֔����y��j��N�g����7�8w��ٹm��;M��f���[
Tͽb���k��%���k���M�E�W����*���}�)��\Cc;kv����S2�t����Q�*:To�VGb�!@sI�O�"ԋ�,�i�P�^��g�u�'\/�K�$��~�=�s(��LT�P���ҟ�Q8$;ieW�s�R�`3�6AKZ$t=_��4+�hʡ��+���s%ǃV���BL��6O��P�WkU�^Jcz@7��5�$����CzL�,�h�k�����|4��''�T�Bo�3�*�1V%�m�B�|��Q��^L�a>���.|�(
���Zlw��i�B������]��:�]�k�O�o5�ۚ]s��C"���:�`���v�ޭ
I��t&F��kPj9OS��� : ��Aσ���*�qfz1��J�j�%�+���~F��d�vաH�u��N������������ǳ6��T����H��B>�c���� %`����>�����#�2�����:�3�Q�w��P��ɰi�'���xR}7���v|a��M�$��&��[�%���9!z�-��j:<�ld�>/d�ʍ�`D.]�Ҥ?�I�l\��n��/�;��~�L*^�u���{�Pܕ���i���Ԯ��g�E��"qzܼJ�>��:�`�@hy�e*��֯,G�K��-���7:���ǜ0Eu�.U�8�
��;2�tnR�¼�l(�+��!`����K:��7"�V@���Q�o�I�0y���w� oէ���C����![����j��"4�����z6^��6>\�{j#�~I߲r��@{�t�U�ڮn�Trc�T3u�)��� v�/Z�@��
d���T�j�P�XP{����1t��q�t9_r!��#����������57uE��y_P���5�(c�T(찢����	�!�l��\"��nc���-���M(�)�(��WQ�cCx*�$�d�t��}��eK�w��,\� ��u�T�5J �LuP�tu�c�ʅT1ģŏ�6�
�JP��+��&(��+F���Iwl��`���^w�0�`E����g�9R݂:��V|���'����	�8��s�-��'� ��6oeə����4��"�{.��@Ǹ������E" ̣�ƥ�/�&�ĀzQr�վ��~���G�A������O��;����P���X��� �jN�3�yܩE-�qa�(EK���T�s"����P�<�U�4��4@P #p��~s����4���p\���L��e�¢D�Ly<BY������C�tr�h�6'h�`��]4D<vĞs\�KA'~o<W3��hW�e�G�t3v������f��Ǯ�:�!M؛㫠��To�	i�S'�?��_��K|������D�r��W(�[P��uK�;7�dƂ�� �%.��FD��
�`�r�F���~=`=�a�����Ŋ2�Z�Om�I��̫xqx^�1$�
�3.���L�^��/p�s�`��>���A�	�oJ}����,Ӝ�mڴ1����['�g8����[�EqΠ>��� �n�C�si5m�(�0�E�iڬV1/�D�e� ���x]>�����W��>�/G�19��c��O�i]���1_ּi'��]�����R�ԣݕ8Y��=։����m�����S��c�M}v�W�:N\m9DB�cr�Ds�V�J��0�y��:���8��� �o0��9�����x�;ڭ;I�#�0�����K��^{a �?'"�f�!��2舀pH�S"��6�uOG�~z:���>K��.��y��N�y���X+F�a�����޶�D�s(�6L��%�p2��B۴'���5�B�Z�`&��l��s��;���=����;�A��%�XV��i��Ͷ��vHg=���^К� @U7
]�U��~�S~ABe��hrf�V���}ܣ���ky��h̽��j��ϟ4ٛ�m��>���r��Bt��ۘ����=o���`��U=K��2��V�������NKG
��0kԮ�|x���J�H���c�U7��*l�C��t}���Ԙ�<��ګ� ��P�b.�V�Y��k7F�s&��Y)|�
���^�T&���|��8⭀�Oju'��[��T�J��s��U �J�~0?lX�C Gs͊o�.$,GLQ��ݟ�`�����O}15&!��P"ƿ�<&"<9�����\�����jLL{��*�L�f�r��=-�<�?X�ej~gc� �wC	@x���zL8Ğ`���6�^��w�`�P���Ɨ�,��^�j�7W#׀��ס��i�q�p�<Xv�$�������Q�g�!��R�����Ƃ��y�_�$�j�|k$ӀT.t�����l��=aeenZ�%|H���f�xH8I����jk��Q6U�<�k�M0�T����9"���k���j�3B���)S"�f�sF�
i�9oYh$Jd\��OF!���7N1������$$=-���$��X��υ=�m-�ԙ)M�ᖓ�R���\�r���wEj�n���x�����P`���@��̜����jO����2���5�����:��O�O�/9�P�ƈ�ƬC����`�~=�^����z��K��s�4�ĸ@>a���	q�|-�|N�~'m1n!$��|r�y*ѧ`=�_�����Zhd�^���sg�F��N�t*cY�c���;�%�̽Mq�����ZR��S�FKU	��1P<2����#Җ�	}�t�!ƽ�Y�q�qN��%����i�R��x���x
�������g�&����߮&OW$���Y��85K2��a�GL��Z΀['i�7q�����M<P��:A���G�7W����MW����202z�+�>�^�1��_0�� �{{�ն��=��5�K��N6��4�y>L�IR)��|�ڮ*�(AHXDe���$��ycK���@�+��Y���g�պ��w79����v��`A�$�dgP�0�[���[6�� �z|9����\x���

�x9��芷%,^��ݽ���;�.�pFLݗ��Nf¹u�هy��UwA[3۰E
:�Vn.��"wz[��?�]6k���piRQMTw�}�ԧ���^p�⛘$^�@whW��%w�UɨCu=�Mʌ�uY�-�.h�#�}<�[���
躗��+}T�rN��J��ҝ%pK��B��b@�E�/q�­��0�Z�dv�����ba��%627$�Sy�8��-�&'G�C�6I�1ܿ�.�����k�ެ��5���2&WZ-3�K�Y��#c�-)t>�(�����;x����txfcP~{9	�p3�7�W!�����ٹL�~�Q���p �߾���ʸ<���&���~MXۈd�������u5[4@l�z��9��#���|Vr�H��7/�懿-���"�!c�r�+��W�.��`�^�M�1^6��Bg�W���Z�+���k���@'�~����܂�j8�<��;;bB,Ҡ�(aPH���e���ڟ"��c�'iȻRP�qڨ%l�ҸT�a�>�����y�5�1�8&�F'�]�����h�.}�F�W�60pP�(�Ѳ�I�k��Ywr�lW�PW�9���t�����zmEPl��1������H����{��]a}�*|�[�&lxS�����p*�5IR�+���-��t�&�J��cg���R�v� ebp�� �c��hU�CL��O���6�H΄2��+�)ě��ꂣ�r��e��֡��2���E���ʔD�#2IN��"6��ʹ4�E�Y�?��L���ߘ �9'�]#2奓�]?Ǟ�R>��Lɛ�Jk�2h5+%t�N��8xiiA��^y��i_����,��'x=���x ���_/au���p����R����ɞ���S���A:ѬeG9��A�53qU�]F�����?W���mh_�ⴭ(�aټ�	�f%!��S""��QĐk:�N�h��k ̜gM��gϸΑ�rR��4�}��]aP�
�۲H�9;Bܫ/
F⦁[q	���ծ��������V$������{�:�z�ɶ�A�3�s��C�t��]
i�D���I�H\|��*5,fGTaŹ{�Fn����p�o�<�7��ċbͯ|�� ��o�-R�&DaK�e:i��Nol������Lk���-�U�����J����`���8���b� Ul�3}�|S��|Ni-#���J.��u�Pxś��v�E�sX�E9�m��iSs�#��s�\�A8-ۇ��3e���1]z�t����3��3��(���?`<l�6#��\HZ��^0����.e��!=�O+7D }�9�Iqy�m;�%ι'�KRlB�0��}&%.�x;���U�T�qq�,t�( 68T��A<���"�J}���0��IU��褐8\�#�gDq��[�p��0�%^�3䎤�ם6�z��V��fKT��h5g Z��]�2���Q�����P�.���Q�\��F��$Y>8��VN,ؕ��b�ws�����-=�v��b�\�Z����wz����8�'�̋a���h0�س~&,����GZ�1v�%�/'�|�3<v�R%LOм^LXS��C��hzx�Ϗ�<I_�P���n\7�-�Kz7�q]������Kٞygκ�y��.�l��J���/�yx�쌙�,�-�2;��X���Ud�!�$�����m׎��9�y6�b����H�}��Ck��y���Z���,�ݜT���@[�V0uz:*���AH"���i��[ɩ��`�C�����yj�`�n3�@�|�E=�Ԯ��UT����|//=� ٝr�^��W}����o*.������Ӗ��9����h��C�^A"��ҷ�ģ�g�m��i8�:�l�X�Om�b�e�+�R��8�nlp魄2��j;�y��B6.9'��H��d$�0F����Ǥgv��k)?6XlA����5� nEX	��q�I6Ȝ�>A�Js��F�E�5OR�/1+m�NqP��.#��涽�L�'��ϛ�%~r�7�p��i�G�i��!��%/�8U�y����f(�����.؉iq	@��	��Ԩ�_�"(3N�o�|���T1E��i.��ɮ��kv�dg�׿�(���g��QoZ�B/Y�Q���7�[h	0#Ȓ�3DDd|��Yڕu��)B�An|}�~��С�_�S/�|�6�~*!�X�{�My�9�b� ����T�\��k(��yIR��8�Ж���1��k���e���b�O>��p��J�Be�W�:�4�� v��������&�,hY��>��m�mo�Z�	�N¼6؈�V��`.�%#BO�{4ݓ�?w!f��)�V�h�����9H���f�Tl��8Fʞ+����,�<�P�P�*�����'�ַ���?Ł�ԫ6��<<{���jz���iS�H��M�H�l=������){̠I�z}�1�^u��4��
����lG��D����d�j8�+��/�U.�ҷ<��)-�<����NCV�<���V���4\i@r:ef�|���1�������k�c�|ш�y��x��%�&%@K��n�S�T��V�����q�-�! �>q�(&���Bb��R��ki�֯)�P�ZGB���	_ذ���7����v��[���$Kp�O2��ѨM�?���M'mn�SquE!р�z��Wݹ��yX� �ݫ�-x>�u�?ၑ��7��6)oR��@]�ͩ&V��>f��4���}�%���0I����� ��ѩlMng��PMNZ1tz�!�u�젚xA4e����"|�%�]��
�p�KE���B?e�k��n�r�Ћ^��nmѭd��s*W�<�����[�}P��m�nҸzZ�ީ�\g�R���,���M#Z���[
�	�͟��sCN���Y�3b����KV���H�47�C���޺g��k�7�YZ"���%���p�]t��� ���y�JWv�h�S ��r<���O��z�T�=qOձ��`��ܫ�&��(�4l�H�m0�QR�I��qS�(��O>�~&O+���R(1�7VP���k���L(���Q�z�O��6S��lW3 *�GF��H����-ճ�"gO*5�v���띦z�f&��:)����<�-�©���M��9rs������+%b��o����"�n0�p��&�����_h����S�̹G8y7��B�*}&���˰�D��)+���<8���׶�(<9.Ap��'h��*�=a�/g����Ki�N�h�J"q��~�@U�HTO]I3���a���v��-k�|�5V�C&�C���ϝ�p���N�8��C���"�Oӄ�Xh*\�)���N/���)3sW�*R��hɍ"�[�"}e��p�3$��ǎ�^o;�~�9�?��0t�/���4����L��spg�k��9Ğ=�p��V���=~2̶�1�Dc!�=���mĎ����xɄ�%3�PqF��yO���@`�%f-�%i�|qiU�M�%���RP�~D�PVj�.�1�ZC�f�5��B��0���}aлG��K,���'?:�}Gz٫�5�{����f��~��~�T��؇�|�K�Fb�Ӎ�T��;[���HT�%��؊u5E�/HE�0�#O[��zָ�Ղ��'0&�o�^��9v�-TM�a�:�)���"K=��|�6���[3����V1�񎬋]��Sf��}P_ S�5�=X�=�m�EY�羊��Ґs�fe�A_~
���X.-������B�F� 2P^�EU��)L�t��p�Y��>���=��� n'5�}&�9_ m��u��g�"���Bϕ�P�H�|}�����M����eUw:8�|M�7��K����x�B1`�j_\aOf�D���ww�� ���eɩ�>�e�c(��!�w�����&ڄ��_���⊭J��Ϛ �.�ۿ��_75i�H��:��:91��h�KoxEGNc��)����F�,|���	�b��_O�+}$3�����Z�][��A��VUK7�
�τ}�`A[�c��i�
�F���X�����(�E�Uʫ���=��7(S9I���v����,�U�^��U�1�;�$�]�l�rs�T�P���lF������/� ����-�Xp#�f,�;L/q���9��L��΀#�Ԏ"���f�����@�Y�X���`l�=ɋ�| r�@�~V]�7l܏9/i2�r����E�i�1���L��Ñ�P&r��H��%น�� ;�Z'ib/�46�Κȟ<s<q��α��*a�~���5i��]���Vʿ\xo|7��Q��Y�=��ck�x��sTs
��2���2�����u" ����T���"KP~1����uZh�{�@a�2lL�뚡z�Ƽ/��r˴�hgm��2r����=�'-X*5���Cj�x)L�%������Yx�	A�j�6�C������a� ���2}�I�:9N�t]o��^��(o4�)�E����pMT�8EtM�+t�Q.�!*�S%��BP�;c��K����{����h����R��~�ѵ�%-�h<����|�u"n,k ��;hy$X��_�]B��e:|^5Fn��+���v8�M����e��S�^����F�����:\��]X���'�NG7�کR���@�:E�)N�ʂ�S�dq��.]�=�%pт(C[%d|�N_g�S��ӣ5H���e���bQY�,P�g� (=���Zv�(�9�D����C;4�`�vR��Z��'-��yq���L��#�����j�r-�4��+Ŭ�ث��z7ߗ��v�����e��k��?{�X_�ڪrQ?Mvh.E�>�����!�t��g�������pɍN�M�`]�6��<
&��H��QdDk�\�XT,��vkRe���nK�w�s{��c�Xcل�&V�`t�ɭv�3�M♸����	�������������Mެ��XV��P�!ޡ�I�@�������H,D�Z�(�(�)���32Jlz�/�
�+�}��8���_�����M���������vI����B�4�,��څ���`JH<��V�̴ߪ��9�d@>ɲ
J��'�*t�W���ֳ�+�E\q�z��ˬ�s�������⬤#(d��Ɠ�.�e�X=ߣ4V�GZ�N���*�u�%R��6q�N��R}��]�&��#m�X�q�UU-�QѾЖ;� G�����ː�;?Τ;PN�c��Z�m�2�?y��f׃�Y׭˟|����B��e���	��Ͻ��@�*ur�WuJ���u�q��b�ǭ�@�� W/�9a#9Y'[5����;���	�f��Upw����OH�诟��v�����k��է�ߝ��~8��5���px������U�yxk�Ss`�|��β @�� >���O3�O��514cBl�[u�¿tZi�g0#���Cz_�_�w�
�6��J� ��ך�6-�$
��õi�u��v�Z�ͽ;|N�⣦X������Ü��$შ�@���2��A�f�i�����`��O�	[�vB4d'Q�)�5�Y����n�}�lmi��#��6�ћ\�8���A	]l��g�cpA�(/�����G��ƴ�_f.�=������t�|�3/������G�4��"�_�O ~2��[�^���~���Nl>����Y����ɞ��4�_��ɧ���ުg���n�N�1/{	J�tW��(B���^�c��[{�6;g*_��^'��Ⱦi���BG��w��hSQ��?nж�˵O��R*����f0Y�C��J�c��&\�/��۵0���*����7ҡ���f���yX1Y���z�+*Ψ1��NW V��s;�hX�6�r�⯁�j��VJi6�R.}HnИs�B��+D �]�����s ���q�]���� f���:^���5z����@.�0Mx���~'�C�/�8.Q��HK�O6�+�6�'�D�)�W\���op�b���f�+!�	ty�{e�k���oT��ܐ�P<u�Q�~�h�$��VvG 5'��(��>AEG��P���O�]��A^)���2�K/��D
�'��|��w�5F���cIEn��~���6�Vԛ�_�n3�[���w)��F��$��:�N�h�ȋ���{cs�pK0G��Ϣjʺ�J�����8|w���k����0�B��j�`��lKn�L�%��&����ElU��� R�[�����K�FFC]W�Q���Z���]�O���:PCg�����S SL�䫃b����~QZ\L2�`j�jUc���i;�i����uo��2u.���Ǝ�M	#�\e�0��<? 6�>��4.�G�B�K���m���+����1�P'Q�R<� ��Wn%5$(�:�jTCѧР�y����;��6rـy�ɥ�5�p�^��a��M9���O�)T���B# 4�O�i};��џ8fU�x�(^�-N� �)FN����Rh�j�r3 5kU!�P5�qq��ʮ����?5�{b|P��@!������{�t�6�U XYS��Ol���$�[�|��]�E��t����/Z�q�ؔk!çЙ{�T ��-���c�tֲ���4��M��x��<6t��T�����z:�5�2��>��×��o�'�����]͹o��[�tj5"�We|[�����hڟ@:nh3��hl�}��+F��} ����w,��0V�>�m�BJk�.�SO�m���v��)O3���J/������o ��1��"������c}� ���4zm�O���Qͅ2 5��s��ǃ��Ig�8}9
�}а��<1�u�L��q��O>y�Rس�cI��4t:�A�9�ܤD�1:��p[t�r9
�tp��B�<ک�Xi�V!�HTcw*�y�Վd�S1��s=l_0):��d�E�+������2�~>� "t�Qk{���w9i���$P^��R.�oeG�O�Y�K�QY�;M'Z�ƽ����o��;��Nݿo͉��bq<T݃�����&���nL�����]p�p�ry�K̨f�F͎2@��x+�=Șa�8|t��C�Vq˟��=$�x@�o�O�� ��h4P���6��Q(��6��Vro��2q�3ps�s`�Ty�8ͫ�TFN����\��[�"���F����Pޮ����AͰ��=�z�r	>�B�\�#�Q�4K�Oa$F��l/��3�)F�r��S�4�O�Ц�����G�x� 0�1�t���W�yqg��_�(�/2�.�;�6c}��M�W��S�*����K�����c�-�  dn�trC�0U7�('h���P1�i��������m�c]<��P����SP��6M��ۣp�����m�OE6U�1�x��o���8�Xv���Puݢ���2#�{��V���T�lĥ݀�SA�Go7�S$rE'�6cPb`��q\s�w�Y�sm��C�3�<Q�2����>�-��ƍ�\�{н�eT�y��Lȼ�+}�fo����2��w�L�ǐ+����~�.�W���]��]��z]���)u�	�#�l%��Q'��J"֓u���ap��/���[�`�;"�4�T�2^�b������O����=�r�|����7�E���$�J	3�F�܍���+�d�P���n�s�=���a#�TR/�NBw����q�|����r}�����㇤;�FgNO���)3�6_���h�v�kQ=5�Ӣ��g"}C-���:qNw��2&�k]��iC{�#0�3���
�3�|��&s��Q@�4���]d:�h��;Aħ��Υ9{y~�u��|.�[�>���u@�`F��T?��"m!�:F�Չ�V^t���m�)����4��Z6��C�[G�(��;����\2�x��JY�b)r�p��|@~E@�m2!]��h	�	-]e�`�X����������#:H��p;�G�8�w��l�Rum/������H9�´�8:��v�ߒ�-���NX�#	�b��8ت`����M>��;�0��c���$���!x18�8���*�$���O4o�%�@Y�UN����%�g� D]���S�Ë�;�(�%��#^s����3��K�g�����S��=�IP�J?��m$&�>fkŃ�'��9�{�,�:��1� ����8fL~,�f`�zlys�$F�y	\�U"g��D�q��!�����ȵ��T=� �X���:
 ��h=g@2��gj,%YH�Fh���Y6+2!��f״n��xE�������ܐ_�[ �ٯw$�Iby��h>�V���\�	-�O~hԳ#���,����E��C������2��{�<�@؉�o�[�|�[�}؝ͮ-ֵ@����I�y��yy3�n�֠�o�2;?n�^8D�����,]l�Z�t#�͡ɧG7��Rd�ǳ�zTʛ{�°��B��b����u�ص�fY�}f0CJ�]̂�ԉoG�N�pJF�ֹ�DB6�	aZ�4�����Ok�W��#�Vz�P��2�TϹ�AΜ@,�`���MA��r��~��9�٠�&��9�e�U�_U%2��"�2S��B�h�F�D�9eU {�p܍�E��X���
��:�/�W2����)�h!s,�C�7:��tы�!�������0�-zF�5�@u���[, N<#�p��D˽����z�h@+jM~�t���{Ć��7�vy+�䑈���'����܁�������P6�MC���ű|�	tF�D��u⍠g���X��'��\����P�0#G_ja�i�F��'F��g,T@��׮��h&�	gmh[�\�����c`!L�Qs��t{Rn��Gמ1"-�s)�*ldW)4�|�-�r�Z�f�B"B�j�ٲ0�7^�_���������l '^��掬7��}��N���4y!�b\T��+ǋ|>n�ϝ`�������!7K@U���F�~.FϢ��)�э����B�8��R'�(���;�b{r��l{Q�T��ِ��g�		xWj,/��]�����0����~�'�W"zGKW�C8&��sʤ��q�؈�� ]�"�/����k�h��2S�5�x��#´w��;? ,c�C���dv0!`���܂m8��0ĺ�n��UL�׭[vk���T�ĞO֥n��R��Z����.�Hpaf<���(G�7� 7j!U��͡�K+���x�
|�DKI�~k���^���h���?Ɯ��"�e�a(Ԅ��eS42*�W$�,r��T�r�N�o���ފĜ�z��D#%��C�&��y�OZ��(M�&�`(O��	Jܑ��w�J� ��Xf�B2�7=*��e���=h�@�e������Բ������D��mѻ��lĉ�{���r��}U����6|�ڹ;��4#�������<Dpp�����ttW� Ʀ���B6�����5u-vb��X�!�������P*�
��4����.s�ű�����a��LO������.I�ďF!0��}n��8G��WcW�^���\s�b�Op-[y���|��b��X���(������}Q��]��	���B��$�1��A��ϦJ��|�x��U��3�3��(����Zi.,v��㹮�K����i(!<MZ�0J��0@0k�zP�{t�E����+�����j�x�^n���>�%1�^�������Ni�k�-�ђ��d*�� vэ�Y�٢��A���6�}_GМ�-H�LҖv�j�O�����:f"�}rr����~m��H� O"���%KN���F�wxX	^9�&����cŎW���������G��2Oe���:��HD̑֭#mE���ƮŦ�5���!|f��R����ݔ;�)�/��G�T`�����b?X�xj�蔥1��2���Y�\5ס5��J~F\���,�[=G�Q����z��)�\�Z����NI�B�,A�9��1i PVV��l�ە+�O��Ku|_Am����e��kam�T�� j�`*��h$}$T;Vtj��j��Z��p��Q�v�ߠ_A粛ndH:�k��bɛ:��Lș�;=��I�iU8�)���Z��I� ���\wI�>>�$��|(5n�����P���*j�:��`�H�1�a�ϗ�bdi^�w��+D	���G��?�%\UO�ɐ���d�E�n���\�����EM#D3t ���ٶܓ��D]6�/���?��j�>�e����?UC��8BF�.���DN�]��ML�/�"�C뫺~%KF/D(�E��  �]'�#v�:�������}�ti]3����0���tҌWD�#u�=�2�.�hVZ��A��Cb�ky�N�Q��M��T/��ɰ����ر��@����5V�stmo1�g���4�wJEl�k��jC�0ȅ�;É%6�T���}נ��8�G�'��Z�e׏��hL���A��=\��/�5�$��:�8��'Om7��=67�� �KݯX�k��r�|.�:_�u��3��ZC(P(ݔ7'���.wr���b�������Lke��C0Ο�B8'h�
�	��P`�N���$(�'���VMǸa��B�#n�r;!M�����U��yaˣ��$q-��܀�8��,H��C��_+�m�|_�h�!�:�X� 	}���t.�P�*�4e�V�i�(�<�5hbڡ|�%"���yC�~�<���>n��F�5�c���X8�}D"m�	xv���7o۷������{�Rs5�3{�)-�n�
��Ãr�!�!*����- ���� t�b�Co��`<ꃯj=��}K��g�]��{2�s�̌r����		�"P�l=]G�h|�cLhh���\Á0�a�*���D��Fu�,w�ݡGRh*9��UTbbĕ���I19)�$6(���Z�C�U�i���=�F��b��虡{�mW�˻�\6���|2�@/捚:����X�x��
��k=��v/��2W�A��'���R(��WgX��\pȍT�r�@��+����<�ꭳ�}��2]���oNiEFv����R����h�[=tY�����Ftz6�U���xR�l���hU�HC�]
$��l�]Eì��H��Ȱ�C��p"4�k=OX���㉺Y8�-Ǳ�OS�߲*ٌƟ`�d
��ٺ�Wn�9Ȼ~��^���W�C��)ȕ��^l�(����;��g��`�k6qC}�`��|�p:�ogSn?kۤ {��7����/J7��R�*��1)lmMw\}ڧS0�y�Z�}��ðM�`%t����F�mˤ�L��
�ɼ����oe���8�ud��NC�V.M��E�ZQC��R��;.�p�w��\E�6�d/2��`���Y���5��./��תj?�h�@�M��>�H'��$Q_�{��H��
G�X�9{	%��θvjӁ%9��N�b��0C�^�Qf��n�#�++&��^(�v#_���"=��hkp'�t��{G�[U1���@|JAэ-����a�R@�]急DS�$f�%7�г_�m=��a�$PR��k� .��Gt'�{\�>9�� 1���+%�!Ɍ�$;���#�:��U������0nY�T3��Yu<j o�aw.�	� �y����(�43��?D?�ϴ��5���t%B<I]\��e�C�r(�V�ad?`�QKC}���89ظ8�U��t�lUO�?���v���ń��yZF�A���p�r�B9d��m$a�_0�	n�[���GO��_v��Oý؅��V;��S��(��T@Q���G�R�x�a
�)/�߹\Gc^�ɲr�m��:v�61U��m`V�N�����ئg;X)�~c1K�!OAQ�q����uH��|��c��.���g�ʕF�c����T��eca�GJ�X���Չ�X���;WWv�_�~��Y��Ӑ��KA)���������4�('�YW~7���5�GN��A�#8�G�`> �-��"�4����δ�$�Y�Ʀ۸�<|q�.���5��Vh<�.��_�w��.�V*��W�s!-�ֽ"��H����t��h���~�QHxW4��X�}�+$�g�y�UҘ܁�P���2\�l0*��C貀�I`��u���J��N$�K�)�C�T!�.}"M�5�x��#q[�}�3"^�FL�y|�J�n�%Ruwt�� �
��"��������:��KYz�\E���}6���l�%���l��A�*S��tX��p^e,� �Z���bhL9��V�O��Af7��x����d搢y\��*i�(n�&b�F#:�d��	��$af�G����1���{$�;O��a�M�n6ܝ�X�-˜�.����M��+���:�NdG^����s*;��c9���,��=n���PSM��?a��DK��gAr�;n�*'��5ľ-�!�i�,�5Gk�ڑߍ������h�`�ku=�`��9;�@�%�}շ��hKؑ@��6�D��_O->�`�<��ׯ��{�?7���X�YX��!-��ԛN�T�4I#�T���쾕���~B~?��~�E�yfmz�k0K���j8-��
��X,_:HDٝ-u�������aY�p�У:74=��T��O��M���М�z���&��#�̱�����t'�*�4)��?������HF�7���]�X��Cp0�����������}g�4�c}�X=�
��!i=�:���BE94͇��~��d���k�bH9�<�$Q�{�=\mu|��I�>��ǰ��q���������H?��(VfB�:o���0kՐX+h����?ql��{����Vj�[1��SK\��	��/�s�U�_
�b��ƒ��"�S=�1}��<fo�8�������R�d�;)�K��N�t����2�¬�-T���%J;�V���8F� �̷�c��sJ�$�I�iŬZ�)n���CU��-�K!n�n�R������WX�ه-wH������$����L�C��{h�gZ��uT�zB���=V�z��"�V�o�мq�E�����F�)��!3i8%��J^M7=1����n����*V����B0�_������ 2�~����}��������/WS����7C��}�g�!�h�Ӈ\����D��~)���h�*Ut�M�fY���KЂ/��A��.ʲ?~�4#�:<������-��"�b��ނ�/��B�����\�>���mI�]�K3�Dl��
 m]��;g�!'�n!�����-L!d�%���I���޾ۑ�KkFB� Y��^�2�A�&zW�
��z�2��b�@ݧ��8V|�:)K%��@s����[�9 ����N�jg�_��U�E�8��bU_�.�{ώ�~d�S�4�*"v���3vb��:�Dl�cnK����A �{=��fV�%�&x� �W�@8G�D9����Sm�������ֳ�5�M��1{�+��FSc�OC�n�In�}$�cn�-;6�R�+�.����㯩"Ml�E+s�ؓ�$H1N�\�����Y>�F>�q<�]vS���Q
/�[Zؖʹ�io���0������PA��2d�t��S@ ��N\@_&٢�d�8Eu3��9��5Y��Av���������C$��T?���+��B2�%OX����-2n�Y���`g����%譌餏�ڇ3M����؃ܷ���Æ��s�I���TT��Q@�p��c ��w~w�4�4�<|�hK��ZO���9g���9�Y�Z�멥����k�	d@.�_�V�h�`�t�-C�ޮ��y8��`��h��)}Z������O�g#W�4���B
͍�^ ��άg"�9���_�ϱ9F�_�eX�N�
�"�x(+�9wo-vb�p��g%�8J�]���bs�/`6��nޢtŜ���T'n;'���^ਫ਼����v�>i�Ʀ'��|?l���."��˷��o��Q��p_,H�3��Vl0t|d���`M9�vH�"/|;P�������1��h�M�������JXV�O�8���8s��7L������FH�9��oN�:���<��'SJᏤŅGz|�Ŧ<g�'�&�p�^P���R�Gm���Z$�w3:�L���I��t�w�|����\�k�3�T�罄��
�'տ�& ����	��2�,X�|,�Ӧ�x7ᇺU�}L�����C@�oGPU�F��?=z�;��z�8���-XI�|����0�]W�@j$��5[O�Cu����t8`�_�j�e���Yi�%a���.�(�t)� �|�P�Q.�ĐoG�oE7��n���`��9肛�Y�@&����ӆ,ǖ���[y
sv�ܺ��}���&�h��Z�;8�qG.gڮ.F䭅f���)	� WdTE�7R�ioNlX�# �6E�W�*	��N+9adV�,gg-V���paAҪ^��U�,�)i��D�DҲZt\��y��8re�~��9+:s4�<F��k��P����h��f(m����Xw����"�M#<�v?��)����	"S�
q$Y�����G���������!��kx���W�!`�ix���e����DAު��[��w��Om�V*����Q���8A1�-=����/��&KH���y�%��W��<�b�״�z�!�n0oOy����R���� 0���B�_.��i�f[E9�X�5m9���W���n#C��Z��*�����)2X�WTN��:0�b��2���
N�n�b��f֩��ér}c��h�%
�d��rH����<��]������8� Z��
�
�] eHޕz�گ	ht��h[f�5&?�^�Uf�C�E�Hh����b��5#��v��������K��`�j����~�nc:�`��r�諩���3\
�'������1j�|t��5gb��	�0����b`���k���w��g� ���X� T
�Ol�ew��ܣ�"��"�=E	�t�GO~Q/!�a�hXwd�uY��)���Kߚ6,�EO��ݦq��&�]~τ��#�C��Έ��Z�7Gr��|5mkn�/���n��kN��&�t��v�ₘï�7�ڝ�nV�AFP�=�vk4LÀ鱡�뜍��7�\A�ReRe.���Y�!)��hY��6�(�
��P#nRܱ����`�j�.�yIN���#�E HUI���k��=u^Lװ	�^Qy��F�P/o�A�6&�̙t�tݯ+��[M���"X���A� ゟ���9�ta�����m��6S���XN	��3IN����Y4o���}ۤ�� ��-�D��S��prNd���"�~�X뻌೪���������RU��X`3�ۃ�+)�ͅ]���2��.lK@��[tǞ��s�*U]24�S����xk���k�2��o�"X����2�~�V���[�������(�?r����3��}�FB4j\�h����4���q�����W����OWR�&�Ze�����z*���Q���R����N$�(SY�{Mor�>���e!�9/�����c��6�������V�hֿ�m2����K�o+�p��$Ҽ��)�t(��7Ѡ�u�bK!��g8�!�����P�{*T1טT��9�^T���7Dfp^�E�8�e.j�qB�ޭ��K�o��/�t��R�.���3IW��q�Ϥuw[��-"s3�N\C4��M��^*�A�%�ޮ�e��m���l����Vo.�4�~D���]�ew8鶰�D<�w�@;�h^�QЈ�$eE�^�灄�2!��D���Q���S}���(DS�9R��%��O@�@d[�ȯ�?��ߣ�3�"��@WO��=���%��P�"R^d���gh���6,%~��k�7����������1D�cf�*��I5Á��C.aW���(�҂d�J�"�۸ gd�lk�?�+��,�����n(1���Xֈ�ဠ��J�� KU�9��7��7�+�qdb�*���[@J?A��N�Fy�-�^��2���K+�C@��e0��%�1���I Q*͘J������!�^v�[:l;���0u�Ɛ"y���2XA�`�������*\6�����-�dU��=s]�E����)�=D��J�٣�����0���o6;K�k��^3�n	N&�t2��pn�֞A��ji�q���+�ю>�q1��C��VdO���]'��{�X�<\�La��L������[7[�KC�fߪ�$���!���)�5�P�
�T�0X��!��Lx��8r�Q���Mo+E	��'悌�`6�~#�6��:B�Pˑ���}W��_ؐx�5gKo6��|'�5�$1��7UԤ��#��x/
�E����N�u	��:���b�y�R�i���6U���?�����\6�nD@�+`w�C-&��ݰ�����'lu=W��|So+���֬I�Aɋ��e�5�`"w��>���EE�g�ІR��e��7��e�8����x���]�Yu�7�i�ԩovn'�-}�|�'W��cY�œ�(��I��wX0R��Z�&W�dO��o��{��^5�u�n�8 K����觉��M�o�K������7+���C/���O�X�@�z ��I�1�)"��<��z���,�Ls�)�IjS�.�O��aJ�4��l��Da�褈1A�N5h���:��j�W��Ζ��-���pm����Q�Z[UpG�n��ȡ���j���6�bc
R�D�}����dF�HԏQ%+�<\r����E�Q"�����9KۣLH8~�ׄ&.�)�ރ��~�f:�0%||AJ����J��֜l^ =�E��c]�}���Â;OCz�8��W��ϫ��{���e�b	�~1�6��r��5��Q1��g�g2���4��E�D	���)�N�W��[1o`ǔy�t}�w�bW�|�&����z{0 ��Y��eX�T�����|1�y|$���񏄩/�+���� ��:�O�&�jo(�wʂ]}A�Ϊ�Q�y$�N��7{���r#�E{�@����x����/�xڇXm9�q��`�0-��u�ߤE��-��y�����u6�wpS�d��=�5��t�&Y�.QƩK�] �#x�q��<���l[*��f��]��*�wH��C��\
�ܹŴA������I
����!����1�fP|�ִ���w�Z7e��Es�6��vC���a��˗��Y)�(�V\�����4�(��{\DE4�o�ۉAʽ$����&D� wr��ۆ`���un2"dÕ��|��d�9�$
	�I���{�rv;�zY<���]?�W��,y�|�I�)�8�_�YG����(G��*�H�<��#x�����O��J�ea���sB��+jg}��f=7��$,��Rwu��a��׈Ҙ�t�G��z'���T�Q�-A�U�r��1u`�����VJ�iCs<5�i���gc9Q� =2���n���s����;�ܘ��9�e�7�d��� &k������UЗ��7 �8}%˖7_58Qp1���Z��j�H	���d������9�^�Dp(�(/�8aJ�Rcl"]���I�G�!�r����b
��9�n�,�����ߋ��ܕ�RWZuaQ8r����[Q"������I������Z��:��M�y�4��?R����{d��P���)cx�z&���H&x���)s9?�u���/���e',W档�+��jx�m6��	j�=������Q{"�&u����vXG�;�%��2��s��_���U���=���j����<���Q��*��P��^_�0�Tq�1�rR1���R5zc����� ���x������;ڭ�p�7�1�.���n��w�n$}��֫�����5Z���6�N\��De�~Wh�P<�-���W��1��^D����o+��_��+���V|n��*�q���>?�4�y鲫�M"YLBs���R��q&�͍��aH�M*�=1���2��VM��L��{��qYQ��!aU���g@g	=�-��X�����m��)�����Gz����ӽ�J�)�)�i�Vb�ɸ5�iz���ɮ+�{r�c�����Y�*>�Ő/�$�E󲲜 �a�O�&i�l��=�n���+����/bW��`R��yc�m�ׇ�Ȼ�D�T-/$��ǓJ�{�b��?���3>ƈ[���Zj��W�v˹{�����H���~��b5���!������5k��)ajiN�{���d�1c5��~)ǭr��%���jÑ���|�d�߰|������{�==���=x�ŬN匎8!�(���1�-f'瑾(,��B�{���a��'cAw;$9B�vz5;ҟ*��ߎ�(A�*[D�wM����r?�W~��2�&�B�v�w��;�Yl�1����Qk�,�d����~?���W���i���$�e�9�˔f֑De&L�Y��y�.�{�%\nE�G���l5,n�M��3�9�
8�w�YPW��Mɐ%r�",�����O��h����3���!���|n"�1���7L�U~j���"�Rj�׵w�֍���S�h�Җ'e�[J+�ֳ;�t	���9w�e�?/l�L;W"z6'T$"����&�� �Sb`ӷ{P1��>G������s)>L�I�P$�g���]K
06�����%�@3֘�%
�y�y~�G�Y�/d~P��ݭe��]�%/�?�e�#uώ�u����rP���a�}�ɕ�F<��U�q����NVX�Ad=�b�Lޞ;~I"�i+&��  =Պw����o���7I�8�mP�4a41�[�n�~����E=��@����YZ�������@�����L����A�'��〄�V)���E�%_`�pN�I�i�� ����}a<�7�2W]�=��Gy@v��J����b	O�9���f�إ�-�.y؃��έ���Ox〚� ���$DD�F�en`�� �*G�p�	\��څ��@W�����M�Hb��2o��A�"���<��LQ�։�}d�Ⱦ^����J?G>r{��o��\K<�E(Y�R���$F���8>%_ԉF`�`�0���VY�&���^�"W������ސF������E�o��1Ʊ1���N3��#�q+<f��a��P�LT=q��Y�Q�������An��<�h�|hHn����C�@�wTH������ԢHj6۲��6'�
����Y��#���>�n4��K`�ڪK���ϊ�|�lت)��݃]��Md՘�	Ư�ؠ��&���R'�*�v�����.z�U~*	�B�%� ���`ٖ���r�$	R�l�<��a�E(���S=,I6-D���6g>�^�F���YQ���	���?�F췳�d�)$�ւѐDݺNUT�z��g|��}.��Gv����.(LBj�,�m5�?�̚���L�յ�e۱AVOg2�t�Swƥ~=��櫢0�,��Xt�`���}��1�U���Vg8�A+�ve@VY?������z�6���}�sߪ���^�]R\��ņ��L>�7���2z\6T�__>铯R�Vn�צ6da���ֹj�g�X�y(6�g�>��Xu��@��[TY�H��MVH��kC��N=`���WK�0�P�'��/�O��r�B�#ΰf	�^7s�JI�.Uf�/��5;K�w���%!�����e��������p�(��ϡ	V�Q,��ݓ�O�3������Q2��&�v���{S *��i$m��?`��h��:�Zc�ס��T��lT�����F_�z/e�Zɟ@�JI6��i�,���aH�~�%Yl��5〣sk�'�\W�I��@uS�M��nrUw�:j���b����ဲ�.2���1��y^�X���a����c)ւ�Ŋ�K`�n_,��@�Ӏ�w|gF���Ǧ3�!hX��1���tq�C@�r�{�=���='2�w�� ��Nsx*��9���:�!��ʟ(Q՛�7Y�R�$wkc��Uxx��Ǥvߴ_�����d�+?H���T�	������>i_쳀�ɶ�z�l�FXG� �%��GCGr�z���XO�5?��xB��}�N�.;�.R�:m����B���л��h���Y�}^.a��>!*o�j���q6T���X5�#�#�x�'��y��kn��-<���r�i��&m����"�W�~����=��	�IW�v7����a�ޑ��s�;م~�A���(�G�N9sq�:�=�i(V.��v�%��-u�S�&[՜׿S���AX��`༣㢷��eFt��F_�8�K{<@�l�ݕ	4x���@��!QR�猦&L�f�f�=�v�7|BH�N���Jzg��%O���?�F���t�	;��� t0�t���
��D�CyF  J�Ȅ�:ט�E��o��[�ͥu�i�uHp�Zi�����$�6E~��6FO�I��0zB޸���Y$i7%!
�Z�q8z�����a�'�6�v���g("�r�[�%B� �j9S/E��0�yX��	{T���y�g�[����SS3�q��PJ&K��n��}q��ek�ts�+g
����glua��y�}�J�k�m�����tEd�Τ��M�C�Z� D�����M���"���Q�g��� �p&��/��e����5S�j�l��J^��⦕Ql�h���J��~Qh��<�p":E���ڈLgGb�eb�`�=�ܻ3v(�/RC�<sI!R�v��[�b�M�Y�a�!�{>O�|���;d���"VSAꎄ$7�lAM-*�>��&Gc��
�
I�(�8Z�$13j؆��q�.�Lk/лB����5Ox�O��m򔭠5�%= ��g���`I�q�`Tp>H���|O�,Eo�FM����t0ۍ\[��^3�F!t7=McI�\h:d�n�M}'�}�>�4�����
�f�����F��{�������lR�Bc	�)@�Xu�'c<n��b ���'�Bl�`%�ȹ��T�p��N`���d�+��b+��e��r����E�k�^��G��9|��-C���IV�����K�Kї{�*�5S!\kl"Ykk�89�R�n������bS� �3����UmU�����)�@q�+���8����R�m�vZ�,EI$��	W�g>q��;��m��W����m4���M�Ha>n��Ȋ�����k�Xբ�H��Cx�4���z��t��xY��{��@�A��^�J�U�p �G��_�q��s��}}ҵ��~<�ӵ_�ӽ|9�"gn�D��Z��:9ߥ�#��JH�:3t��K�/�>W��5�5����*���p�Mh��q{�@��JE���;R�<R8�q
r#�@W�@ڔ}��,4}���Q�Z�R�+ V�M�n���6�fq��Ò2)J�9�����ק@9���ںc�'oԹ�C�d��9�)�y*�Ymdz�l�Ye]�}�7�to�`�Ӊ޶}
����y�i�$��ɱ�4;d���y敚6�xg�������GU��y�N�����u{��K9����FG��j�2�[���P-�Z{Ԋf�Q#����Ah5 !�o$0egi'�]��h�l��*Fe���%��P`BZ�Q�u�Pv2W��ģ���@�N�d!QW�p�D8�aS�f'�=��_{;a�c�q�@�5̚��U��K{A
�^^����m�>Y��[�[HJ�On5HTg���#Ab��'Lҥ�;v�4��Bsv�l����LF5���Eѵ����B\��x��Z��r
���W@�q	8��f���%$Bw�n�����*{D�ɕ@z���E�O�t/���i��	��$}���1�{Ge�A�s�1�����vH�~��rJ��F��,1Ɇ�e���A����ť�=p� +zޫ�B^��u��h���*~' p��;�3G�M�P���S���߱�T��;%K�x
צW��B+ A�eb%n�+'���P֐B��O��f��r�ڮ��C��m0UZyz�"߅3D�kb�U"�Q�w�\��he,V��Q4I2��
`�tKP�
vN0�4���BЯL���'.=�;|ǝ�U4��0S�r��9zkY�,Jp"��{��O�s/�`| �1  ��%]�ݶz!D�Nm�	����}�_Y{U'�����B�"�Q�/&���^"���u1�4�N�`��xvL_�)
�b{hӾ�x�m� ���� ^v�4����y����2K��{�!�"�J(�.l�I7�#���,��=P��o �9�8��)��TK��8�i_/d�C��e\�q&��.�9!�-
���=m�W3k˄Q�@?��8X.n��xB>|������Q��?���k�Ɋ7�PN]�#9�_������?�ӾwL�&��tΠ�x��������c���k2-��t�㤊�j�If`WzI�	m"CC�øJ��ӵ���QY��*�Yr��j6>�(�\b����g��r��O%u��»�n@���G��(G�C[�)�K��2B3�eܢ��ws&;���>�@�S+y�O��̉�෪f�K��A*�1��g#��̯���^^�`�P
��	��˫>�-Tbr��t2�>!�@D��r���j�K��h���}_�1l�u7A��k��Y��}=��7R�&�A<�"���G#��M�@�3H����dg�������=��$��-�Lh	��A��~�B�)�u-��{�U>b���>.~�8�T@s�E��vQ ��؈Z������N�;��0.֨�O�nѡ���6_�7|�4�4���-J�h�B���ݞ>>aPu͢��;O���5�C0$o��ƈ�!���ܩ����y(`��G[u���M8��5�j���s/��f�2w|��iuS�M�gF~C5Buu�ǎYƪ~�,f5���L̒ڹSIY��
\%x�����?�G9_�ڥ�#=��H?��a��Qʭ�GV���K���u{��2~Ų:�;�T����(M�p�7w���S�L�=tHMC��.Y<s����N�,���)3��vR�r�VK��b_����5�+DC��i����s\h�D�4�*h��QK��n o`�re�+[;6��:�f*�aB�kV�7�Ќ������_!o�r���ݨ�<��=�zǢ)�	���c$+@�K�9�xbA�榘�C�k��,muMt�	lx@Rt��t��M�4�'�!��W�B�K��unZ��u:���A�o�k����+&��U��SPn�Ds�ؓZ���v�cx$i��"=gO�.e�$؏2�^0^2��
��ES��������d�]V�'#�e���zfU�A������B`��S����^��!�H���Y��#^4~$c{�bW�4����GT�Q�R7�Y��]�ub.�أh=1�y���K"nʰk��[{ebj�8ۢ��Z��:��w^i�j%ȴ{UT����ʥ�>Tm���N�Z�q?�j-!��Ù���w{�A2Q���,��2?*	�f���l�tU3�2�cs�� pr2�}z4H�e�2��>70�w^�< w0=��G�1*�t����η~�Kis����_m�W��:�}�乑���+J|R�;e���?��䗏P����O�ˮ*�љ:�SQ���	�[%^P���i�!^���=�lrA��ATGG$=<v1�P��		S�!$0EʙSq�hvi\Kv��3b-W��kG|����m�8�"��B��)mq�j\�p+씝K��Ğ`U31$A��'_R��v�ZdV����8v�6�h��%	���H6*[�o��t1V$����O�����h:{����5TI���9br���0��!��|�Т����Ybd#�53�����̮:���'�3��UQ�'�*N	��5�(�PP�s��O`V�XJT�ӱ���C,��.,�3�|�y������	<j؈Rz����'���J.���_:�C�{�gȟ
�D<���`.�{5\�O�O�9M��F3#�ъ��.����D�#��8��{���\f�.��y��Z�>��,[ aU���t ~Wt�����p��CC���Ll�o02�����-���z;�_�r������D���Í�JF`�b��/�_�}��D���~``�O��(��u�z�U1�I baA�o���P���m6��6��5-h�9�Ff�רj	�8�ں��7�t=��9o8Q���
Գ���[^��z�0ڹ� ���i�deӫ*���/�8�y�Ϋ}[7��Y����\uJ�l}0�$�?��4ŷ�&.�t���qJ��{(�̳�Xw��\����B�ӷ��މN�5CTw�Ċ���������~�\j�у��.nί�.a(TB���ƝKu�;����a�Rئ9G���<�&GL�!5�a?u�G��#�w��u8Mh�M�al,��e������������	�ר����£�.�o� ��T��ֆ���W�k&ǹ�E�gL���;��u��2��(�IW���Q����ٿ�Z�z�Ŋ5[������&��C��H�O����K�$]�j���2�V�	�챍
J<}-m�"�.�l,��ұNd��,��Q%(�
�B}�P���X�FUgo8�빾o�����"���p�,}]��3w@ש���k4�o�nP��8
�����f>��c�}���,��F(�l�(��!���?b�$Q�}���v�}D�h�
�6H��#h����R������ֻ01o��i��HZhz�+������
�#��5����k��M��ߛVUa���O|C�a©��O���X��RJ��h��"f������f�A�%쎾\��'��%�#��|fX�)�1�~������E����d��^�Q�:l��	���3�<����?m��t�=O�{��I��ۻ.��2S^�f��P��wcCKGٖC%��l�~zS"\�Yk�Y�!E�Ӳ� zYŏ����	����leI��|�_)쀆��Ž�;��MfO-'��	��3<���V�g�Q�)#���U�kU:�L5���	��E�9��#�ۛf �bÅ��ǅ�rXIp�-Ç���<�2�c�gP	×���A����R��1_�`֦ޢF�\�p�p�0��Tg�P���|�qŨ�zy�͔�K�Vc&
�o29Uv��6u@ޅ�%� ��g��!9�VT���U �b��jd���g�Ծx���Z�
��a$�g".�'�`&�;��a	C[/R���� �]٨��(N9U.WF��;ֹ\d�!$ *��XN�b�w@��u P�s���y���IL;Qʘ����x "�󡥋��E�Z������GMV�u��ao��8	����D���Q�a�3�X[oܗ�ɿ�i/m�%g�c_�������'9|�U�T��ڐ��|H��7l\��¯��{t�uظ�I��8�K9�O�μ�%���������6l;`m*ܝ��%>:���$��i���3kgF��e�-W&�2!�U1:O��rY�rt���-c�����7��1(�*���C�z',�K�����?��T��x!�֏��GN��ӤQFYGlS��$o�6���L�=}J��p.�� ��ѷ ����t_�8MJ�>�a1����.�3�n-\C+�5�V3@�E3о#n�C�R�	n�Y?�ܕE�k�	�k���XՁVo��X���ۙ*���q���m�.�8Y�)�t;D�*JFFMZ��#P��zK���2��W��;E��4Jv��ٍBq�1+av�=�0�UOS��_���u1@�O��.I��~�R�?��.Ja�A����*��K^Cu���sO,~� 0g�7Tߤ���̤n����5)�5��bl�L;�3��#�S�I� Ҿg����p�� �)�QbȤ��bx�o����* Xu>��B����^x#��c�Hn1�<��G
���i�.Y��x������NGk�`FDB��v�]8�c��Ћxj!�I�la`~\������wWp��pMMd��� iz��7{T�u�=�e&?�,ίI��ޖhÇ\�W��!�SDu}���E6��Rq��"dH��
�^�-JB�	^�BD�d�%� �t�V�^�wT<�����ȣU: 
��:@v���).Eݳږ� ^؛󑼙�'	U�Yt�����p(g%=Q���_;��|CRvD9Q�A<!n�K�u�LͲ7�U�B<��HR�,�{(�'���	I	�&u��暗�րv+y��I&��!��&��vc�(�vb����Ddw�Kxߞ����n�F��#���|r��T�}�1�cbf������]D��q�A%�Zj�y:iB=��	�Vqe����K��D�/ݚ�Kp�#�!���`��]��*'��Q-;D7��z>�nO�*���<�)@�y��C���H���v�����/��$Tc�	T�Ui4�kMj9�������E�F��%FI��HhSZ-N��bz�)響�?i�薣ZS��D�1�Ez��N \��NeO�2$�$+Qb2ZS�Lb��,Rp���`���>��Ne���h��Y�_#�W�itPLlbQ����H%�g�0c��n>�4Ȱr}��,B��Vqs�7����	��;C�^��ڗ��y�QӋ�cV�
�s�ʯ4 ,��h��{1�"oj�t���b��f"�u���{��F|}�U��6�kg��|�{�����5������hT�:���0�擄8_tL��j������:~� �J�))3�չ�j���v3(0<Yd%>�%h�]�aM��k�i�9C 5�PX��W@�[:�6=
;�n(����⨯�<k�F�t��z�]
�(G>�	��_�*�ZG��ﴲ|_����e����Z�]�z�#da�13H�� n���C����\�L����`-W�sA
:��k� b���W��k�۱�~s.��2l����9�`I�Hnob�C�/��A�nz�I��?�5�3F����[�U�}q=��ğ$ �p{7�Ȱ~�K����<��%����f�o�a�r��S��T��oO�N���D�S=�w�S33n$S���VIHs��=�@a�=�����};�����}HW���eio˪t��X�	�N8Ɓ3�J_k�]�M槨��.����\����͞���u�(F��Thy���m�W�OxWb�"[Dbc��ȉ�#���e>Ƅ�p8o��З_ ���Ĥٚ��=������t,K9R6Q�N�Tņ�nsk����
�
9�+�Pz�V:��j���	�u��xhd6�5���� �����c�������u�E���������v\ɷ-{������� �sW^Wɍ�E�i,��bo:ެ��F1+�d��O��9��CL���-HE'�R�cQ@�&��L�:˥��{ip^���l ށ���c��PS�ҡi9�s�:d��>h*��5���'�5AfA�sCX�*m&U�-�2�e� ��^wmhxm��u�Z�(�x��嬟9d��F��������}����I'7��8���mXh/`cO��B����ڵ�K�|2V5c�ax�D!�ٕm֚���E���!F��P�O��)弃\Ic��+�Z��~��{�n�����\� oRN_�x�ٍ�UW;�7453��j..��9+�_-��XLʘ33{%i��y4�8�H6���<�^�~"ȱ�x������͌�NPڬ��$��Dl"U,���*��ƴk����k���fė*
0W@bS��\�@4��pX��]���)Կ�샷��e[I�÷۫��[ψ���.�R���֔�Ҳ�o�c�f�Y�Tq6�9��]pKN-�.�N<�Z�ٗ�j�c7;�6�J������!,��>~α�9�O���9s�ʢ�D��fs)�aS��>���љ�B�݋#��(Ψ˷4�UB�q��}9"��ف��Y�r掠�ðy���Ho��=^��u~�6�\���C,�!9���X����� JnG�V�:�J6Q���|߉P��!.�>PԖo�|�����C6��<{jl�������u��æ��>L*[��n�d�i563��:�N3a��AHOM�bt�	��ug3���0@� A!Y�+$� �8A�!A���\�����{Sx��%�c1��S�I���:����U�*h&T�9;:n�/��z��n��kuaեk�P���6<_Z�C_��5��vP��
�Z>�V�y���!�<�R�Z�xL�B�40���?JK/�$d�_B@-�f���̭O��rBd���i�C�T#Q�|����hlW�q�W��	D(zDN��jL�:s�w�;�0�-�[h������C&����c��������:.9���Ȍs��3�rW�Y�m��f��Qy��:E���*\��,&�M�t1	S��%%4�5BP*^������8k���&ؒ�`:���$��RV!���n��q�Tc��*
�%r��dC����B��3|�d�8�ㇺ���.6�<�B
{��rxgX��=O�J��|?�­ɟH��C�'9�#ǃ�������m@6A<[*%�YI���'�]���:�����/<��59��%L 7	<K�}�r�hȢ�����!�9��W�o�X����ω����cr("%���
V��⥄ijNvI�����y�������`�����.x��jX:}����AS�PP�(������N��B�X�-uJ�s��y��@�u���o֛�='��1�."R�?�>�I��P��b�����vŌ��g息C#�Q��T7��;w��C�IQ�jqA��)^�LMْؙ_��T,���݋��꟒^�V��F�ʞՖ�biWEzirk�����3���/����a��"�-�? �#�d`���s�n{��3��"���[?��k>�]wo�넼����K�,�w��s�.��/�y���Kx�]���<��z�$ $Q5�̦�,�Fb��	�8�~����GC��_W����ԁ���ڿ��$�Ӝ�nm'm�`@�z�@�kB�+��H��5�"92���_��h��%�^Æ.>^a<W�v�g7��vh�"a�Z��1����⫁�ڣ�(��Q�|	#�{�-���楶�Y�N�ɺ1�Q�VC@��P�06���-A�ݧ�1�k=,���Z ?��>��Q�S�МP?�nm(�����`�x������b��CB��B��w�[
�����\��lpaΊ����ʎ�g�]�g] �����\��xC�U.�sf������3{�b����5��E�W��C��O�*b�<f�'��I��↙�[�R����6�*$������^.��b�O�@���$�8��Om�Za-q�J86W�`���;�E@�yM���U��7�\��je-�T����"���W���w�Ϊ'݈���%����lʡ_��񔂤�Z.w���.��q����e���;T����tO\TZ��'/��=:Pڻ�gS�����*[�4�	�*pd4xɤa"@�^ �F����IP�&s�A�H}>���aQ7���t�~�79ڎ���\8)��1�u^�4 y�Pͯ#��Łq)����r
gk����LȐ�y3#ɀ/�~�u��u���a�t�*Z��h��0V{�8�!~ot��W9������p��jO�3�J���N�f�*�8���n+����XA�U4�-����!h����@MŻ�-��/���I�x�G�� ��^��<��b�Ѫ��"���w���7"������7x���V�p�S�S%U�6$�|=;� \R-�Q7f�w�#Z-X9�y�[2u�!���)�QL���4'����a!�.�����Y���P��w0�C&��ְ^߉Y�ەom�ĺ�/���=�
aD�)|����3��	�����D�����p�<1>�Z�I�DR�ʘ<
l����A�o������+�;%m�i&�Ί�$Xӎ6�I��]I�V����z��}�i��Q%9\��:�~/���d��D�_�hn'�-�frZ�XW�� p�_���My�x�7.�)���R��%$1-�l�;w�8��6Y��잿X��x��+�(�mzn�S��A�[�[��~u%P��4�z�t|)��d:`}���3D�`X�p/�;�2�O��2pV��;N"'n�ǣ^FG�C]<eH6��ʠ����Z���|��S]�����{n#S�wЎ��ra�Ȼ�ZC��������u`�l����] ����6��:`���Vȴ���y3B�۪4�Ѝ1��̅s�N������JO�����D��ُ�b�G�]JN��C_xm�ʔ}	�r�I���;�"pb�m%�,�g:��?{�S��6�����5�0��en���(^e�w��±���y�u�1-���:0�����-��3k����(j;-�+���0T=����,��|b�#�e�!r$P�3o|�k�T!�y�Ũ8�NWH��T��4n����Cǁ��׷D����;`����sp`��Y�jݥG�מ�ӡ)�`<��Y�0��0iʦU��}a���Tt�T�߂�W4a�p\Kc����y��	�,m}��X����2�W�&/���s2�- ��YϨY%��
=)�S��^JG�p�H"feH:���o��"aǄ�Ѳ
���������%�U�v�G������}�Er�N�i��~�qRI�d�ےn�8afh�t�3�ʘ�H÷�
r�@.:��6��
�`�j�d�y�~h�?^�V�-���c�.�FG�L���,�6�,���{�|^F��^u/E��O�T��6p��r��n���Ĳ21��a��w"<r��z��N�Iõ�$+6Π���#`|�ޯ g`F�������E�=�O�egԀcA����8���U�
�lw�Q9A 	��Φ�!u]s��l'�3�}��Y�X}���zc ̈́l��/d���K��A���!A��Qv��~ 7ˈ���2��eP3�}�h�1�k���Ļ�8����g�����Ռ�r&�TPR�\���k�� �@����`��mߕ������#ɺ��}O-��L'����s\�qk�)y�k���h/�IٯF�(���O��&���p���Wu$�����j���=I*�BD'P�IZ%���G�J�ꆥ"D6ON��<���*ի/�\_����҃��`l��p��x:~v/�����u���ET�,��x&/�iQE���X���a�� ˙����Zڭ?��&7֕-�ʐ�����dR���ȈU�z�Jw�6b�A��T<q峟��/W=	�EH��z"B �8CuOE_ � i���4�'�6/���Ą	�v��-7�h%a�~Q*��mV��f� Eb���
Mh�C;Q{5���6�r�7ĺ��'nˑؗ��X)@2���=��%�`W!�Iw����4F^D���$f�$Dw���'�W�K7�=�;���)�-a�芍YD��$w��Y3[z=uSnS �^#�[L�D�(�_'�w)���E�xl�)T䅞׀
��p@;����R�TM~�&�q[/R���}��3���]���n��R�]%�=F������;��f�ɟ`���f�c�+�t7)�,�e$m�FW��>����,���ç����C213��L�hai�ўs��J0����ziڧW�y*~m���&�����3�/x���2������}�B�gw�4k�o�J#[J[�+ ���;��D�=��d�QĹ��Ui|�%���ú�z/�ÝXh�������$��ܕ�d�G���uw����@%z�ݭ�ኀ��;Q�o^�ti,>
8+j(�f�D�5s���R`m1>���Y�̰*4���5F���?�.�d��E�Ω�Y8߅J�a?���N�q@(0*��S� ��Sn��W)3��Π�%"�"c7-l PR郷͈�>���s�'��%/�f�����?���>z-l�����$F���I�%��;�-~�Z!��j:�(��$av�e@X={���<�����܀ݘ�f��Ƴ�A���.��#t���kJrY;�rZ��o�v��yd,C?�f}��M�ȵ�Pg� m�|Ez�e��K����&X;�zCv�C��t,�JCP������MȂ��ܼ�������}�1�^��=�ސ�>��f��.lPQ,��u±s!�Jsj;��f�8�lV��!����I��bQ��E���c�"�o��a=��ҟ�j��Z�F��f����rc��$�)��я� � �l&+�7�)�>r�Y���7	Y9����I&��_�W�s��ǅɻF��w�}!<=�ᅆش��ΟcN�����!��N8;&eq6�(N,�'�UR0,�����Gg�����ϼa��9�O�A�82������(�3 �������3W�v����C?3�M,����)��A�"x�VѶdi�͓P�"�Q�у!Xbq��Q�ݸVF~��b�fJ�JZ�Z)">hl�|��mUi�f����#���[�n�lT�J;����smu� 
�ڱ�K���� �uLs��Q�@�0�V̱�Ը����T�G�ߝPS��g&����Vf�C��-C�М��w@g&�,���x����f-�|
U�&�-����AY|��P<+���I����:���F�v��s�4��OsME��Î _}�$����Ƿ��*%��%V����y.9ku�iZhy�U"���8�\�!�45ig�&&!�7)�qxH��d�Z�8���A/��%hW��`��ع3�i!�����xu�BN{9#jb�i�n�S,��y�A_�:�t���P��&��[7,r���J��x����0ŧ��Ԏ�w��ۖ]%�_�G�w�g@�g}' {$��tTw���(0/U�7��{��p�?����-�0'��p6r?��V��9<Y���,�0�ݲ~ApA����/KyL���w/��������U�o���%�#�Y����=B��+�/���5��������#ݴ���?��࣒�Qf��=��n�t�����>��ٺ��?�Zj��a6C��Wd|������jCxoX
� ܈������@�	�h���C�4����QL�@��K�5P	�Mچ���խ�w�V�z�c��/�\ASw��;�	)�<�L�ƕ;��,O~�lŃ��&P;��CS�f�uWc�ʑ��HC�	�@l�������,5��v��b4��y�%HY�a�*J���8���	߾WJ������g���&(fI�>%S�8r��������6򸺍�T��#{YkOX�D`2C�*�����^�5<1%�;sp� r��?���GY����|z)��y,���vz�O��� ���f��yڛ��܌|3�g���I%����ԏS=��:����P��a�c׿^[�xL6E���]�eA�� 1�͝��G�Q��H���΋��r�v�a�&�$���ўP�q�wm'#*|3y
�K~�ޜ�y�4���miH��_t U����V!�>Z�y��#\���w씬�}64.�/<�����O���q���&#̇�"�Y=b���*�� Z���81nF��[/�7U��S�F��]�_���E��C�� ��6�C�R��]ћ�-9������t��:��M��oO���?p�6�s��؈�<ݱ�̫����\���Y��2O	�0Bw����&T�������'��Jd��]w��'�[-j�i5B<+L���n ׊��.n�$%K>�:�خe�wBW�Fv�U �d�����
,�Q\Y��;8�ac���[�U�yp��HpfM� z�s����[l3k�"����8���B(T��>�UH�?�A��g��p=Ӵ�����Ӊ�s}|ѝ���t�:���?�[����s]�v�B�N/ݝ'z840�ms��PpV�kUN��.,s�Y��/�k����9�$��,�;��?��:��s|$��ʟ��h}lj��X�)qr����u�e���ݱ<�PH��x��X	T&��b�a��V�Q�{"�;T5`gpA��^*��%�V�7��E���/sFr�7u�X�k�(?����0�VZV�-]�
Tl[��a��'*�8�C����}=?ƦE�!��ńN�!eyU5���8{�QJ�&#>�Kbg��M�k�m܀�-H���O �nWW�l�#ƳO�CK����Z�n�m�����h"i�a�U�! O�K/�o<y	b�i�;��ٶ�<_	���==���W$�˟�u{�e�M]��u5�dp���>IW2r�+�6�u^�ң/y�c-X�h,M�1q]����a�`��J�;Q@��`����������")�%q|�k�^�ܪ�h+W��br6��E`�w]��{w�u�b2�~�u`uB��g9NAs�W#��e�Vl�i�a�i��x�΍�r��D�f�ii?Mb�?d7��RO��b��	���ݴ����2F�;��
?
����*��sc!�?��Nlzh�(�j�)�C�F}��U���_�� ݣ~��X �o��;S�ZLl������d��2��f��.���)���{R�e*��� _�g��q ��F�ײ����;Ҁ�T�xʆO2j�-��Q2xA��'�1�m>u�Ї����R��L���|G%��"fʍS�ז=���,P4O\!bB
Z�C+e�ÔĄ$�r���*k�e]��~�h��ƙ9�f	@�X#]Bw��#kl�D]��9��,xn�;d���C�^sA 	qF�B���/�;�������jƷ�F��t7ǌd�ߤ!e6EV;"�v@��ŎX!E�.�L�	cMe��i�vqg&Nچ�S�+���V��8�w��AO.W�Xuj�K�K!/O�*������B� �����&��qC�V�U!��VI��������c��S��^ɕ���%����BXT�u8SW)^+t��@{ĸ�:���bq��l%a�����N��H����Ǌ�hIDl�yT�Ԍ�Z��v�����,�P��=z���:
�%�+[	�M�L���hN�����&�g�\Y�mc�ќ���4���*���Y��o'(;S���Bx�B���aM�&h;b��.szY#�Y[���K�=����sH/Ʋ���ސt2�D�iJ��\��l�f+�Q-�9�9;��g{�]���ݩNJ0eJ����D���m�0D>�-�?�ǵYF����N��$^��Fխ�	l��z1����Zy)�@M���(8�m��qY�ax8�)��*�W�v�(���x��n��D���1#��x*34Y���	D9� ����R���.�~%,q�6u0Uٵ��H�t�	�zՎ�n�������h�~��ir�F� ��ߙ�\��e�U@ϑ!$!��Bdb%]ޭ�[����	�2�*9�U�G�jG=G�����jE|�sI�"ǐ\�`�S<pM���(+�R�� u �,x���lX��2��JQ��ls#R`^GB�`�Ӳ���
3х�ܶw�~��%���w��p&�
����R���@�Aj~h���ɉsX5,�3#�8�d����TZ�^ߕ���+^V�v{�tG�0�c�O�qVٌ���f[�[��Z���:�8�q�d�1�+��M��m����\昷�y7��c���O=1r��[.x�TR����A���p}w_<kMB��3`�m�����ӎw�^d+ȭz ����g̵�Vy[������V ���+","	�=��uO����x#���mdދVE�������sJ��X�'��07r���,.8�<9��tq��S����?�q� @��M��׊G�eL�ED�Gׅ��z�zzQ�y^x^$�}��"7�.��C:	]���?t��K��+׭gQR�a^��w6��e�z��8R��<u�ncyp9�����,�5���	��^Tv�}⡊��x�+O��L�KkHg-�ٹ4m������_����OپSB��R��.&8-�a�LPV:>��w�p�0A�F:�	JWM���[�Τ1�F�-��
fGǸh��)%��&{T����,��d�zP�$�v��l]�ȼ�MFn�q��s�	S�N��F�H�:,��ŅK��r����C����,d��Q�w�H��X�m5i!�7]Ma��G��ϥ����-���2��|m�69E���u8��~~؂��)����q8cT�u�zY��x�<��X-��v/�mQ}t(�Z� b�=z�E���1ïl����t��}��&D��η��k���H������hz���?�e���nc�uC��n��`Uzxg#V�IDe$!J�<D�_��	x����z_�9wn�3E;5}9<kn�i�m��ɀg�+�w�ч��1�奟9�� ��,;�ӻi}�͆^r��@���b���Y#C�_r-p�mP��g+�.�7z�m��sIRj��I�^����s)|��_�Ϡ%��;k�խ(��:Qqu���ۘ�,�B�i��DZ�8)����3u��2?>*�����Y)_u2Z�_���9���x�̙"8?#}�Cx�vl�s�لz����,������P�kBW)�"dh��K��Ȫ��S=H��GI�s���e���p�</����/��-�9[���<]w3V,M��b�jF��DŦ!i?�����m����O2C���kw�P�1?p��RZ{�fH0�(	d}8yI�P�����^ܳɜ�3lc{�=�Z�"�}���b��]�"�1O����o&��<c����'� �i�K�*��2:��!>�U�U��#g!o�K}�Hܧ��/`���n��ե����hH��3z>��-A�Q��o�FϥF���5!,g��v��t�0^�Z w�3���t� Oe	�8�'�8)a�Jv/#�ÂS��5�ʪ&��WČ��d�Z���L�'"��h$�Hh'���`���j���}��(+��OBdD�/����oBB�j�"����˥�\J,�z�t�w��sՏ�Y�s��v�81HBاr�W~x���vV�gfN�I��+��\~�2&78>۫v�������o~�r��������� �3�T�Z�;����;��VX����y<,���S��m��G����Q6S_�6&-̸���S���q���-F�k������E�waT����v�3��2�jo��%���Y:�.X	�1s"��n��%ʽh$fZu�Y�K�>���?�l��r�Q��m����V�K�	y'2-��Z���^.��ݝQ�|���k�M��ƌr�r+���/����9����v�Ѵ}75Z�3c�Uh˚o�� �A�|=�l�ߎ��9y���ƛ A�|���� H�2|�b�58��L58�%[�Iot9��K!��}1쯇��--�[ò<�z�rE�Z��L7�
�\�#s�c�ɮ�)���f8�ϔx�U�~��\�UH֯������ԏU���ナ�7�i�yeQzgQ
o�+���ᾞ`�����ԣ��~F'��5;qpr���Lp�+�T�v���if�"�mnC��c�����p��U��}2^�P�.�/EG|���>/V���T�Y�#��liQ��Ǝ0 ]y��J����Kxq�L��H�q�1�η]��s�x��e~'�4�)��/�ʮ??��*WeB(2�L<O��ך�c�ӊJ1�����d6R�}g5H������y<P?	8G��I������������P/=��IT�1��@��84���U�t��4����/)
90��֗��R
�?���0"�.���ً�kE��[�p�?� �-m��$�I2���k�m��8L��M8�Iԥa>l������B�C���m܉� �����Yl�>�x�ޜv����>Tq�֬���#����;�����k����׵��(xT���%t�zb�Q4=�!�����V�/����BEGjf9b�	�)C���a^.
#qC��2rsL��?Hð�9��TH�i�mZ�K���v(8��5qO��X�	H�:)����ՂO-n���4�us��&��	F��N|���ID�qZ�t�5���55�� �/q����<�
Q�!e�'ТS����d���a��9����
1 ���٘��F�5�U�2'a�A+·�K�K�d��|���}b㙸�X���A��!;�)�?��"�v�N��z�׋i��/F	�A��+�Q����38O�ղ��~�z/�.@}&/�����������f����
��0~�֐ȋ����~�s�\S���h��r��{xO ��Ai��:z��Ț��L}�}|g9�am���K�֑��uy�'i�Ay����1�P/�O��a�U1䍋�Q{��~��0(G��'AAV}�4we
P �c�*ŨL�� �8T@���i����H-�1B��$�!I�7�|_NhypH��s�IÒ�C���1B�bV�K�]��ϟ�t�
���J(xjzH'�Uw�4
�;���������W���i�a��첨���ޖ[�\�4 �IޗK-�/o�p��
���=��GՔ�Nk{��|���R�����!v����K��E���n5��:z/��_N����3�?\��ؘ�-"����Q�y�M0�t���E���������%:$����T�I�#�#@tLʔV;u��h �����?M��trN� c��	¨�I�Ƣ��K
�p >���E~�a�l��qg�?��㧳۬e���x�%���؛֯ۉy��r��1��,��_$o��_���$���Q�4�1�w�,r�>������k�L*jU~�_��Ł�-���-�D�(����0*~�Рh8���%�"}�}�$�W�H�z���PCއ4~"�/�Q�&���R�ќ�E��ۧ`rF��B���pq;�%���>�!M}xq/[�F]
B]T�^���⡸�l���}�~�{hV��-���i�ov�>��wB �z�,��r�4��љ�C5�7��`9��a��>2�Κ_�r%�QWO7�̲�'�n�a୴�5i�9Y��q�蒡� ��䓣c���vu�D_�OE�a�����{�����ʊ[��:�r�$�����<9�h햣��t<GK�%�z!�{'9�&cm��}T�B蹷���=�t[�fdw�D�g�q�L�]�)�����}D�	��}%�Ќ
�Y�X�%l�����W�ݦ�lw˷I0}X'G6�\����,�c{���j<.��|�!f��Ȱ��S�߾1�Ԝ��g�?ԙ���T/GfZ(^�ȇ
�+η����VC�f�����	}����~ۙGrݘ}��$�#��HYB�$��8��L��
�N ?�`�㞉P���
���<�N���|r;n�V���"G�&]�!a&�"T�C�#P&�jX,�(��@1Iȥ�[��<�3t@�����5�
w��/��}��b8-�m�<�����gc�Qjj�<��$��k��^4�Wc�-�&��[�I~��wBz޵����Wj�Q�!��G�7��ģ)m<��k�*�-=ֽ��^Z�|�i,����zzi���u^%���Y1�T���cs.�0�h����H7=	�~��k?��Gp�UE��/q(�K�r4�[^n�uJ�06Is�+��s�8��Mۛ�A����1�V�M��j6(��e�Lk�V� 銌0' �L�ta���I�WEF�8�P)�a��>IJ�|��� ���w$�4^h�2p^��s�SdN�">I�G�k�����\���� �g)Go�O�d3/iޢ�&b��mE� :��N|V��#�wћ<j'��&O����r~�Ҙ��eX�Tl��Q�i��hR"F�\[����K_��]G�K �i�R�'k�&����KYJStW�o�<Hw� �ȓ+�%��G��cs�).o�\�D8�Xs���*�e�~����pZ��,�M�Ww��XT_#2�
�u��8��GC��׼N,N��P ��*3�&�9��~��W}Ҡ8�N���?xb�-���kta^�; ��cZ"�NeB׻�9N��7�,�F���:�����[�b�P甫�&�v �MB�;�q�{RU��'r7G�:��e��V��d���S'�J��x��̱��/#o��B��RK^�����v��C�&Z^'[I�f���Ē��D�u����`=+��ʨ&B��x�C&���%I%�*�R��gŷE���P�f���f���:�����k�lh���I�&�������6�wG�b��`�A�4[��	Ue���} P'�Q�;D�{g�\�Š�S�⩹]�-�50��RySw��y�M̇�y�&�8���#�Qjyѩ��`0�(ꭇ�s{�� �n��2u�u*Hd�^��w�_@�0�W��������Ec�����Uw��iT}�ԗ��r�q��k�G!c�`ݝ*vK~X8��z�H�=�p*��ԫ�l�d���.�gv�w����5���0��  ��I���U�Cp��k$_��7�"�Px�����Xw�pבE����Du#��"~�&��l-��x��(���g�$5�uaP����wdngC 
���<�(������ݩ�5����2p/Rcb�4�o��KJ�H<�C9:I��+���^0&m����U�C��@��*��F��7�ؗ)³A�$>�&��[��w�7F ��*9~��I;tsM���K{,�2�r��n�m���!O�P��Ԥ�S1�p���Is*Ճ�����+�yOa{�M�8�C	kb�D�/0��|0ן_�f�'�Ji�����\mNe�s��m�W�M������7'��/kUtf�UES��hT-�������m�̅q��K0�mn~"(#F4�3�.|��/�5��L$Cvk������/#��F"�auZ*���$�B_T=��p�e] ��Y��4��5�K�����xu:��F���5�ja7Q�Z(5��-��J�l�n ̄���	%�a�oֺ��>���7��m�6�օ�� Љ�f���p���w"w�-��n��=����*8�@�v(�`��m:���5~(^�ij�HZP����
�3��2���d;�	�냪������*��ok��<I��߳��[�N��$.���p��|��m/�t�Rռ.{�4�d�{ԣ2�3>x3��I���,��۪#o��K��MzSڠ��f3���ұ����f�[B�A�P{3�9��0�z�56�F��'<*�Ci�:��ؽ�D�����?'\�_Gp㵱��\����������O�r?k��B�e� �](���{�OZ�_��~�p�gb�&��Q~ׁs,��n\0(���o�'J'��(\���|Bk�>�iT�G�����!��^�.yc?��-�0\���|Ug$�;�ލ���G�s�#�������Y"lĲY�o`+#M��}�b���2��>�}	:��ȃ�~δj�3�0U0����S6m�?�.4ղ�;������Yt>��p�p?�Mrv9�s�{t�	������i�ZL�� G���yd
�i'���>{�+��q�2ٚo���O.��ym�l@Ϸ�����:[[�ؽ7mZ�VI*��|\
�i�w͛1�u��~G���[���V�A���@���%�1*P;^t4��������v!�,ci$a����Ѩ�a�oc�������\���v5�|R�:���Q$@�q���7_�T 䶛��SGR>���̚����E,5s(6���a�����E��F�������f8�׀� B{aJ��f�!X��`a��w`�3��<�a��1�͖�^;L�-m\��ޛ��e�������Nl�HF q�V�ܷʄy� {S��9
��+Ex��s�9�L�mQA��E��䔲�icw�������$�$1X,n~��(��l����	Z?�bK�����%�K+����!%� ����6��-�3�����>q+��gO��Jܣ�ᡟq�f����v��_�
%}f��s@Z��U�1 z5���ݡl�K�/�'���H�$;҂�}%v��2M<�؊�ڥ�٣!�\��n�r��')a"�&��)l
���cG\��qC��D�>��&�l��^F�'�
o6,�=A���V���q_5���B�@�z�&����YN�F��Ҽbq V)�t�k�YAbj�!�NF��+)Y���č������3�5�+S�A��m*��� y{o��P��`j�i2�O�;���K��.�xa��\cҬC�@ �â � ��Q�%�� ���D�j48�ۗ��E,%��Y��Gګ�p��Ko��q-ܾ�Q�\�h7r�o#ӵE�dԆ���-i���(�� ��%�N���5��Yt���҂c#�� ���� c�f���U����Rp�Jյ�#;Eh�
�� ^c|��qٍ;i�S���c���ʁ0�����X]�v�V3��x>-�+�����#��3U��63f��c�^�-������c�X�	�jw�a��A0!��wǥ�;H�y��oo6DIwvA�w�X��Vi��T��-Mt�_z�q���:)�`�� Bɜk����l�8b ��)U�UJZM]�2���竞8��u8�JhJ��"�K%o �`1��e��+����e�u��YC��()"�ʲ t��@���'��q=���U\K_s6�ߘ*'���a�A���U�+��ߔf��\}ƒ�/S9��T��3,���G	�<4"-ڴ�5��BL��r�/�S�s0i��}Y�mkXw6��j�9P��.ŧy�Ґ�X��t#0��$�37̜[I��%p����U���A���)p��T��o:��X��)y�diD* ����>��'���
��1Y���(Sp\J��.�*������u^iÖ�<or��F�V����M�T�(�0��Z�v(UG�I�J���=��Pқ���D/��Ҭ��3��`{�\]U"�td!��}��%m�i����Kȧf6|B�'�ӕDR�O�\JW�^�s� 1�9m��H7�(ȖP���wn�#��!z�N��99����HS�(�D�y� ��|���M�?�dSl#��Y�=<��BU�\muRԧ��Sb�M�V���JՂS�!h�|3�2lL��ߠ�^)6OED�g9ҩ�o}[�{Պ�@�Y^v���:��Ёo��@ګ/��H۫��H�d,�|��Lu�7:�;߹p���F�11⚭*g�5�;��wל�&v�3Z^�NY���H[��b܅�2�[5�Wfj>���Ԕ��b����^�2\�����Y#�J˄$]s�\1<p��{�	�J4[���wDo��z���Tf����ɼ:RT�t�::;k�Wg� �Ї�k�����E�靚,��������*iQ����Mgn�O��9خ��!�3�l�n�?��C"@9Fx��d4*Z�G��,��^��su�[��f�M��&��­o+��_t�(Fŉ�,���ھ7'uP;W}d]q���9�l����S%;��+J�n��N���Dh����BE8c�{nh1*Ҋ@3�=d�:m�������;'��Y����c3������ˊ�^j7Vi	����Fr"Cv�f��Lm��"0���(�D �6]�`q +wl�Q/7�.&���g"��pQ�q��:��U������Is+���@��V�R��\BL�1����X1��7��M9{;�d@�y�ƠE�a�׎���J8֞Pao�^�1�گ���:b�C�3<�|O�W���U��rD��D��)h~�>vP��fȉ|>�z���օ��y������'J���s�K��.�K��x¿�?ѐ� lS�`�RE��ᮇ�%�L����A�T©�$22+�ͩ���@ѣ(>�N��&Gb-.+�3h��x��j��ES��\�
D�Y	��v�O���{����������3����Vr��N��3��M���V�0գ]{Б_����a\����t�?�,buJt:����\�D����-���w��ٛ�� �/�q�d?ܜ�Y�iqGI;f�F�+��g��[��~�^�1d�O�,e�bnK������B!�����d֠�TaP�8��I�1�,?y�־�M�r~?����WD�{W���x|wL��*$;T��]R��*җK�`������2Ĵ��iU5�j���A��G��J���P}tpsW��4�a�v�8%�1�P�'��m#;�m
gy�v��+0�b�!Q��pٸ����v3#����h���GH~H'l������]�V��K�n�^4X��ZO(�/o������LHE�	�"`����V���'�xP܏���l�O�>��$���(��oz��V�/9i�H��;�Y<-�6݌�%x��O���)������TΌ��=iK��G�n�T[\���T�9&ȵ��={؍�`^[�n�� �������I��ӻ�j_7�{��ZU@��"HTq�fT[��8י������#}>*Lv�D�)ˠw��)��Ɛ�����6T�L��g�'l�T���0m����9��#G�#��,M5p��0�Ķ�ug�a��ݩ�N5��A�e
y��313X ��y}iC&-���%X�|�NP\��A5_ �o����,���;���Uo����d��m����Eid�*��ʶ������jf3}���{��7�8�c�F��Ό�*(��O�N'���r�j����`Vr`EX�4�>�Ҟ�Ĝ��Um����90.w�ໂ�swl5�u�PyN�_4�����{�i�N���B0�Ww��$U�n�*�q����$@#�F(�����w.�N�������]���&|�@4�aB)�����)��7gJ�6�nY�6����Lw�:X��"��b?�v�m�T7e�cؽ�}~��J;>����D˖t��h}��hO�c·���N;�H��Z� u7�E��D�L[۞c(����K l��كV�R=�CY���w�Bjg����:�\{2�Qa6P,�	��5(���6�?3qx����!i��Bڴ:����������5nb���`�/,v��������-��2��~���o��i�`�;Tp�W�eC��P��]-D�����lm��uN��	\����6_ �����;R&X4W5����~�,eߙ��"����E��5�ЌP+���>.~E�iUA3��ٙ�����9��G�4<�r�ľ�^�al�~%D��j���j�D�j�ā���>�7�ôRO�l�`����2�l����a�{�}q���R�"|5;9�c@ؑ]��I8���˦(v=&3"�ep���\����&=�ӆ-Ą�]��x�b=Phf_�Y������c{Kz��p�Fi_�h��0<��G�_-I��B��#^�Je#�Pt�߄��Ug��wؔ'|-�	��ȧ �ɘ�ԍ���GL��$'ǒ��~\�!���M��Z�m���%�٦q���H�i�̧�c�u�d�V%�#��t!��(�h(�`XB���K��gAX��͵jpd���G��8�MY͕�4$T�+r�d-�
2�'6�c�����X��_;_a��(O��nם*�j��}�>�ĀS+F.�*
M��������~�/�L��h�'�흻KQ[��7��'������;{�g [��:�Kf�q����?�!�2���V�����I�e��:��*���A&�_)d\��¾�`|�)������q�"�QG���x��5z�{̫�Ŗc��|��m��n
���5r1v)���lEz�>T?��,�N�(���]A�-^���(!|uC�'�-��qD��P�.�����8�̖�M8�5�@�N؟�s@.{nR�~�[@�|ᰦ��c��*ŜK�Jj���&՞������e���ugȟͣ��l��7�k��XS5�*0+fgK�Q�|���'�޾����������ۜ�j�↢*�)�����>�]@bYd<C��k� &�:#X�7��7�4�9wv�Ik��gYFS	�'��c�D�w�����w8ǔ����/C��&��y?L+�,�%4�n�'u�����)��.��RS	�6���l��X<��=� Ƞ:L(s��Vgca'��/����Z�`�?M����A��鞃.�����{Q=�-�����,�D���3-)��VE���=R�!��F�U$�?x�K�(�9U�6E��~���m��"�j�\���Gof��.����a�CIvj��^;�Q- �}�9>���ͱAL�ؘ���x�W?����lx��UOQ�Zw�1yS���k�*�_w�R %;I��]��	����m��:q��3w*��5ޑ����`�������6ѹdҟ
�WA�`�tV94��:@sF��~��WK%Ra�Ms�'qg܇km�p��\N� ���x:��b�K�%�Q,#�e�%���<�`h�5�c�N��.�����4�LR��P�M.y�/�Ç�Ҹ�����)�+W."b[��?�k��;� �{J$G�ƴR��;-�9�($ᓄ0ߢ)��j�k��I��ɘt��H���y\�c��r��B^�"�"aW�A��ցB�|�g|)]f�S��G)�<��˅}����*���c�&���U>I�\y�_  K%"�����tmP�7<1]oh�H%7�fR\�F�<��ĩ{�yk~�c��h�noe�'��|�xv�D�Ѿ�
��=(�8�E�a(M���1���?\{q5��>6��%A���o��d�������d�Ǫ���#2C�0�g�p!{���G���Ŷן۩��`��+G8~,݋��s9L(R�g�����/jBx�$e����{��J�Z�h2���f��]�-�4���;V�b_�h��"�_����8�l$�ÿ�2P&��|;>�er8�5!j��z�]t�1�4��{/E����
�m՗�N8~�~
J�L��a<�����ˁ��C������	�Ϭ �3�֪�sc��-�W�K����d܄�v�"T��]��X,�0�'�����%��8|���w�q[��͇$��Y0C�*�*��R�� z����X�p��i6�н_5ٗ�(n"U%o����n�>�!G���tx���E���l�7S@��GWc׳�=��T5x���-��f��Vv52p��\��w�5��+�v庮�ͫ��"�t�<i7�F�|)ȩ#�l6![�`\'��S8���@�G���=���C鱞��ϲdS�����Eh<%����5�,�����/����]��xC��g2�.Alʮa#�����U�ƺ���,��?R�/c'Е;;`1b��uQM"Ę����ݽ�����~.$��R)5C6���ړs�`*s�|֫O7���� ���b��i�oɤ���j^�%#�S+yIm2a�_�#b?�Ea�4���CJʿ�����:�3�����=�º���ӫ�E�?�O^|�~ ��ϼ�������z�'8���ւ*�є"����V���o�F�ʧ0���a2���!w���F>�8Y��+�,0|{�X
`�2oͫ~w����\1c5ޜ /8�<a@(��G������x]٦�D����4��V��Y��{%����I��Y����q�X�[��
�SX1s~V)��>el�b$t-������x��+��ٻMZ.������n�Ʀ�p����H�� _C�'n��M�)�K໅����#�N����R�6�#y�]��0Ʉ	��״�N���!�x�@p�&T�{�k�?0�U�$ ��ñ�`Nh���0|֣����"l	���r>�w��U����+Av��	pF��S5�qT�e��W��x!�R���y�v|t��߬�q��I�0Bm:�*̤P�d����2��4�o)z�q�&�(��?Be�ס���1o��]H��Ty���G��A�z:���P2�k�L���ʻ�0;J��ΰ�1h�I�)<�#g��q�j۞BR�	��\�]B6�%�7��k׻1�{�pl�ѵ+���9���p�����~+)&�E�]/�IT(��,B� u���T��d�2�řc���{�Q�n�pi�Y���&�_5���K3GB�W��w?!єP�u�X^�����u1�0NԼ$ٻf�����Vy�h�4�T!�^ڦ)!� ��]����b���n�x^:
s�vW܊I;Y�u�Y��x�;˱ƎyK��̥s��a$��/8~������U, �}�s��Mv�����~����,f�Di�WRrHn�z��rh�i����4�jB��)b�x��	΁_�R�
���2�����h�5��H����#��d�|K�����k�6�~:ӻz�͖.���-9��m�"4YM�u�QL������L0�$���
��L|߄�fX}H3�R��c�?R�P;E�N¼@�SF�9-5��O�e�z	�d%|(��ks�\�aE�`s�xv_�3�f#�"�vf�[�v�KW�
r�D(�0��T�TȞ?�fU/Lc-�)Ya"��sQ��T�fQ�R��#��Aq/w`2�|U�N�9h�B���r�&������4r�>v�Fp�����@��� _xW�Yc�����}�L�y�S�(!��g��{��l򨒼����#P��z��������;c�Ƿ餗n�"��!�lo�p�'*���V��#�hP�;dٝ�$κ�������k� T,���^����0�ʻ\ӷ�Yӻ�#�I>��͈[���Z�E��"�D�m��g���ɀ��|k����eӣ��<L��E]1�`V
D����9x#kMo�UR�<fZ�4	+�t	����7�!�n��/�9.��T6�OV݋��d�XDV��Lk7����Bp�O&�.��D2}$Z���2���'�ʘH�6:ǁt�R��>5*�v�7d^̜�$�ЬD`u�W
|��G�q(�B�$����@�o;"8�_냹T�+X��#�q>"�p�fjvn��f�>�u�tq�߭�����,�s������ 5}\4/�*F��Ux�!��T/�h!�,��&��? ���wvP�Z���k��𙷹�`e���3[�5M����r�ජ>YWJ�%�]��̦����sd��^Q�@A�5j��~$I����,_@�ܱ?4&
r�-���4�����AwJ@|�F��׽ݗ/I�!!���O-�.y_]`V���]̤�k�=�PK�A����ݏ��S���|��>ocb�
�}w�����0�K��?�a��� ^{�#�<)/�X
!�H�Fq����	��z���_6r��^���B��H��|K���	��s1�;��S���Oǽ%�T�I�}zB�E���^=l��L�>�2�M�t�L�\�]���O�M]>u��@�����	��+r�Nl�Ӓ�`��o�eB����؅�	312����?��V��4$��u�g�v�*���h�Ǡ/���Iآz� .�a�g�K�z�h뷇g��,���ɨڿTz��bߒ4k���)��
@!җ*ܚ��ı��%EJ�O۞��cx����@�֟�6�a ՞d�王| ,"U��l����'����r���6?����h{%E���� ��ѿˎ���0
�]Aoe:@jJ���C#�b,2�C�i����Z�j6�$p����[ŸX��!�0�� �W~%�C�Ѭ���w ���l3S>�A�$!]ȳ�ׇ���$T�	'	��x%�o��/�B�_������x�Ƃ�_sE�L�����4?�h�CB9$����`�����7��J���J��1�@� ta �z%R�Ӧ��C��L*]lF�8��it�ن��>���%�+d��Gz[����#�意E6D�D��e�X��:b9)�c��3�G��`��g�������G����ȡ<#�B����O)F���Hl�j#���E�ܙ�YGh#wE��i�-�G�)����/��+e��b�����_�h�ۧ �VU��r��:�]��3���������}�]��U�\`R'=����ׅ�5׏���k�@���/��h�B'#����]�	N	i4�h>�$�_ּĹ�n����,�4R|X���S�m�����zQy���ӛ�Y�QA�yL*»�cfM���e���y<i	)�(���6x�����$�P�٤���C�w=&�0��\j�r�Sbb_�˯�p7b�i{SW��K6��Rn�u�5E�X�v���J�]l5��f
LPn�NPh�Y�_�t�Z�����j�f���d�yѣ�,��`w]E#�]�;7�.y�����l�ŧ]�IH�}�#���s�83��ɚU��b�E��p�Dhړ�`�n�f�@��'��`�L��OΜ��c�͘�R�kŉT5Z��)���u�I,
ԍ�
��$��Sm�}^���)���y����3b?���w��MCL` ��f<B�D�1�H^�����ǡ��u�L��u��e��y�L�7d[���V��iY*:}�ѭ�f��K�(�$,�	�����gKy��|�8Ku�-�v?���Qg辚�5�;&"[�����Y��@����.V���0	�Y'}&��� �Ф��.k0����$�l�<�%�3��w(�����l�a�L��M%隨�r�ur��5�U�<�!�<��� 8ȼ��6�P�-�$2��3�S3"�lu(ٵ�����51l1z	�pƤ�5!�������%����&���'K��iZ� y�Uu�i�;�+��g�sMr��Ɉyf�b�7~��|��-ż�����n���T��G�>��q��s��0ζ��k���Ĥ��X(�C�W@�<�_YS�����L��RϦ3�=�E�ѼO��ep+�K��X|�f�G��]�	�/��*������Ӎ����6�m�8@���~�+�_���A��2���\\s׎��&m!J`�H��N�7��q$i6���B��siȩj����Dw̪���f*��IݲnFL"�,hyO@�My:�	��.����#���#J#w�Ʌ���K� �P> �؃�&F����>�|�jT+���zꄲ�߶�oUR����n���$��F �_�0�hD5R���`�C�������������Br�4�=��1������&Cr��<nf��D�b��Ŀ�"��fy�M~��&W_�W��iy|z���1��ݪ"��7��6QYc,D���V��ڥ�d\h�M�)6�i�>i��r!�N���F�b��[��}������NC��b<ǅ�Ԇ��V�ؒ��;��ڕGe�pP@��u*Kʕ�x�ʔ�
(r$�Z�QDa�K����D�f�V�ѱ�O�l&�?t���������s�ɾ$8{�>�-�ۑ��x��;bE���HC�\�i���Q�&%Y�2�w�Ԋ%ƹ³r,l�H{����Gk���*������H���.?�wj��Q��1���0pK�ب�ۃer/�_�ɷ�}����Q�;M�n�e܀u�~Vb0���7S$~���>j
,����[�Z��'�:�[�����ƴ�u�7�z�K81$��[��ܡ�~l�2}cS���>�W7q�C6����ဌM(�q�P�Kst��vm!w���s�~����E���_<�mk��q���Y�?W�Zi�.�.��.K���n�G;�G`�T�^�B�G>��Я��r�"z�J�+d�nJ�4q��Fi�O�0���h�dU�r����M8���]�:�ZKC�#~3*���Ԧ�5��ᬍ�$4#�i��>�D�]��������B�Ul���,ZA���8�X�;���?P�՛�w��ҁ���)���A�|���Ja�V��%[a:i��C"�Z��G��=���[�λ=Ck��L�O��Wn#�:	�c��/�ʺ��ӵs�1ͯV�0�VC?��R��9��q��X,h�F��� ���p*=��=��}�����<��,PG���4�Pd|m4B\������E��>�ڭ��K9Nq�N�%.���^�����՛�����~a��E Yb�:�鮊�Lfq6Ld�E�%�s�y�ޥd_B�C�%X#МXy �k����8�#t6��ﻎ���~;�&/<E.����N����΀��Mzd� ���h�\ƽ}���0�3�=V��X>_55��)"P�箯��cEPn����/¤�45���<��ml���j(��1�>�0�R�����Q����=���ӹ�g`%B��]�}��c���+ebTVϧލb+'�d�-\�����tW:}-��+�B[�ʫm"�$d�m(4�F� =���균L�/�1@��wS�v$q ����Y8�?H�t�ŉ�C�W�L�0��
X�q������S�L���� ZaJ��XC6��8�潒��#[ E>GV(�{c���1�����)�gpH����Y��!(��67_�QyP�v,7<��G!�3R;�")�GQ�I;����w� ����o�fŢ5h����.��7i��@f�{h�5��g}�=�dG��d�7ۺ�{��o��z���;�&�Yz

<�;�A#f�)5���d�������6�
E(�Su 
���/Ҥ\�����:@ ��u7<R3����N�P�So��MJ2,m	�S�1ء�Zuv��t�]EZ�J��}�	C�F�R��[�u~���� �4��q����̦6MA�ܖ�!U=�5K��c�7�@;��v��C�rG�sQW
tPҕ�[Ή�
$��⻍sXwĴ�<�5�l.��y�k�i��]���6#�϶ANb������\I�s-yd<mz<4��,�lR��^�s~DZ�,qxC������a����q�H�_X�
S��SJ���V������]�-<��ٿ�VWbk�������V��\���`����ｍ�l�&3�)��Ӱ�MN�
��V�RU��rP�p�!�ʖ\"ҙ=��>��.x���<K1oXs3��q�-x�3�8C�lZ>2���c�3�`/j��+@!`_���:t ������3�~���HE|#�R1��4�QM?�d�9�x�6�����l��J��jZ@x��fӿ� �2W����EA�c����?xcY���dw <���ݳ�+8��
G��o�y���Ix6\�QQ��r�,h����jEH(��*sæ�/�ĄȾ}z	3/�r.�i�80�ij:h�۽�&��tt�����m:���5���䢡(GX�ur��vC��HB_�n�%���ϊs>�kp�$G�[�{7sd�E�Aϣ�24�p�G �l�ց��dr�� tZϓw�3�!' �����l��gm#�`E�MjuǞ��IvHL9J , �`G��t��1ˊ�m}ՒA���;��Z7���:nB�4�^Bv<��ڗ����l�ib���M�E�t���bVRi��W�R6J�$e�!fUH���U�ůp�ժ�Z�
�I��`��m�o��ٱ����ޘѐ�z%����K���4<��t(��U̩�žQyG�WOE�O��ݖUd}��O���8w�l#���|r���¶p����\6�V�?G���J��)A�1���'�"�d$��;��p���~�k�R����+��>wN������8�Vo�w�o��!5;� �K�_�Ul ��Zi[>�N(�������V�ij�k�������J�<X��}�e6�C}�|�n�E�^XU��/�v�-� C�R�����1�m��Ko����Y��g������ػD�S2�(�DɫF�kM���ZF��U�!�|����_	W]��hq���"��KC�S<^h���BK��B��E���'Yy���+�@'��������m(Zs����>*��fG�=�%Q��y�v(�BQ�J$F8	�
���'���Ei�]1�L�1c�b�sΞ����:�����[n�v]kN�.H̉K�*����%��Uقd����9�M��ˆ�8o�����U��/��}eA��y+7�'퀟�E�J��;�Dn�Y�-ܬ�t��B�k&s�H��|��q��%չ��A���J=K��m���7X'X��f���k5����ϺGna���%��@a(S��K*�����
�׳�V^9�$�����x���W�$6�����܀���������NĂ�`�x*j��6��4FR�;:TV1� G{t'#	ˉ����U��H��2y(�砩����'>���ǭ�ַku�G�T2捽2D&-g����rO�\R>uf���VÓt$6b��2Օ"ɋ���\Cb�������o\6^(�CG���>ל��Gغ�uּH[Pt�����P����_5��I n>�琬⑀�4߹��J ����|ͤz��s��i5�d�NKt�*��� ��SҒUZ���=J�"���	�8�̈Ǯ�"�r������c�t�H�\̈I�ϟ@�s��3,V[ܻ��p�:��yd�����{��Ljw �咴}N"O��翉b��[R��pC�f^ӀI㍖9�)��h�S�Q!�V���^�Tϥh����>\$��v�e�W[�O��찎��7���.���-8����V��C��Y�6��)����@Ǽȅz\����J΍�&l��*xM_9��b}��D��{�P�dqӡ�vP���g�n/Ш����b^l(,\�\gNuٳ.Ez�����cf���iB��4*ϋ=�׆� ��5e�Tr�)%�,]~[������+6ʵd(� Z{��?jrTuܐ`��:g�@uDqD�8�š���&����Զ`lG�z>}��-:uD�M�-�n[�&�K�\
+GZ����ڟ��!��?T�I���e�K�.{��8�k��_��k�������G�/Jg!VML��F�&�5���t�)n,��&��9,���
v���)~�[���z�	�Cz�3r�+�_��l����K���1M��Qv�w^���rO"��Zp����f�Y�pB�^�^�M�<�2�	������� ���@�[�8��X7�l��ݬ��5�8H��U^H��	����Y�����~��$z�8�5r$���|�I(�8�k�N	�xSc��'Q���1�÷bk�⚤/[d^��ޣ��ڿ�Y2�j(� <.�e��2=&~؏���2AS��-�$���L+�z�N#��| �U�k2@�oe�"��P&�UL��"G�%�6N8�'gq���"�vK�g������"��A�U�H)!�S"�~�Q�fz)O�փ�uy����F=�.�i�v�c|�HԾC�Y��h�C�(�Ex��Ӈ�W�!HC����zjX	Lf���Օ'Ut��ߡ���Z��Ԣ��_Ds�o�LL�0^��b�!/����4��#*7�H�T"�\���t����=l��Ľ��O�!�Q�D�TYŪ˃�ȅn�"K��TSD�?Ҋ?����L��hD-���q�*{����:�?������x']�f@@ln�7�p�fI�R��sD;����W��ל������z�:p���`�KJ�zE�%Lyy�'�$�f��D�o<�v�
l���e	j��<�2�s.}x�����瀛]��a]��tg(���#y�%�L�$�5 7i/Q���G[��$�]e�-��nF��8W�"�g��4]�L)���J�*'e|ђx�gq�8W�t$��}���H�肈����'��%δL̳��\�bw�ﾯR%���Wyi�dl����̰6Z�Bq�>^�&��e��Cq>Bt6��,#�u'��<z��.!QGw�Ā�'�z���R��U=���`����,A�w�Z7tȎ 憟�D�V#?S�/�����:���R��g>���k�݄p�G�}��痏C���]���vә(����sz
��8�����mtf	QF1~Fs�<�>y�sg^�j
���u֛4��x�t���z�7n�J�"���iG��d���<�O^��uĐ�.m�~�z5(:Ɓ�Q��f�ß�\By'Ͳ� �P�QߴH��n���z��^<=��f�H�]�Sa7f�[�i9]"߂�^�<6�e��NϴUc)�l�v�F�"#������7�@�.G�����-O���Po�z�}#���^�l'������2���ٲd�!k�z����o�rs�y'Ⱦ�[���E��&[��D��W���}�HZ�=����U�����l֏o�)Ԓ3��9m��VQ�$�k��O�Z�sĕP���,&,"M&t�}�4 ���㟍��W.jNd*��W�������I}�M��HB���Ƀ��GA^*�|h��9w�0"(,k`�m�P)�Ź�"X\Y#��/e�+��8�����n䞦�l���GJ�/��� l�u .��B�k2���r6;��A�V+ZN�Kb��Z8%�$;��nE��_ɞס
9Bʆ	i1'��.䪂�09�LHlT��<-�)3�O� �3���z?K�J!P� .�**exd�[�ɗj�&6I��l��ψ��Am>��}��r┗9������8H�x|Sc�ϵ�m�d�!�F��I�0�}E��f#�����Z1_3jG�!�퉗��nl0��0߳2�F�J�
��C�	Q�@"�i�A�:�O��0^�W�iK5�4��^0R٦J��֎�����mج�r�BY���ڌ��w�>���$U��r0~�0�8{�d6�Yyj}g�����0��m}_�ʣ�d�����x}��y³��Fr=>q'n��o$�-ˉ���|4U��ɪ=^BZ������2�s��>X����c��~7�)N!�p&�J`���\�4��csG���-��4��2Fs�!j�^�O˟��px/�	��P/�mI����Iq�?]h<�b�����45E�d� � �c4�bΪ>P`�{�ˎ#�V��Y��;����e@�H�}O�z`����9��`Q騉�K���RF����
�}�|.d������eF�d����ʤ9dgC�D�i�ރFo����W�zL O`V��;SFM���a�.}� ����F��j��~�j{���
9�v�x��q�1R���/X����[��6f:ӥ�L��Sp���
�� ��1RVuQ'#|��9��
**�n�%0��E�B$���U(�"���C WMcʞeP_�Op{�|o��.�K��\�֛5Ҷ*�Fs_��[���Ŕ�ekn!'�xEx��[��lbh��m������ގNr��dp]�C����C�+��߸�bg_�W6�W��>�����^F�IU�A�(�=D�V�W�T�4�JI��K���X�5~f3ĭ��ׯ�"�隝TW�g������x>��נ�>O�'֥�aH��{��*E�	�#J_;����\,2y8�Z�������t�9c�e��F�o�T�P���c`�js��%���s���� R��+v}����$i�0�pxc�@�q���ND-�'ʜB�5�6�vpvjx)Bl]0Y����9�D���Ey;D�J�D7�!��}r2R����*��P4}J��Ӣ}�-���K����(2j5����]��ʽk��}y:m��*�䋾0X�L?��=˟p�n�T����Z��#֒C�q�g��"�|p��rko�|C,-@�\������~Ohr��v�S�]���@&�/�-]Ym�w)X�ض���qa��H"�f����b��:S��]���	�4��gJ�'����d�rl���~��9I~��7�;x?rX��~�fST>�N���ĩsC9���T���Û�3"�zl���c&2��>����{�k�6*���.�M�����ʾW#�d��!V�$o� �+�O�aJr'(h~/�����C�1#=��q�6�IR �[�>�)y� {L�~`��lQz�R1��yf���+��lӑ�l�ќ�f�O�v�KYv��" D��ፏ뷹г�!�;^=�3y�;xb|���^Np�r��:,zX��bh�ܺ��������[�d�z�b�m�m��/4�j��,���v�
�P��ʱR�_>0��8�^���ƵQ��F�:2�� �����)`�0R��C@��Jzi�N�^"�����ٛ�,�"��9�����}z�n�l/�2�����<��S}�ܽ��6���J����Dl_X��F�vF�r69+���)&����2�	�3����������C^+`�!�Zƀ����AB���I�h����'k�|Kej]�� /���E`)��貈�L�U��<'=�Hᗕ+��� �������ې`��^���)6>MAZ��M��On2�@G��İ Yk~5�����m6��d�}��*���*�zcv�5Ub*�vO�)�vwa?p<�=�+zt�M~n�\v���ʛ W��ۊ���� ���I�d�5�-����zHAB���) ����%�hP)���9�:Jae[R �}X��W���3��(�r������#m���hXH��;�.�s��6U�n!Wþ��Xw}U�z#S��.o4�3�yie>��!�$��E��C�]���E�h�#�Q ��ۧ�wє�"�:�
G [�'}'MH3� 0T�7%�(�&:��uWOj
�z] Q����7ی��.N������$����1�3}�g�r�VP�i�:�(ث-aI��d���ɧ��x�ۄ��J/X��u���N���iU����k�~��	��%XU0qxk�G����t�KM�-�d���|�F�L��F��C������B��s61ۻ��0sq*"r!L/�sP@A�q-�k�ɚ�y��'��P��֬s��']��m�#�,�8T�g��=����ֻ�Z�*��Mz�]ܥ�eê�< �����r# _2<^��N{����boN��b�6"iY��sO;��(�K�09�"�b��L���P̠��3hģ.!8�=<��5W5+���A�@�i%���r[����S��" k&��:��R�/^9�Q�6��w��w�:j���`]�S�ن����.�.�gpp��6ѥ*�Y6�#�p�t�-$�w�Ȇ Eˍu.9�����!��Ǖ�p�#5�Bm^�6��Q�\���k���O�
T��칛%J�	Xrc�쯓�瞮����T�n��L�`�f;O��('e��A�jKG�M>��N���ؤ����:8��T]�IQ�[����݈>;^�Q_�6#����#i;���\�(�
`���?+UV'�-4��e˖8�K78�S�M{j8�8x����*f�
��U5�P��[h�h7��z�����U��J~̅�P3��
��͝%A�Bd� *��=�{4�G5�~s�5����i���g���v�a���ǖ��q�Cc^
�T���7)kl=ͤ�%ڳi�Jh�uU��$�� ���w�`�.g���E���tc-$��������f\�]���s�HA�}M3Z�:�.�:��ZԌ��=�Ը��fh�&��o���פ{�)b��8G^^�b�����[�#h[?�]ò�7i���kZ���e�0[$BY�]�"X�ot^��Q��/hcs�aR{�������Wl��g]:��pkX'�nkA��r0�+���:A�8H�Nnv�P�n��-�[m��f��^w?]8f��=0[�;��|���0���8��r��0���x�)�m�J?.dJ9J%�[�y�(�5���,US��mo��?w�_%�����y2{H�%���Q�%��+����46%�	Z�^l��[Xo�UMȲ���S��c��y���y�EAY`P
���چ�3H6��xs�Y�|�a~�"D���(���f��]˧}0 ����w��gG�Z�e�F��/R�S=�\�W,�s��/[�UU��,�o�ƅ��蒣��48 ަ%T�$�}�@v�-;ia�e@��K׈�=שB���������Jۍ��U� s��'H����da��VI��iS����<H���b��r�+D�,����ꪈ�(��]׏Dy���ӌ}f�?�t���]���_�˰�u�(J�,�	�Y^/ԯ���G��%�QsoU�#u?b���@�1.K���D�3�!��=[Stt�����`�O(y��%Ey\|lj8�f�\��Ae�T��&��0tIM�;(��]�T4�$��̤����o��(�2E1#�1��ĵ�k�-ҽ�Q�3[:�*�fbl��nNb����/X��l���$��P�W��S��-�Gg"�	�}��!?���ި���f�ٜ�g�U���}�Lq��部���{߾�df~�_�v�JKז����Q/����8�R�HRj	 AQ2 0E�x��LDU�N��I�넓��I�V� c�r��dp?��!����Wu����p\��{E!E���ec�áȰ���h(fw7 ��j��m��Z���p�А�p�hR/Jd���y&<�j��<♧9�r1as�Z�$7P�������?�mP�5�z�/m[`I�ɝ"M���v	Cz3#u���'�2~N�HɎpֻ������4���3����Q�6�1�h�nP�m�
vX��T���_�1��S�ǲ�}D����1'�iuT���>{G���6��M�`�?\Yo������&��Y�4��K�t
!:q�<�T�٘K�g	���"�GH�N�C7Rs]hr˾m|�+I�@�/�����Һ��Ar���cS+�}��(pP*TJ�R]Ͳ����jH^xS(ʱ냸�� �JʇT��pYF�:ڱ�3��5��.�id/��9��w�a�hn��<rC�i}d�Kű-n����	cjYac\ý�����a�jo����F�K)s�oLq�ǣMl����N	�;�9!��/6���"��b�a�.o�[�J�$��1�':��H�
¨���SUJ/o��㱀�Y}��ˮ�Fb�)�4Ο�6�=�A]��[������\߮';Y�ѥ���8D��S?t�'�ӗ���B^B���8G����j�>og�_������U�'���t���\��0���:�V��TJ3�����҇�E�C���&H745^��H�G������V@H�6����5$^v&UXh��/Ao�T�ǒ�L����My9�	/���"�bvoMރ@`�	_f,g,�uq�O0~cj�\��Ѡl,8�U��{=Io��cd���q>_b�,��c裴���H`+I��b��Nۡ�!pʻ��D����g�ܣM�pQx,��,e秵��q k��duͼXl�{H�^�;�VucǶ(
�nJ��R���`�S�"���YPu'�MTkXoT����˩S��m��(��Fu���o�_=|��@�'�nD����-��-�%��F����>�-ٻ���5yO�iS�����W� �]d�j ���}=T�
D9i2�=�"bPs;����_z/��֞��@3��`B{��)M�\C���U��b}�zݹ��F�vаWa����oMT���_ۣ���n��F>�}��?�)�x ��W��'��Ȃ�t�2���c`�_���(:G����#kIa��OJ��ض�l ���\L����fSX%�s�e�����5������aI����S��fT(���
wX�8G�,�σ,��pT��7���JR���鱑^�&Az�9�w��^�W�c$���.�=ɀ�:T櫿�+�`_�(��X�/�(����� ��Uxֽ��C<�o�d��,���r�����H5�:a��C�����O���W��[�mH�U�c.���s�p�
c��]��!��W�}r&�:9��	��c�8�i(p^I�[�m��y��ڔcb����70tfR�1;�Bϫ��?	z�K���A����H��v�[��`t��ߝ�;����V�ӄ��dE��Y��C���ZMv|ֱ�3��d/��z��r�V������DWz�V��*xN�F2"�SiuV<0���.3�)�8�
%|i��pg�#�����	�",C7�GX�v�(�͂����y����Χ����]���Y/$+Q�s+�%�{�