��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�#&��#�<�����;镬���IӒ��wf�����`��ONl�C��>�u�0�w�S.Th�dMy�|�����i?���$��	n#��͈���jUl�f�4�lR�x��6r��X��SH��l�Md��v��L�����<e�"��!��%�b��~L���djȻ;S�w�b7��B,���F�(P��ٻ����G��{�S�}�9b>�%6�?�r��9�8p�o �e��u�Cvʘm§�&_Gq���\�y�b����A
�ǌ�G�Mٰ���H�s^'��m۹������Mf퇇��L}ƙ�7)MZ��|n��I�5�3�k\�($�rhSת�Z<Ey��g���={
�<Άv�m�Q~���ӕY^�j�9x�)�MA���@tj�q�$t8,3��R�v�Ƒ�>�h��0���R@N_Abu����|�/׻�Dwwɬ�>���A�0�cHF9փ���.�i�;��;5�<_�D��ɓV3�|k�6B���+�㬄�Fу�������T�*R"54>%wߋC>6C���X�,��d���}���V`�j�S/Mz'���@�^�^���"WTC�ch�!�Y�q�ޝy��� �J���V7���e��T�TE�T�>|�el�-�����J�qMp<f�slo�N?��μ ��s}nh�AB��C"k�7*�}ݏh����?��N�d�2��j@�LaI���p�c�8ΐ�~�q�I����̍3L���G�2�� g&\��+�!Kq������ɩY�,�@��`�s�S)7RR\���p@X}9�HD�'[R�#�&

<P1\���`Ŷ�F6?,F�Uԛ������.{���P��h|�%����C�:�.�+�Z@���Ą������a�l�`jf��F�-X�{3�]^GK��Nf I�I���j�G��Tl�c��z ������)Ҝr��ߜ�9踸]��v=�����H>Z���!:�&���@1`�h�m�a�����*t$�oz�����v��p{+�4����o�w�y��ǽH+�أ�h���7v˥���i�^(l$��<�����*�����@,1G�*��\q���vEĤ�Uk�j�ݺ:�gSh�t���
�O��k`�^D�B>�cv�#���6�
�4[�kUt&���RHv27g%� �&�1$-�3m�҉�Ƹ+�ޠ���·Fѓ��[��+ӎ^�YO�&����hó���I��(=����K!�]w��ُfr٠�)�9^&yggLc��-+� t��T�Q6�o�3E i·q��
S�ќ �l�ͳ���������)��w9	a1�S&}�n��IE#��ƕ��uV�yJ�Qه�UM�Ny�p�W�W�n9� �)����WΡn�s��6���wpw�$a�#�7 Q�v��_���&��ʨ&?��|��Y��?s��x�-�K1 2#�B�j��ڴ�vF%~�Va1a�^M���4�ոs�O�J�����-�oq��@����[L�^"�S�F�7,��Adfd�Es�J�����C3::%�RgOb�y�Kऔ���+�ERs�s���@N�!W2n���0l�gxf�����\3^%�yj(e�me��yc�ť~��J��8���/zՂ�������(�:�*����
�mL�pC���,��������J\���aZV�^�d����v(��=�<�o��gY�-FtO���Ĉ� ��4t�zi�zI
"�o��␓��.ޮ	9֤�BM�v�Jc!��I�-e�g��*˜i㸭O�oss��17r(PBLJ%������|-ޢJ�*���r4v噱�d��G|��_5�D�TB�-0�+!���f�yGP/J���R1�b������6w ��z���g�W!���N�J1�Q�ܓc�� �S/�m��')4-�T���sy}��8� �L�v�2��v�/�W���W���Q�g�7�A�XX�[��' F�� e�)�$'U�q���=�f��-ȅ�S��t�K;KB��n*��I��S8fr0[��V���A%���n�!�pgΡq��f��~\	���9���G�PS��J�Ȁ��;5Ө4 ��w�e��w��&4-L�l�ԓx:��4���F�d=f}R�*��2Ɏ���g��[xF���i��U|B���M�Tmj�1�<Ϝ��jAY�ѽų�r��l��?NM�?�o.9�,y��8mj� � �A͠<d�$ؐ�u)��Dp�J@3��zj�ի&�{N��o�R��'��IZ1O]���� �#,&�� ���{Q�F .ۆ�
B3�2�C��{p�N�Ϥ��K�����!�Y�5�����lv�Z�����	iJ�]Gnc�*�;����'��m<o�l��8�n�ʯ��m`O@�a�����h%ٱ�tH�9�bX�����ɚ�v��;W�L�ouԝ�j��$�Z��,.�0��\��V�C,���KR�*A��#<�>����Ӽ�C�i/m�Щq�������Ǵe�@����t��]{fAB�Ё����;}2�ô�&U�j����~�$n>�<�L�T(�D�d���޷q޹pb�B����c��V>5�M���^�	$aM��d��4YΌe�FSͲ���ʄ�p�^�r{�P%磁��T\2`pI�����k`��L�X5'� �5���p*.-o��!��0���bӽ�]�_$�ωE�D�j�[���7�!���7�voЈ/0l�w�F;��!g❅Hst0\|Ӧm�Wɍ�~��.�p��n�_MW� � ^����J�	��]K���2>]T���Ӄ%�j@:�+�����ڑ>�W6�(��-����0�z���i#Ϥ�p�"T��g�'���YCy���)A��}�����z��)K�y������xiD�
\S�|w>D�xZ��UDG��L-|����% ����5I��Q�H�B�!`�ˑq��OY#.񭿨%�3�'��K�JU�	�B�����t�ىk�5}�RG�
"�)�B31H���_q�~�s���\|,B��,�5����zڮ�ih��%�����{��9쬇�>�9�atd�ϩ
�?�ij�Ÿ��~L��)��+$��p+E}s�FY9�^ݫ�i.MB}=��_�ր��7�ߌE'rd{Q�����eO�$�W�0���Y�E>V@�N���.���I:'^��O��e���Q6D��=��ň��n��n7yM��a��9�����26��5*�L*���QU�ʗx�=� �1�Z]��"_5�#_�VK�Ha�rY�q'���(�f�݉񜄍<�?�F lۨ���y���m�:)�o�	 ZD����9QR�W��5Y��{��-��K���:������;,7|��'G�u��T�6	��v�����H��o�-�2�{Z �(�E ���HӺ��m��5D��S��/��j����>����?��bV�5�_����	�TŤ���4����q��c��SG\s����L���-��;Uz�}�}r%
j8TL�;�St˵�)���"H��Yx���c�4]��x��od����
i\��C�i��qk'��Y܋�f}Q���y}�55#,�~��~�K�;����Wqjɋ��*7�[�����Ř=�f��
�|Ӎ�/Ю�%g���Iŧ}^k��Ol��t��4T���sYu��*{=M`����HDGl���c����$@ b��ao:31ݏ�e��CT��:ɷF�`����fW����g��@���$�`��tB�����8B���K~ѮX��M�y[#��ࣔ�)0Y0�]���F�ֆ$��E���+YU��% ��Xx�R����r�	��2'3Yp&��8�6n�?S��$�=2NP�����G �y��k�nX�����mYRNW뉑����?��ٺGw�lȋֹW/�_��@��9U����;�`�"T�9//)��#�F�����w8�dmI�(���D�ռ�Q�~-DLQ��j��������H�ƍ�\������y��]i_�--���p��9�!8Hh(̄s-׹�ml~-߻��$?~mQ�Y.ki��~&;Y��Bc���L�i&z�I���!]��^�/�*P>���h<e�"P��0���n�'R�%���_X�4_�X�t��xg�2�-�>��;�I�E�S�e���v��`�q���4���zjeK)���̌��WB���r�_�V,xGEv�7y�i�����Y��-��8�,�u��kS�ƨ`�`[1��ìg�s�m�GOxzr��4e�@���N�~�(�O�S��v�E�(.˚��wn䋈K�#�S�j# ������T#~��Bƴ��:!z��
�G^���Z�Դ��q� q�bjʋ1+T')����X1'���%L3z�YF�VLA���@BR��v�v���p��zH�R��=�^8����1ZD�1�&�95^A8�Y�(傪A=�*��1e��͋u����iGQP�]���eaU�Z����tCz� ���+�;Gr��U��]��h��0��s9��jW���IT�����o� �$}�OX�d��?�W�[QppL��<ER�l��V�}�WÑ�����;f��CB}Ji��x�춝-�n�ީ;��4��� -�BF&�V�6Z�@��av�����	z�c9�ޛ������4�!q�,�r��'HIE������XD�ob�fb�S��r�����U���J%�~>�KT+�kl�A�y�7*?.u�Ң��uu`���:���t:ǔ�,A�+���`�>W���4-J�e�(Y���
�LbRk��T'?H��qF�.�3���7�G/t��:u�%Z�L�+�+B9���W$����u�c�������W�$�x��m��]qQ�M���VfK�y�2����cȥ_��8���,/��A�������[
A��I�5�ó�����[��q@#���`\�D���|��T��x`��Ml�)�Z,�����e)��Xͳ\�Wa���ewk	�� �s�N�
#���+��,�h�Sh\��W�/=�?��Q���NaSQqU��h�K]j�ed��~��������8���ȹ39^�vj@�x #'W+�-��fe�fb�i+�����6l�ƄX�E��`c^1J����K�╏?NS�m�~��`��S�W�q�89߈��"�q���=�EF�m��Pf�=�D���"�*�i_���J�!�g��W�,U�;��o����%�NM��������z�ڃ˚��9jT�{�P��*���㞓�<PQXx�2IIÈ��������g>���������a���:�!�E	_5O@i�� �Ԫ4S�T*�;8�\���!�o�UW���m�{p���h��(��U�ph����ၫ�'<�jra���i�{�:����G�J�L�C�.�0��p��VQ�gec��7�����L�X	%��^6��������U����r�*���cZ��#���X��T��=B��l�+��q�"�>A�5�����F]d�)����3_|UQh�VZxk����\�Rx�;TL�*?�q�mnQ�(���y_��|�c����T�)���)�x���.O��_�9@��- �H)�3Ce����9�-��BPT���L�Nr�)��$�Q����Nז�O�Y���'�o�>,c憼�3����h���^{�Eq���V+P����$~j""�3�8#��_D�Zͤ��t×�V�np��t�3~;�3�w<Y�]Ts{�����\��
s �mfn�<�3��|=⛼u{��4�a3��OR?�-�A��z��E�#;mA�Zc���`W�I:���������PE�fW�%�h:�:�*-8������]p���[qg&E�����۰����(E�i�<�JM�V�$^)a�%���`�Ety�(ከ�n���q*[n�y�,�/?�P�����H1��Х����i�U�nY��i��"l@���]�w�z�	����6��5�NTD����V�dqۄ��x��878AU44/qF|:U)�2����;b�"���0f�#�Ɩ�'�Ci���K�H��4J<R�M�6�q�(CN,Y�#��.Gv���wHi��I��d�L�f-N��T�c�A\L�%�9����$=�ʹ�j�w;�^8�x�k3h��I���Y��������;Y/���R��$�»3]k�۱��-����O���=�j���sd-Y2�T��NV����mB�d�v�:�����K9�H`J�En4�i]��..�r��h��������5�ޕ38 ��a���B��oB�.��>b��>BkCZ�W%!�FI��t=p��mM5G��j����\�4wU�)oJ&؝�r�����D6�� K/{�D�x��e����B���|��3;c�w�H;˹Z7^�����O񄭏�SL}r�$@�Z��	�&�S��D ̱�c�"����	�X�8:4��.F���dqO?�u�R`H /��B�̌_	42)%0!��A��K�)����PJ�L���Ƞ��7���� ��)��)Qe�O �HC�+�԰��5��b��@
22v����V��p�#�^u�!'�$���_7��dE�i�3�oϜLQJXH��&���6�c��Rٜc*���,n?v@�{a�,���bo+�6n \��!�\ɘ����i$��u���y�j��9ntu�0��dg�o��:���؃�e[Iq0A���.Ŭd,���l2>��g!�c�c8{���wevy�D�����*�_u����r3���5�����H[����z�i��QO,�7���Q�>+��9
�c������Ӽs� ;���%��������y�X�����xF�y�i6M`�ʴ����v�O��뤝����2 .���+��H$�s2�3�k��5��Jd��VʁqY�� X}�̈́#���|z+?5���X�B�1�G�%⻧�%
����w��������ѧ_���tc"eF�b h�� J���<��Uu�h�4����=w�)���{��3�x}X6�G���t�E���%�C�(��J�\���(6�F��B��s��;6"8M<�q�Lv��Q��C�[j���wͳ��5��� $��ז(9S����nR��c��tY���l�s4mg�7S��rWѕwO��`������X��k��ƻl��!�G�X��u�ʧ�B}7�+����Mz��'w�dd�2�@�/�w�1X����������i�C?>"���U;Y�'���SR���y�Ƃ�>I��W
�r
�(v㔅���<�鿋:rD���Q�)3Ǽ�Hw�\`�W�$����E��H�T����M�6�N1�n`�������P2-n6R5�:s�5�vz'�RUV	��yWx���$��|�t�k�ny���Y�u�?.dZ�P�EI�m.���H��t�Z�MR^�. ���Q����]��Wj�?}i��@�Y75U����gދ&��&�;��Y�)���E�X2�(�NJ�į1G��}�����k�	��Pt�������l��[�ȃ%��d�����E���"���5���,���Z�n�BM�a��N�����NMUv���R�n���"���e�[����-7Hp�K���Nkh�����!'�Ӑ���A�����t/D7�U_��rD&���D@����P8�oç�x�=�%�582nۂa�D�Y-�-���qh���ņ<�rK0+�p@� �* ?]���� %������b����E��{8��ڡ���#(xJ�ą�=���"�R�}�Q�����c�Pv>-S-\\��_w�*N_*>������$tz���H�=C�,>�S����79��:$�\1��Ұ��5�@�X|��e�O�P�h�#�K����������۩����n�r��=�ג(P�}��T���j�������k�zPQ�&�>J����Y�@A�۹��Ԋ�c[j~l�؍�1�wPQ���h)�$��Q�XT�#�ޅ�����D;�7��y9���qy��(&,B�Z�e���$�v�W���EX�w>��0���(S�N�����a���Nv�M�L
���g84>�(kOKA�?�p�ƈҎ8����{�8�.h����zeY����'��B.S�s�Ҽ�7U'/S	4|H
��Z\v��d>fw����'��3�@��f����t�ݳ�8k&x39�b4R����~n���=�|XU[o��
�{6�?(e��dS��3�rc�A�:(��#DGP��pYnwR`T�(݀gD�'� 擽�3�����G*���u�f6���d�/��Z�T��OEW�Ti�8��0�csS`�9'���X4�U`�o�$��l�f����:R�/�R_Fch戃B�0?/��iJ�qƪ����X 5$�Ef�� �{�@G��r!��6�k�� /�յ�-��cg���d���.ĄF�����-�
ȣ��.4Y8C�9������9+�����$4���Ӌ�Ga��X��X�ݝ\�v-13�������Ͻv�
t��{��o=��V�\�a8�+��n�e}��s�m��.�"��Mk���ҕ<�_Xz�� >~�C�AhB���-�I���D'7��k�U������Akr�
� �H����}�?��I�Z�����ݿM-o��g�9(�u_X��:��1�z2S�O"P1�p4O\�(�ʿ�j(t�rw��0.VF��S�6ƅ�wܓV�٩�5�,��x��y�����`~o�drr�Og���zN���{f]Qd�G�2^'�+stЀ	̏�!I��IK��:}��Mِ�L,/Y�R�*��x,��N�u��l�����֩"� �@���l�������,��l$%���Vo����6��Ov��&�`�+�߶��1��%]�Η�U���wQ���T
�Cy	��~Xa���ǋ*��:��*�JȘ��(��� Ӝ&C��O1�� t
����̎�-�c]G�r���r	�QŻ�ӡ�+�!bw�q�A0��EP��"��)����@eɎ�y���U��gx����`BM�����9F��W��e>\��1����i���!gv$FZeZWT��f�8�o��X�n��;��֨?��G�L7��hoD���<'�^� H�kC��v��/�[<x����������)���Ƕ�bs�*����xv4���}��k%X	����s4Y�҉�a;"�9>��o��F�����F��di��:��a�P��b9��8O��e�2�W��l�Ĵ���T"�c�t�s%&�_)��T�P�<(���~��g=4G8���� t%�Ï�3��f/{x��h*h�A��;w���t�O��%6'��%��x�j��f{�����`���p��?rFd��k���Ԥ.а��!�66� G�� ra[�zLJ�fI������������P$r	���R��j�z.�a}��_��  �j
������Kϴ��ŝdE���@lķP�*�|��>VH^��m��c6;��m؊W�)��'�Ym6�D�&'L�h�LR�3�J�ծ*��pɔ>��5ii3Ro_W���{yY�]���X��J	����t�o�Lj���a�p��%1��l������K�{Ȫ��p�Ә����P"ͶK�y	J��_�%X�pT?Mh#�{Ap��r�[)���
��j󖜯��_4���D�R��_m<	�ĞcJ@���P��/:��Q��ܿ�����wF%;0�&}is+O��;�OR�NE+�&�ߏ�
�^t"����DtP���q����i~�Mw�a8�^q�m,m	pӥ�<�%��-���=�e���*k���'>�T)���W0P�q�t� �[Z���HJ0����ɒMc��Q/"(�J�6�l�b6��1Y_�	�P���i�,�M9�J�ꭶ���U�����>�9j�J��ǋ�B �N�=@KW�E֯�v�@���0�	T#3 HX.4�q=�@B����Jf؎�ֶ�O���xw�CH��٫
bx�܊��N�Nc"���҂��a@O|�x%o��<�5��3�߬~&ล·�AQ媸A��dF��XC��B�IhY?��U��e[vS1���hI��֌�{�r.���wd��Ƅ~�H������;M��wO�K��e�a�Ѯ��dV�ȴS I,�D��Cç� 俑#��>qN: c��_�2� ���̣9�����T9��l����U�s�`���67e:3����֫���{�Q��-D�����7��TT�.3W'Q��'G��D�t����G�1��Ҷ�R�0�s�dW8���+��h��7�s���NI�hP�Y/�>�\xa���N6~��J2�u���p�f}�yfWou/]]��[�"1k���#VO谸�'ùA�(J��_�;�����x�/�]ǽk�%PsRכ������Z�~��:��v��t	䣪
a�u���o���"jByEItϿ".[p��d3A�^�$)�
��=�`�#�u-�� W�љ]y����f�����E4�9�v� ��914���)w�g�m�u�,۴$0��翓�`���l;P�'4����&@H����!�I-��#���C�U*�?z�ą(�W&�ԳP�*���u%���iR-�o�a*�Hť�f9�(J���BßM0qhA���as���=�2m�.�@Q
!G���V'�Ǔ�	ͦ� ���"�'[��d�i-:�^o~p��V��c��P��%Rj$'��P_M�v\y��gT�t���c���O_H{�:�NQ|�Rw�
�_uQ���H�&tb]�fKv�9��a���������X���G<\ErUv�/�C��V+`���y�@˾����nV(9FR��.c���#C_���Xg��l�Jz�Y�1L�y�Q�&�}��΢>�-���[���?iF�k��y@��qT�M��F��  �C]p�d���-Ηz�r}�M��X�=D�_�����"F&�Kق�ו���i�ekL2�ɹ������U1uS�F\�8r`@�{gO=ߵ�z������������+ �*ni�����.�\�
���5�)���f�֒w�r7���-RK�����?w��
4_��< *��v�-�>��l9/���d\a;@�b��7�~�n[��Ͳj�2�?���q˺ޑC���9���I������&��F���[ڌ]A�4�*�SU�	��y��1'�.A��W\s�wΙ2�E��+G�Kױ?V�Ƚ{%<�*y�u��yM}W�>x�H�u�_�#���i-�LD>~V
G��&��B�u��j�3��������L	G;�(��*��z:?΅�@Iz��nAդ�"'o���t��� {��6#6Xr_n4z	��D��И���`���~�V쵕�Q_�^Ӊ�ב�wZ��Y��bV)���{��r��_��f�s/�3��7���ZT{���ms�nm�� �D��+-
�������\I�H5|�K-��Z4&y⏊0h�}r��,����}��+����^�m��>&O��Z�O��!=*c��&�t	�A��P�>�B=방6�x�s��S��p�����J=��Y�Y"��M���W�H:�S��v{%`I���Q�-������J!~-.?�`��c�"�Y)� ��I��E��4<�0���l%vGл�s���#��OB%�N���;����tQq�-��u8I�������������I�ۢm��/E�|�&�Bߜ�&���2�x=�S�yL �1s�v�-�JF<��g]�݈'M��7�Q_3�8��iUVB�w��_�I��L���CW�!�/���R�s�l)0O�s`�&��-�*��d�B��S������M5fA��n�4�P���nF��(�?�.?�0I�	��L~M���v� yꦲ6���6����|SE:B�}]���㞑c�:om4�N�*�{`�dm�؝�G+�����ɚgP[È�L�fr	1wS���l�L@�7x���q��<�q��U�4)�w	%�s�=�Mm�&*7�}`[OTc�@U��3��*��/�T��
<mP�N`?���'��^�Q�Z���H��"����c/s~g���90���4#2�O_�l�/2S���?��V汫[V�\�;mt:#̇���-�$%�bˣ:0���`96o��5�����ߣ�)9C<N�1#5���'ϥ�^�
7���W�ȵ=�e1�Kil��%��1��1�"�9q��45��w���H!*R���pop�cT?���H�������H���[��h5��b2�/�����X���ct�9Of?A�Q3q�
B�A��ٛT��y��Y�1rl������m�_�6��0I�������~���-�M����;d�I�ݸ�����7�̸� ,���'P8��t[��~�˲-����>��!!�c���`���,�\��K�br�X�tH�D���tή���'��y�#���q|�NV��G���d�b`T�~�}H��F � �1�^/;앤�B��ؓ���j6QH��/R��fV�� KA%�U&6�s����j(,�Įh��u!�6Fk#�ٸc,�
O�B�ȫ��2EbXRd��4J0V}�ږ\�gOw|����TG��r��<�]t훃��Z/��KE�8Oн'��؞����H�q�}�.	l��P3-,�S/6}VY%P��WHX��!-��y���� �-� �������N�Dp�X�A��z��i]����פ�ar�UlϮ���vE�B��S���DvRCK��h^�d#f��'��|�L�C�j���Qě���'����8 ƞԙP��Diİ��R�c�i&�`�
�c��&�����p1��r���3���S������@�z���W���E�ƞ�Z��� ~��f���RȰ��KJh���kU"�Q��N�Ʉ��7.{ID����b��ުt���	���ȵٷ4�aT��z�&��GL�&��Gӵ �R�'�|�ڻ� ��$!�'�oI>K��+[���G��5��oX�/�hC�� Zǆ)�1#�J���\]Z�]�s׽sg_\��A�U��8&f�2d��-K���@�EjAa��F}��&\��u��.���	q��q��[�h��ZDAL�2P~�d��7SH��o�F܉6���CK�D���\��̉�Kr��]�N�D���啼���Um[ ��՛h��z��U�f�$��a��Ȥh���~��e�:3�z�;�>�hl����t2�>Y��ܶ��y'J�<傓��ϲ#�iF�y��L��
�����5l�{\kO8Yb`�H����FR�)o��A>%S�l-W�l�.U�9#Ζ�.��s_ p2@���9���>&bN�|�P�������ִ/��C�[�!?D��/x<�{0�\&Ⱦ�?A
��0le��j!��Ǭ��_���ŧFy�e)K�QThE)���������	��Uu�G��=D׃&�Sc���su�3>�������qi6/Ms��T�p�&���g��y,���� �CW��3af��?�����Ij��fU��@%��J)"�#�d �ҙ��AS&40�Cp%0�K�da基��|�i@8��v�O�fз	�w/�
�?���g<�Q,��,i�Z�����!��܁a�� ��,s����/�U�LR�����r��G���[ߜ��@�2�n<$M�;&WQ:�����Od"�K���&���.����������:̪{N�}L��#� ����y�-�$��_�.��MRQ�t�*]cM�ݝ��5ǧ���Z�ů��rd�֊d/Cބ�v�o�hVX�A+����7l�L׀f%м��ASp��?������Ҽ��1���� l-�f3�{��L�<�6]�#�b�l���#@F�4r�W%M_����'�]��D�f�46\����K�Sb�7@�H��H�˂�L:�@�t���7���s�"�#Y�Q�yL�gul�4�惞��pU��i" ����{9����籖��q"�����1�gN��&��y�[��j�ʷ�DHKV|x�B������Ro5s���&a\�nI8� ����5"���iIw�FS���������p�}��b����=��;���2��<Ճ�FH���!�]�>�nWel��@m꿥*kb.,p:v>EDY�6�g՚�~6��E���K{S^��:��"��q�|�"��Ш�hӚ���T]��$���`���J
o�%?<��+a6'q�(��D@U� �f�'%Yl���y���@̋�e'�.@_�d9����S��.�3�^_�<=V�J�ͬ��:��'�b����~���-�V����9>J~)�;��{��B؂��,pa_ߚ�`@jW.ϸ��u^n���e���$Ӭ�����bSB��ϛ).[\r.����jpF|
�ŬK��N&@�(���8����>���[�!X|����~�|�㖧��bK���ވ�v�خ�Ѿ��Ðd����}F�m���#�aMnX��]c��y���G�"�0��¦��@4&OGO��;4a��b�~�ks�MV����a;���o�F&Z6;�3<���LB�uYe�Bc�Le��)�لuE��k%�R�U��5��ds��_�X�d���o�3t�	k��������L���bٰ\
5����d�kݺ9����X�e�͉ ��yݚ��uW������i}m��?���;KQAcz֘���� ��v�%�#\���}��˶ϓ|?%ϳD�.F_�aoI1�uf�
���Ӭ�־�n y���|ZA�B�͙�:�j����yD��F;1�