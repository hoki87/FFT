��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ���������./���+��`�OR�/��c���D~��I�M�,[U�yWw'��R/��ԏ���nˊ�ڣ��P6BS��	�=P��Qae���-����;iY��ϱa��v�)�����
T��)�+Ƽ.�M�P)��By�q�x��H��ϴV�8^ʱ5���D��[M�;��el���4d�{���5=/�+��=���M���U�@wHϔ�Q8�(B� �'ڬ�AHNu2X�(x��}T��K�{�`^i��?��f�z1R�tx	�}����r��#�}t%����a�Hq����X����&ZC�Z�C��	������(Q�7px���4Mg`�e�bN�u8G��� ��z��bn2��ȶ��H'�3�ªbp�"e}X%�E�G�X�V'��MiDc����z��I���c�C4�N����A�d6$��Ӏ���!�� �Ø��\���`�H,I�!���v��$�ӿg/�@$�z�
6��r�������&a疵Wj%a����א�t]��W�+���n���\�6�Dh�O�oJ�-��c��ҴI�k��X�;C�XQU-��Ǧ��z�Y��LS-y��*�]� �>�HAk�^=�Z"g�."�
�A�8����a�9�^}�`+}��NkRj�n�&yF^���'��X� �(9�``�@ω�`d���/�����4a֩$�gz�������o)Lk6�s9b�7����n:���{+[iQ�aB8vd��!i�Q������w^�٫�Gev_�N\Wl����zO+=��=aH�{�����[2.D���$�`2T2ACJ85�yҚ�p4���T�&誀ܚ���3�p��&ѭ��%��U�j���I���2=+K8��Gw�WT�y��p��`"}e�}��y�툂��d��yp�c
l]A��~"dҦgm?�f�y΍��B��Z�8�s�?�:%e��5����x�<�\�M��6;��v�����M�f&w������9UVB	�r��j�움��㠪��7g���Ӷ)��c��,R -�m;���h�fQM���јVYM){�J)�$$:%� @�
��f���j��� :b�]��9N��K�aI�k�?@[�� ^MV��T�Εy���PVt�T11�@�H;�҉P���2��;g厷�����o�|͚g՛��L+��~��{֠f���D�T�q0P"L���i=�{)rj@�{�k���~�GV)�9޶T6����}�_�W��(B�)��´�]C:�v�T�C��ڛ����&#���Vz߼�Bc��Ȝ�K�g�R�8�h�a192����#g��������+
ѐ*�a�S�î�!%�{�2z��|!��̕X�'�ne����� �{��u�|��&6�g��-`�fZ95uz���LG�mszHL�<��"Fl`(���O�r1��G�{�A�Qc�)P\Ex�����b:�vqx�B�f�Z!�����l���w߅5t�ΕS)���єQ�k���C�g�"\�����BW4vS*��3�	��Sc�F���K��u3	�]���g��#"��7W����s�b�1m�����2�����J�pS� ������r!�ūǺ�y��>�$���۹�R�7�O�`�nz�I��1����BHw���"��ĝy�i<w��"���ۢ{��/3;U.���u�ܣ���:D�-���a�c.��J��P��t���8Y9�Fs������7��w�JA�p-�K����S����3��\��VE�(^+���t�Ib��G���0l�'������>Yo�G��f�!+�[�h�H4���`�Q�Q_�Ƌi0��K���#����n��% SW]��b$���`��I?���������+��蹲
@_H|L>��mx���*��<��ᱟ�^N��x�������*`��+��~X8a������%��I#�sѦ��| �f���!��)�=M~�p���_-�F�1]*w���*����i�����Mo�������^�f��(u����8oya�,J��:�t���xZ�HO���˛Ԇ�ـIӪJ���Vy0��^PծX0%��p�!B-�9�Qp&,=L�q ��n��!��� 9���q
��PްG�I31�5�uwRt'�'PTs�լ����
�0�W#lQ�[ϧ}����WY��=�7�ս9��H7wA�uu�}G��c;�8�g�����v���CV��#k�#ͫv
�0���<�ӱ-x[�{�{��?sA'x�y3�h����#��T���C�5-�c!7K$$�*��.���l�jH��:�!�J'�>��徑o	��N��$�r"��`�d����� M=���Λ"jD^9���
��&%�x�u>HF���Cjk���G��^��t�=-� X����FJ�TW:yg�W��!��_u�IT��|��.Ҕuv�>S�9�O�
+��A�x��QZڹ�R@<w����u,h�z����޽G�/��'.Y���8o�;��~v�sN8�I��a(��-A��i����n��^j-fN�c�S��w&�X�۠*�r{{����t@�"��zΏ'��ϿI胂����Ae^����z�wFJ�����J;�6�+5�6�T�&�/N9��ז�:��Ѵ~�K>=8����O_����X O��-Cg�c�OY��"*���y���Y�ξ4�9E�(Φ}ȴ�7�ƴw}��j\DW[�m�E��e��䍚&��K��[����B>%S>1��J�has�׍iDoX�5lq�s���(�|�7EK# )�I^�D*^���������҃���%���ch-ж�qO���Ć���;[�'	j��J-�/��y����um���I#��T���=�� *�v3=���u��_+ߴϬT&l�`�vCw G
�m.0��� )d]�QY��)�q_D�5��xe;XĜ��'��<��B�h.��p�e�����{�����U�5����l���Sr�S�WR�A����o%��Ն�Q��׈��%��ZV<b֞@�#~����F�-;n�Sўt2��K���η=�W�t���]ʥ��t��d�ĘٛL]N����S��d���D��~�k�N؅#���y";�2l��5����r-�?^dY����f�Y��I��>^��^ubٛ ��VbHTb�ֳ��`���|R݉�2p�Mt�D���m%�3V�Τ��d�)��=X��8�BTb���0�}�A�t���b�ߪ���P3V#q޼��BF$;�&4���������a�5Ksp�"�)��݇(�����UW�.'�'!@ ����_@���������h��E>���&�mB�m���J�i���4q�> � �tP��m�d7�w���%�l2P'p�3��"��ӿC�:3�ݡ�]����pCyʔ�h�_d&��]��=#�ha���1E� �� =��G�y���4��(A�9�%E�]9�E����s�4��L����4"�@������k�7\V����e�W�X�-p,�Z<�鶣�ٓI4� ��+,z���Q�R0���_���(��Mq�w�eW�͑���}'ul�_a�������>4��شU��Q*��,
+�I���hjۇOpq�3QU0���U�Z�@�SfD�����M"����O0�n�����GԮHi` ���=w�˚�@ǘV@�zy��rW'�N�6<�Dƹ�l$Q��*�ZhєX�X�얭j�ѯ��{���,�����G��Tզ��V(?B����}�w
����00$q�����@�*�\� ֱ{�Z��22�����<�խ�v���%������Wo6a��M��lƫ_��������Z��f�G�e#p����N���ML�*�^{�j�C�I�Tz<��,~�@���wn�Z��;��Y�T ��t����^�n�{�fk�Q88�%*���S}�#�x]��B��#�w�����íE��M���*�U=�!4�E�nVB]�؛ ���`я�Z0�δ���K4��������� �z�_�gH���-���*�����������5Sl�-�ɲ2?��7��� W�AO��L�/\PH܂y�"�B��<�z��-�k�T��@���v�P��#R-�HG)�}p��,?u��4���d�q���w��ri#��D(K��O�'.s���mjG�3�M,�oG�LGh��u\7�����|��ځ�!����	T�]���Tdʩ� <E�P��8�L;)��0^��WPBPE�$Yo������j����w\5Z��k�j�M��R���2fF)�_Ȉծ���yТ@
3�z1n<{7g�	:b#�\v��K�tvD�/s�3�]��� �`��m�V�q��b���Aol���c������� ���=̀Զ&�MU�q�p�W��o�0��c���\��Z���iW17҆�l�cӶ�&�~χ�'$��o���H��Qv��>8��`����H�(=W�(���9.�+��Ƒn�XTX~6����"t�Hh˙��7�d�D�]�}eu��E3��p���D/��Pn���	}e*�5�'1��%��Y�Β�h��9G�Y?��ƂW��q�c�w�OɁ��~g���R9���r���1AB1������|�ȔaW	�f5�#�мg?P~Q$f>��d�')=R)H�{�v�esNM����h�[���CG�p�]'bQ��[P��^Bb�%#��������t�7�Z�$�p��n91����8w�zt�jq>qG���D�o7�Wlx(�Z�H���ˮ��s��W��&L�*�)�Xp��$Wf�H�f{?� �rƂ{���ed0̩¹F����U<�;W�Vqݮ�C�B���[�w֧�/��Q�*����G��fO�D�θ�|��h� Xm�����#�wgt��,�i���2���;oL�(zM�C[��?���x���Z���*��1IhT"��� ��):oX��|&E=���$���1� �FVw����[OL��݄,��ˢ ϙ�;�1��%�\��1����@!����I�\���yQ��Q��
u�>��3����dw������M�}sB ������y��8ƹ��R[S�o�-=�䨝��SXt%�Fߤڧ�\�8��/aΈ�?��+vx2���҈J�b�H��S-@���5�QpO�:6� ��P�톒��锯N��,ı`5�,|�(�5)_�/8jyӮ/j�[����Xn��k^v�����w��`��Hk \�9����l�X-����C�fh��9g�[Q��r�c�N���0n,��NKR����Z��-�E�x��E���UƉQy���N�����,5^%� V7�|�C�Ƴ]_��&��3�R2����,S6�)�H�3,偒�F3gȦ���>�_A�Z�����G$ܥyuU����C���>ɕ@=tʊ�a�IG��E�VL���AK~ݘ`�:��8�� ��䖪)ad:��؟��V�:������1у��Y*��gi(�+�f�ډd���&� ��!�&.�w��>8��C��2hͶ��m���8�y�H�K�������:��u��3zy�'Ew �mEu������W�kC`��g��T�gi��&�"	����uٶ��g�IYg}�P#K�\b�W&�M��0���j-�/)���>W��/�2ø�9s#0����7�w�0�q*b���.�)�e� �}h��mr|9-�C-l��R�f�r-�\eD�i2�H��;�(�Q���eR��q�p?��
\/+��+Jx�m�R>�n���]�]�=�o�|��w�3�k��|����X�u� ��V!`j�Mbo����k}�}-F��7�H�%��=����������(����8��0:�W��I�����/�~G1wJX��bsU*=_���G�H+��;��V�g$F��V!�ZD�[жo�)�N(�6en���*a��{���7�'��ЯcR�#�`�������wϴs.��A�\��2�'�ϧ8���I����NϽ�l!ae� ��;��P-�&(`��㔙�_.�?~@�]���*!��Di�T�y�ȉ���Y�G�ayW�+.�ΞvCRȲ°|�W�V_��E�>��FdU�8�0�*޶+�i�5W��$��޶&�^�p�_�7��(��f��#N�P$�R̴�X��wIŝě��a�z����.���3�k���x}z�����[-��Y�rM�D|���[�5L����R�
Ρ�3�vf�g��_WI����?�+���4��~Ŧ����V8���fTZ	�ɡ�+���������0zi#���k�6dd��ʎ���� ;$�&����o�i�)���\&�(�����	XzyB��L(��Ư�b�k�ɇ�QehDm��.�Pbd��&�Y���D�Z� �F�p,���ܳ�v�i��z�h#���/T��)�h�;�T��s�էP�K]gT�x.:k���ԹN�m�xD�wX��Kƴ�EH'����9C^	{Z]g���R)���k]�^�/.<��p{W�A����OA��l!�|"Ts� ����\�d"�N-1��.M���}�g�4�T?~�Y�&equ�>���r���'�2n(9�Y>��jj�m��Uh	�,��y��K������O���4ޥ3���t�-����4��vp��:L��V*�������S�bD��GB��#⿹/j��^�%��]g
w97�.C2T�>�{@f�@�1����;���.5;P�5���10>(�b�=��H�}&`N"S��������G�8��UJ��;7=X� �+�}Ǻ�|��Ɛ��Մ��zn\!����	簶��C��B��1B�u&�>��ӛ��h;D������(n^����0��� �I�a�U�o���Z�"���$L=H�g�6h�T��Xi�ܸ�d-e�L걜
�2�CVj��V8pi�����4���(�x�[.$�����>���(�(���9I�l� ���iS���)��z|Ȫ�y�x^+����R¢}���`=���k�<x!�_�y�Jj��y��R[_ϪI�����l�
*Ё�[0����አ���)j����k率����N�i���3�r}���*%�ȑ��A��[`�������J)��Tڄa�zr�&�B����eV�#\iU5,���a(��S�����8;.�a�!�ɣ�Y�c�����?[��ۀi3j��5�D�:�+��:���5q�u�'?���I�?���1)�j��WM4��H5^��ô�1�U6Ȩ1?6����<I�m���$�k�Eg���Ϋ�Ͷ9�H ��H
%��`J=�գzRT��O �M�P�P$!�C� ٥&Z��@��ʍ��n�e���?����Գ"��YG���lW7�ƴ���偰?\����[�ϛ��z��<OB��a0�IB1~Ġ+M�f��Q�$fQw%Sృ���-ѣD�ħ&FD��{�����g����aP��+����=�#��
Y�֥0��Jl=Z�,i�\w�C�#he63	mY��I�HP��y+琚Q8a�4�/�=�MW[�Zg <~�����ĔԞ��!��Y�^�HH���� �/%�����H�0�\�8щ�b�;y��M[)HE��DT��:����Ujv@+��6��U\�2�x�I����e�4�|�>2�I6�HRi7
þכ�HK_�tJ�K�ws��l��;%'�-*��P��+�����/d-iD�l!���<�d�(,�D���� Я���������s�`FB+Ã(31�O>�u�,�Axdu:a@	�p�Т�B��	P�9�1�H7%.������֥���/�?�|?���^'�u �����.fǹ�
��ZI�$͇���˅P�Ͷ9�9&��\:8��R�VKI:ǐ���3� �~&����m(B~�F�� �)Ov~iTƯy�o�w��+�O��8v̌3��)�I�q7�h�.���!B�$^���\��	{������Ž��8�_�湚n��O4I@ͤJ��+�7.V�(q�EQ�j12O����k �ő�^��qϪ��ANu�"���I��]�&�N
W���o��y}���q�
���\�|lE��V���uO���L� v��]���[ރ�xvL�?��~��K�cJh�|!TO�yo�t��)& ��Q�S�tF;͂��ڕ: P�-�L*�+�d�+}l��nCK�4�eֲQ�*�] ��k~��@�����V!���]��фŤ��һ�$��Gt}u,!}�9KZ�X�z?����Ȳ;Y�^wB�;=�}O�}ɸ�,�.�@jc��gJ�n�I���C	�����q+���}h�_%����(�C�@����oDN�� 'W�H�7[��$��N�n��q�}�!��.)-c�9=G� L���{���Z�2[ɚK򼧻������Y�R���|����90uo"v_�o����gy���J��O_�����u+M���j����?T_�v�el���߂\h]"ч���e2L0���]Y&�U�5�<`J��i�Ώ������p��b3[�d�p{�ާcg�y�8��
�M��3�yi�N�j�����`8�0^���{s�	#,�������.�D}<j�dqB�^	���i�f��W�7�*�)�QsqA�YUz����|��.��i���cڈ�#�`0���E{��L���;�4+��"����bU��_��xt�R��	��Tϥ9Ñ��v�m%!a(!zd���JǨs�	�Go�G����Q�DUO��ځ˺-/Uy��ƚ�ǀ |W�:�j ��IO	�qt�� �