��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ���������v�Uյ]�Քw��'�����u΍�=��_-���Ӑ����O��I��l%}G��$͗�T�'��/��m�wY�b��K�	h���w�M5KW
����c��[!	(���%�B:�$�Y���x^��mD����d�(����H��X9� -0F�<��D��Lh;dD�!xi�9���n�ٔ)7�n�Bf��q������^��\��S�G�9x;`��Fa������K<0�b	͚�x��ݻ���ۃ����=����]��:��f���ǐ�H���<��}�(wuC�M�ϛ�5.�d��w+��c��R����lqZ�q�'h�nE���ـ�'�:�B���$K�b�XG2�0P�UA�d�ަ����=	��P��'��)L���<H��@j7�N[�΍�÷��]U���S���b@V�c{)3z���br�5Jפ��)[���u= Ԗ�w�3���!�)n]Y�� r��WCK.���R�{���w�蝪x�U::`�6���M
Ѝ�n�m�	a�\x�&+���}�#m��
�iJ��яǒ�Y��:t��>��t*t��R��hLpcr�l$�$�&�꒚���5�����D���grb�#X�K���9&���W�����޷��I�j�` Mu��Ad��#��Y��[&�h���H��6_�
���y�WXX��c�� ؉} x~X���v�k���<�e���0��2Ն=�88'6�9<����_�n����"	�۰��&���XH��l�oEq}ssHH_���9�\�]e~Ug .���Tb����5qu�@�q˷��36%����_@��+����f9����ϋoEoa��#�29UZ��Yf].%�J\u,�������5Eɓ?����&'W�a�����0�+�r;m��Q��ƀe�i]�f�t���GB5�"�ԥ��# �ʈk�$���}Vt�k���\�S��Y���̅&�Ƃ.
���5��7�Mc���ԑ�I�:�D�r�
J��8}!~
�$Ss�1���!�`��㖃m�S�4��c^�]ٿ�@b�-U��i�BM0�e��%�7A���hAV�_py߰Q^(����UY�?��"��Qǯ�	�JqL(�Ipr��)F�r��#q")(iȋHxck+/`z\�d7;�4�;�{�"���#	��\@��a�N0�_�`b���Ҩ�ܕ�R�(9%�N�*<%ojZZ5�_�1��n����Tx`1�F���5CGK�A�+d��WCYPs��1�c?�OVMr�<��@��+�O�9琉|����f~Q�����o���֦�-v�{�m7�b��%Z��F����iU�|m}i�P�Κ.b��-��Ş�P�Iu�ed�f�0GM�U3%��!Y0Q��1:����XdS]vR��Z��ۤ�=��nR4��^Z2�~�M�6n��(uv����?������>�Pvh#;3m��2ą"���U��^!$�n�	�8ʌ������m9i܁�t�m�Zх[�vxz�Z�]#&��d��F����X�;�ʞ��ͷQPO3�i�^}8nk��gk�q#��}>���B�ɵ���}'����?�\������ ߞ҅:Ϧ�2�(5�C+���d�2�=""�
��"�y�[���ψ�թ�xVQ��x��4������1��>�j�F�H�k��twaӕLmZX�5����z$�H����Zc�z�%ݍ9ܒH?�c�a���G������=6k�#�x/��d.'� g��0����56����O.��f%@1�Bܿ�x_0f���A��bT �Z�N�@1(i���Ѭ���d�S����$� �sH���7V�����^�C!���\��a��"l��F�8K��c\�
��c\�������Z��#�c�9Z ݹ*]��xڄj���F����>�fɛzY5��u����ZW9Z�v`�w^v��	2�q�h�*�ܾ�&]7Ճ@mz0�OA_ <�y�ٞs��7�4�D��ԒZ��p��Zo���4=v
�,s�u�����^�U�@���?��u��tt ��1v�Xm�MO�QT	`Y��L��3%�4�﨡KU���5}=~7�Zq���ьb���瓶�VY��	�
V����̵���:�U�G̅N��\���Р��6wB��@��:1<�Y���O��lJ3D�z2�x������˲H.���%�ـ�:��Ra�'U�N��$�-�껹O�bc)�/[�7FZ+\�q����4$(�%�5ܒ
����a�}�딛Q�;W�N�y�<1a���S|�_�Y����<R�����`��C3%���)A.���ehMDѧG	���(�z���V�M��"*��u,a���Z�#_��)5@�����c�5&	�ô�O��}���h�{�5*;�"�ko���B!r�W)�3�l��)q��P����Ua}S�Ӛ�KXz�Ã8v���vb����N��}����G��Z�s�\�Q��c�ӨC��p)��B���9n2H�N����ۛ'�4��Z�mv�ЙJr�8/��L¶= q�^@��>���ږ�O�He��Y,��l�,nt�e���hTy���o1���*��򄽦e+>�5�ə~�E���|'KׯνD�#ME��*�"`:�h�%Y�*7�H�h,4 �mM�����^0o��i�Y�N�C�{=��ҧ�:r����&�ʄ�����Ӫ��Z��ՠ�����U�EI u)��v>�2�g-�P���wZ�8$p�V��4�$��o\iAU�^>�[Ϲ�XIX���;��9���MǊy��[­ȼ��^nG���$����~2��O��(ϋbMP��$�{�m+��Cfk��c�lҦ�I]��6Y�0�}���.jw�Y#���غ�q��9���������Pa��C��>�?�bн�,�َV��+��ֹs�'��C����)$����I�0sF��+-F�:���A�ÐU�X H��»�BP�!�� �b���4�{h��AU�����*�f򽫬�BsEeUR�80&�&�w.��v��|?�\X(���)�?+�7l"��W�@2�-���\��+B��M��7*�;>S�D�I�����(��Ly���j0���hl��Zy���J�O�c�=���e�"?���W��ıM/=��\��������H�� �^ۨ�УӦW�_<�ݶ{v�`�=o��m�����|Ʊ�EB="ԕY�����Sq*b�o�
��i!��#��^ѿ�$iڜ�i̲�Ȑ�� M�K�/�Y/0ꁡϐo'���َ<�n�壿���87HSB������q�h�'�hYq֪�/�E�e�݂�I���E�_�����v��@�����{�P��!̞N7�2����O} ������1�;���{�ʺ_�3�;)���*�AwuK��c�����_a+� ��ekm`U�����Ej<|X���� �(�����eG>��,�9��h��n��b��/8-:5�%i���A��Z�HˮT`W�A��?a0� ��q��@{j��D��m�0�v��[��V������xҏ����⠞2"�T)㭜nK�s�X̉�����5��Ssz�Y8�#�|�h<N>��^�kt�Sܠ��/Pf'�D�1�.�P�u'C8�$�_�������K�4�z6�r��0�<���`�<>ќ�5V*���	�^�9!�x�zc���Lؤ�zw��P�tS�v_SG�y��l��v��������{��5����c�2E��(Fy؟�Z���I��%Օ�	��ջg{�<�}�^cՎ�G,���?�6pf̎J��L�;�R˻x�����\�\ �H�"�u2w��uőN��<7j\_�w�DD�ys��P�Ή���(����;lZ2�@~���h�{������c+^6Ʌ��r�)�L='�F�8c�xM*��&y��#r�8���~��k�ࣆ�+���<&I}i�=�D��Yiւ��-\�t�tE��k�O8�-�����M�J�G}Q�z�C��3��U܈���!P�2l~o�f� ��i�~!�;��=gN[5Y��zJ^�=�nZMKG��y��Ɇ�@*��X�)k���ȋ�n�.D)��P����欋��ik7O�T��Y�j4��{�+_̇�g�k�{8����)�5�����6����'��œ6����'�&�zsxc�חJ\hu��@�]Q��qb�p����:]vǪE��g�����U�Y�L�8nh�W.�ol����q�X�U�BӔAd�s�"�@��3�9'x�@��s��-�#D5f����"�~�,���~4�|K�缷�d�����+Zf�=�k�2@,���<V�x}ѿ��N�$��㒲�#͈��h�Q$�rδ{��3�~/���:o�OĘ�7������\���P{X6����]-㱸�0�c��X��NHd���_�yr�*S\~B���&w�BX���K����'!�("K�㡰YU��g^���\�C�&�(*+`ڱ��ՠ��bw��$�@� ��i��G���B����.�v�gR
7�<��=Z,}[��գ�'���K�g���#�u ?�wbT#Sɹ����AX��R�z�B���@k�dIn-W�r�`ʋ����N�,���xc�EP���+YĹ��eQ��1]re��YG� ����A4��@;��>� ZC�B�Ql�=o �����4�	E����»Y��K&7̢�[�G���_Rew<o��Z�?�*�.7ԾBj���}7E�ڇp|�e�_�ʲ�ZmL�M`����^�i�Ŏ�������3m����2���(�j�3���Tbw�6��c�}���Q���}�i/�iSk;d�A��Kݘ�;6�#��zP7�MG�6_�.��z�3�7�ݽG�B�Q�NW��PMB����q�;����󱉻����ᦿ��,�g|������8f��vɐ|�-�e-�q�:+�,`p��Fd�K����,U�)�z��8�$h�0���"��I@�cִCJ���;vD�*P��8іWj�%�l��g/�6)r(���Hv���?"��g�|�
�X������D�,����Oיp{Հ%���s�N;KS��V^�<Q&�bc�e��qq�ZZ�?/!a��y�����M-�k0�1����NR�k0S��)����V��x����C/,Ϟ�pu=	�C&�_w|'Z#����v�^�TI���TBE&q��֢S<�������_��PV�?3�N��'��b�41A�,n��VJ��X�|nP05�A��������h���Z(�p3-Db�8p���~%����K`�1̾nH�a�+��� �LTU�d�;��#'�FG�f��Hp�bOw�O݆nD��-sFD��,$Ҷ̨�"<0�����򟼗/�rT�+�T��� `�HH���.>� _e\�?��lKc���Zx�>�;v��x�h�P��R�m'��O�/��&R���R.��n���;t�"�*`|x*�['��(�(���KUΤ��TF$�Ė/QԄ��X:k�-C$����,��ހ�CCw3�0���FWs�_�m�ο�nmQ���c)DE#��/)kІ�3���-��f쌓3[)K��ۭ�R| S�%%;�z�lGO�8neˊ�:���h�bd��M��ǟ�v�uʌ���8���d[�����xl�<
?�ؼgc�М�{"��DF���#K�{�#�)I&3I>�o�*�V���I
+SKne��/������Z��hp���1�M�E6�난�_R3A�Y���#��Y�;��d��5x�M`�н�1_��>���u�y������4<6���t�R�/D�~��%QI��G���;� P�ܦ8�f��Ufi�Z��*JO��tR ����=�<h��2�<WY����?�y�U��;J�yC���������MSZ/��!?u"�XZ��d�d�J�DO���B)s5���F��|�auDЁ���\(HL�FT��3U��7� ;B��[�̼�a��4��mP���4���}s�;�?8.�Ҿ �N�Tɸ�y}jvYW	����)%Œ�Jm�Ly;���ƃ����>x���S篯����j��LO>0�X�V|���"&ˬ{5;%�v˧����8��4�&A�O���@mݭ�\�U5Z87��R�crd-r�>cG7p� $ڇ��`����
x��=���x��g'��$���|�Y'��O�~��e��X������*b��G� �Vy�"u��e��p.E�҂g�/w��#�۬Ў�����ɂ��0��?iS� �����ѐ�������E��G9Z�3>?;ʞSġ�	M��֊ 'v�M��fuQ	}\���5﬐��ؑ�aؾ�M��{��MY=�`�NRf�/A��H�1�H�$���"0J�#s�O���Ke�H�z
�a�h�H2�Y�ŕmߑ���r�9/+��T��`�*S��D]�Ca��o<�QYYV��\;���L�J�V�u��k}R
�$#�`5��J��>	���vV#�ԃխ�LS��\��aDh���?��{�k�`̂�!�-	�G�)%uݩ�ӵ�������F��v�˵#��dF�}��Cm64Qtj���2����w��1-��b_4���5̎�z}H��Г�{ȵ��-���>Yd4z�"���m��5�p�MP@���M�Xg����>Mv��H��P��h;��T��@qx�o���ľ\4�����h��m����.����^��!ms��S��o	)�p�ˉ�e0h#���u��E�3]�OO��C�$2��.O��7�J
����L�ĩ��� �W�qڑ��,� ���jN]�����L&�0A�p)	�t���@�o�ig�����N��wH�q]����s���r��ȳU�>�d\�E�J�>fAMT�O�a?��i#|��:�0����Rx���py��l�4ϩDW�t���8�N�y&"��i�;���(��z���/dj��	�Yi3S*%���Q���ܸ��wG([��[�Q��n_�A��-���P� ���_��N�m}��� C����ëw�e����6@�HD��/9�ݹ�:2m�ϣwJ�#�n�N��J`ѐG���H���gDY�!;�C2Y1�Xjb�c�Bn눫1���7x��G^�'��u�N�`Z���f��.x��C ��5�1���}�YR��h����.m�;̿�:���8P���P=K�\a��{a ^�f��z0��<`���t�X����&�y�t�j���|�Y�ݻ�J]��D	{��Ɨǖ�/�j^O��3�ްi�0����7�A��W/N3�3D�/.�^�4hg3(�f7N��z-�
# �ն��WW*('0���J=�k%��^-�1T� �mM��zA6��f���v���z]t��`��(���#l�&V�D+Y�Ȗ#@���%��be��煤�Ѽ2ӧ���'
s�������}�g�f����=T��l �Vb��&u���x�r�6��1��5��8ˋ���Yt�+q��"ܖ���#�9PXk2�f��&����'B������z��0���A*���
�`y�>C��ޏB����~��q�B�R��C0'JO�T�aM�̧�v�́�v�B�1̀[\(����k\O�~��P�|���/R��r{��W�(9�mɜ�>Q>l�q�a�{���<=�y=0/������aOw�f �|�R������4h)��;�#:�M2�K�N?k��k��
i��.����0�"��o�jdx�҈]�d�t�����#F��n�醲���lc��3���s�7&�Z�N�G9��nJ)d�"+�lԄCWɶq�B�v3�����^��ʾ<e]F�]�LKare��۶��y��.�j�|�}�}9�����!ݫ��k�>>��6 nq��M���6��&��)B�g��T����2?�	���i#���0�UM9�m�k�g� �~�N�Ṕ�H�T�G�����2$�և���,Ӫ:KO��j�d�	4mN1<:'��s+v0���M�V��1I���]�XVX�Q�J��.�c9���Ǽ	*D�v�k�s\�-�g�����q�h�>>U/m��U�Lj��jYz�oCN�������{^[��oT��7b��U�+�����O��Oۗ$��E��#B�}��s��m�N:7�«�'���	��,t[� =٤�5 �eW�{�8ߓ�a�;5�(��K��׈�V��t>|9ؕ��KC8��͓u�'I��;#M��<:jǉg�`	IbW���te��cX��`D	�Jz���?���T�fh~�n�)pv�+�-�=�ז��?�O��~P�����y�\$���7"��F�3+�K�, 4�mdQMV������'��+���~��)�,�D�b�s��K�D�o���qD*��eO&C�2���4r��C�$9&�wF�j�;{_�p�<k��)7D�r����;r��5��g�f}ۄ�i
J�,��1����T.Q?�i��,&��!��$v�;hy`?��䴔j���Q��/3���d�P����
�Fp�Do�Hn�?��Lv����!6Ş��A<�HI���Y�㱊�٦K��x8���0Gi��jX+_�i���*Ex�]ټb�H.Np��FW�W�'tcε�_@شS6Ħ�`FcM���=�s��$.��N��B�Y�������o��('��&g��iyՊ���ho	���2�͌+9��T���s��Q� �����Lo@q��	��Z�bF)�!lج�B��R����¼1���N���&j��薓C����^��-
y3��IF\�d|D����F��`�B�n�R:awD��¦��.�*"A`���`5s�2�"*�Ϲ�jk'egP�}\b���*�m���9�rY��=���V}��<c}�#�#^�ՉM���kt*�{_�+�>XGlC��)���r���"��a�O��!�r�w@�K�!�ԣ�<��_��R�"�,%{Y��^��GKS��-���:Um��q�������O]`͙}=99ފ~�פJE�?0�y�"�=HWެӕ��}�,�{ꔡ�ߚp-��Wv��{W�)2cv��k��hf� E�����:9�� l�uC\P�[0��뀅<��%��:��Ѹ��ME�d�c �6Fz��a�QG����s�6�'�W�x�$��lKډ~'���e,fq}��D-���m��o�ӝ�@�]�I�����,#^hZx��M�����d����Z�"F%�@n��H���&(�&�Q��r�q<t���m���^�ET�so�*)e`��9�k��īN�p�&9��#\���pQ�&�(3%���)���q�D!ib��6�C5�׽\�6�ی��+[?/����ye<p�֪����V&�(���Z�Bu
N�~R
� \�2L?l�4�!����-99'�F��k��7�6>���&e�ǜ��V��Phj?��7���@�UUҜ3Ɗ����	���R�5s���xM�+��g%O�Z��y�c���G!5F=d����QZs�Ň�L���sZ�*��/z�=Z�7�|}`��փW~"*�*o������B�2r���G�c���\fK� ��w�n�.Ps�b<^�I���0�Y�I����Fy�6�<b�����g��0�ކ��r���I��5�����h�g�È���A����ѹ���1��Y�N��h�Q�c���"�����%h@���iS�u���|~)'����N/�nD�Ő���Ӹ��KR�r�A�bP�3���g;K�%��{�3����Ղۑy,�2��{Ή����oN�_�M����K{q4��3}�L�Im(4�>1{GW�7�.k��Z2*�،`���i�� �����PMh�����kHs����y��[	!���U2��_!I������i����V�F���0s�..�N0��S�ɴ~�fv����O�*��/WÃ���l���a���v?���w��r��v�C��3l�T�U����22�=D�z�9KK�[ �_�O�h&�DB�t&A��Wt���ߧ�
@��\Ns������u����֬�F`�\_���g�*�aa ��ڭ���]nef��(�y�D���s@������7��LOWK�.U�ӕ����+�>8�\�u畦���'��o�wP��O`W)�@B��sI�%�־��O�D=�Fy�z%�����	�c&eڋ��xG�Y�9��jg&�7�WR�5�!ID|6Z*��Mh���{�,Ne�յ{��mܹ��2�mz��QQ5"���; ��	^�nr�U�,�;�?�_cB��Z��+~a�ʸW��]�w���#0���o��Qkh.!�����Sh��	���!����T�?39���k�F�N�߅$���Z�4�.���**�����y>PA�컟 ,!�C��K؆Ki����
*L�e�ne�i���o����mn����b��� �eo��]DC��<�����,�y�F��eO!���m^W�S�da��Н��2)Xt��%R�:d�KO*,��J@�������0h洧7[��!0-M���#�Ex/�S�_;�Jy�炶O����?�[h�8ᚲ_
�}*��4�?C�臌�Tݩ�E����"����q�� ~��t��f+F���O�.ħ���}_���H%�e⏆�W�ۂ����:��'�_n��bn_r���UO��+H����Q�-�ֿoE��.��IZ$j(�jVrF!�)�.�d�v�v�<�5�I��L���^��s��T8���{'Oۆ1Bg�=`5�FP�>�S�I�)>������"ƊE��U����I�6΋-�l-���O!=d2��%�d:4�؏
7`�D��c��M�����0" �����Z��
TQ�ϳD���g̛0�a�nwJ�)[�x��U�����f�\���T-�t[8
����lӶ�-�TlX�'��hj��JAa��ȓU�X �i�*@�u0������}�-�r��%�`J^)����o-Ar)��TE����:����ѩ�Yb_��X�j9�+J"�#�I F#b�BB�F���G=xA��o�z8���T�Y���Jz��Off�u|p% A���e����4Ml8�К5���e��\G�T5��W��o�--	6��ym�,�CV��"�w�
m��nY�Z�Yb���tl��R(�B7��C"R�8�UѾ0@a�9��~�����dٱE�^O<�6B���� �d����_I��V���)�p�΂YIu-@n'60�,%��+�./gz�j#|�jacz6?�]N{I|Rb��xd)�~�	!�n�	�^HT����٭���e��C� �CW�4D��1��WrOg���o��Eب�/zK���B��HV��wӐ��7��$_�~�1Σ��?���]ww������fs Uf�#WlG*���{$��S�p�d��w���C�bP��`>Qo:�.�X?�aٙ\:�'�]ds~�T��������/���+~�bMiu�?��=��s$}QH�}�G�rW՝.��8o8係:�7��U�F�#�]5�'/��o��q0«]4=ڈ�0ف�l���f�s����CЀ{�?��s'���A��'�q�����kZ��=��0����lXt�?��:+��$�D���Ҏ!��n����053Ji�aw/��F���5�HV�pt��B�*��4}􇱑B�T�>��7]5�J�j��z�z�k��'���o�.�s=M��e�mU��N���S�0(�"P�y�К!��3�EH�E�H(fY��M�J_샿\KESUMyBT�T.[֡�|�>P���r<�7Vtx���GT����y����L���p���f��:��������\1��=j�@'�5��%8�t������cE��w��ۨtˁ�@>�D���Wѡ[~qkѠ*:�-g�C�k����8�fƦ������Յ�Wu{,L�1�E�Y��
e�W%B?m஻�y'b�G��v5
ײr4�;�q�~FuX/�}�&� ?Օ���.�5|�>|Nn i2+w�Q�D�ѻ{��a&?���:��]��׉:qf�kT����+��1�g���ho�ʹ�]>I�?L̡t�����G�������7=�	��+{N.w��؏�a�zϚv����"�sVK�M���$m����	&�5���bԿܿ�x�}��rz����63�ɧ)I���C����vtV9�%?�c3�PL�U<��@�L��$b�3�2����a��VL�R%��Gu08�1Q�H8f��GӚ���2qbP"�c�l�����o8OV1�_`Bc;/Gl���-�S��{Kח>������H�������bm�FGN��'{L�� �}�:��}*���I`�z��$$s���Z�K"I�e�3�mw�xQ�=/�)�eG*Re�Yb�i;���u�=ejͱ����8��E���	i"�s��W�x��Ty%���;|���}�Q�V�D_���h3��N���T��סd��pP�X���n�{�w�+ȅ�Y^�d�xb>(��Y�Pr���|y	�J]e�N��!΋|��/ȠS���,����n�d;��8j)�3�~`�$�  Ru��u��R��h,��[�������O����ě�NL��έ�K���mU�5J� ����u|�%�dNx�G�P��eߙa�e�e���?�p���IK��g���������r@;t4���[�)i�Y>�e���4ϲJ<��)c;�=�f�T�q�� ��јL2��n��@�ۡ��F�4�9YLP�U䁞���K���N@>*\E&��%��?	��O�SV�^�d���������5��lOC]��)N�p�D�Qn��gg�S���;BԿ,�]�k�R���R�
�'�xԳ�^ً`�
+\�]�)82�V#�pF:�4w�/@v�@c0`'�A�A��S�:Lݓ�"܄S�C}'"�6��Z�(^�n9b��@V:�q�k�B���#:�RV1�G�7���Z ��d\Г�"T�!�Cۨ��s��Q>�����!Rᝒo*���M���}L��
��"��� 7�y'V>u��tF4�u��zQ��([��[�9VP��7�=�-��rF��&LM"x��w��{S�^$�+��+K��q���n.h���Y�$�0��30�Qcˉ[��j�5B�ʯ��^���~��Ry�G� �*�N��>�K�����ݷ��͖�/��2�e���v�e��S/p^��
���,�����mR�[��0�bT%U��=�SR�)EI��L�9۴�U�����,^�բ��-�$j�	�"�H*r �]�bK�7�j��h�1~E���-�H�z�0r�4e�U�>��_ѩ�(��Аw�c����e������S����:��h}���yA�"A(V��*���3�ܚѐ=
�A6$�N23�kSW҇�h��+��5�C��V-��ng,W�1�E+�������ہ��T��0��K�Q�� �y#0r_uءwĈ�0��+�Gh�D�jH1T����־�)��'�s.�7��F:�&��5�=�A��@���� �J�%E$##/���Js�\�#�`�������q��7x`�^3�V��Z�mvI�e���Ua�M;;1�yZ���R��O��>���K=@X�|�Sv�(#S� �jz.��)|�Ǔb�O�/�d�3ͅq�MI�w~UA��C�Z|�&�VT��`�~��w��Õ�
�lkģkOR�,�	�ƣ�*���ȱ�n/�I�?o DL��@�'�gp&`2�J�˶ RK��3�vе�Ff� �Z�!���[��߯D����ؓ+<l��'4��ZPU�8|F�`3T/�pw��b�qs���O��_���J���Ax�z�����B�_�P��ަ��uģ�cYW�Dq#O�]��k�25
ֆ�f!�n��R�Y**1Q[v���ż5FHpBH!�Q�pbߣr�z<o������Y�B��T�C~�	��k��� �o���gq�b깜�m�H�����^O����A�n¨��窼~�N�:U�ԧ��&D��W�qW�7�̥ظ���I���N`K2�y�q:;S0�@���s��c��������X����K&ņ��/���j�G�蠂F�j~Mܘ�Xr� ;��]L���şH?l%�9ӄH0�qCP)c�x�i �~���R����m*.[�
���4#V�bޒ���}>+9�w�i�Ý<)~����q>�b�R��2�N}����3�݃n��ۃ����v��i��������\ �+�q���XZD� G|"p�a
5מ5)��(�z]�%(��ι~ծH���:@/�!�h��q���G$���b?<�$~į�y�ڰ�)
�s#��j�,7
�-��|��*i��=��~r�8����G_3��'�*2'ˀ�G��:m8(���V������u�>��U�$j��#'y��ľs�Ǡ�'�SE)A�����ۗ��/� ~�}b�U��)L�?��n���r����S��}p��@�6Ҡ��X��ue��M�Ux����ΐ:��(�$D8���B��!�uiu!�����4�� F��d��zFv ��yu�Z�nE���g��OE�W@�Ш������(���R)*j�+�s�9����.��g)k� �7� ~د�m�|��W�����w�甭Lk��6��mw�i�q A���ev7�k��q��n����*\������ү�4�$h���L�����T	��	��=��-��g��y'Y�,�F9E��ͤ��do��!c��P����h�|���?yͦH'�}G�ѬIUj��Ԍ��T>C��	L_Y��)ֻ�H�I�8I�(�N��[�]�a_�?�rʘ j����T/���ܧ���w��@X�F%���ee��~������cON�=�G��p�0�pk�˲���1�
k�P���u���=��6��l-S|��q0Ɓrk�>�J؁;���eRR�Vm-��BW()(q�p��e��>̚.*��Op��u�Ȍv��+a~�t�Cs1b֜�N�uԾ���m��E���-��T��"~E���:���V�/��c+F���.hy�v�$��ȫ�8�o�3��$��|C�H��Ȝ��KɺR�'S	�2-��f�r��<�F����}y�R� ����e�R�X%`�e	<s=�p~�	�b�D�/v�{�v�*�@�L�<a��B�2X���Xn�ZzM�b�]�����gf���[Y"�k�@,g�ō/EI O�\Kb����G�$ж�\�.�L����5R���XY^w�đ+o)��ߖ��D�LbD�]1JBmt�G[��s�»L!C�Qܛ'G��q�8�s�5�i����('V����葏�F�WN����ޮ�,��s��P9��G�D`��J"�s�da�����=?F؍��/q�&޿��>�gX�j�ߢ5�E`�),e���LR!� ��N�����GuwQ'>�b��*�ϣ�zmݢ+F���^�ƕU1����)��X��@U7���!WuM�Hb2��7�$)3�4���dne�ܿԑ����K?,f��������1�}�r�|;j��`W�S(��]"����},+�\\;����ZBB��u���~V#;V�!��x�-^�+�䍦o+��il���zb�w]�}J(�0x�mV~�WkE�Ɋ�lRL���(ķ��;��n�ܻ�Y�FzB�S)"b\�{4� �����Va{��+-,��D��A.{�̊U��-�:[�r���vSy_bT�@�if�U�ɰ����Ї&�B��A3�|�!/>l�9�j<뽝�:N��溃��/(� 'H�h\�Y�'��⠌c>Cv��
N�{�c