��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ���������k��+�h<*y�N�vFY	�@"��-�:�Uؐ��8ʄ5Z�B���Tf�e���}Y%��D�UK��%��=`'먪�����GR��ReY�(N�h�G�5b�؝B��:W|��.�g@�z��Ё!������9H���L׳<��\I�azd�Q�1<<E9l�"��D�-[1O3]r�x�7�{�j��R��J��,��Y���<���--ƌ��]�ؗ����0>&-��~~ ��ŷ�)<{�"fV���Ar$&$z���-Ol���5���B0� �$f�����i6N�U��nЧ�<��7�a'���f�[cc�]�R/�e$�>K��ƍS޵IM	*�7fl�豊ͧz0Nu�PL��$V;'�O���5�C-���l��7��vw,��e7��!�˚@�����V,`�|�z"K��Iw�V�M�P+�ۜ�Y����@���T�fnUG5���%^.�H��~���!�y��h����jGy�x�&��"��t������`=�c+�p��~e��jE6"�e�����3ϘV8s���{�7yYނ"����ǯ\_ffAJ�!P%�DMNW�+����⥌c4/*2��(���*�y��{Z�2���.m����~��!!�ݿ�wX��%)�op:�a�����)~�	T��k�$zhe�nZ<�������������֟��0����>�8� ���zk���;��52�[AD9�S�>��T-�UᑵiB�q�8�-�}{���E��LDk��ۙ���4�G����A#����>���ݡ�Dw^P�05A�x��ENt(N"�r>�i��%�>�����K�)z�h8E_Ka�g�kV�zz���g0���Y&��Eێ��賏%�V��	���\5
E��x�����-[�_Z��,_��e��ՎA�ai�i��J�Q%B`cu�%/�D�_o��lfqt0�٨[��]Zь�� [������{4eGXu�e�Z%���V���y�y>��Ha+�gx���o�Ͻ3N�rBux��fa��i��IcI����3'F�:M��\=(#���1���cU���@��ܶ����8:]"G�(P[�ӡ�����}
[e�M����G)�!��M��'�d���:���C�ĞR���u7�n^"G���I$����iڰT��,��~��p|z��CO�rn�/"�Q"�����#?8��/��E�þ�Z�`٨�u��q���y��J����p���	c^ �*>��a�TE2��B��W�2�^�t����I�$V5"PJ���+�rk|�F}Ix��L~vm�L|�����k��)di>`��k�_E�Mb��\.��zj��P��<���������O���������!F�
��s�As����5�/���~�A_�ņ���r�'S͂��*�]��O	���wV��4U��Ms{z}	\-�j��� ��4.A�1����d�@D�����a��N~`�s9�jC�x��!$���/ї���5G޻���}�4y+rc�t�����R9 _��%�����=����8V
�nIP�<s��%w�b�]�=2���}����� X�0gi}V)��R�P�g�I�Sp:rzVh_�0���P�S�7���n��SZ��9Pz��x�_�ɧu�w�|��D�4˅(R��S��\3� ��0�Xp����k>�.����F���, �)��w�]���t�&\o�~�lH�����3��X{��aIҿ��<�Uih���l�|c�~�����5��l;�|0��;c��j]���!e7�:�� ]�4�6�ێ5����v7�]�c�Rb:%z�i
<�$�M|�b�]��{_�Đ_���0�A:�e���Sy�$�Jx[�?0�d��J2&�<��s���f�"!=�ew�V�em螰h��)!z1�#����1y�%��j
<���^bҺ}�������J��#�ٴ�w��a�Ϭ�ހ0O;���.>6��#_�l4G[@<��kk�|��Q1�\G��=�k).�-�Z	*n	�"�w@���]����Y�B���4�5�w��SN:BgM�3��J����[{wv`\�$��0r0���yR���9E��=�Ң2{/���� 6�M�X�4�5a����<Gm��xs��Ic�-R�D<x�Ӵj'����֤ ����~kZ���U;�~�s���2���!�{	�h[Ҍ��AÚ��,|�J�`�Ԝ�k>��y�u��l��΢Ap��vD��N��$��+�T�z�Ҥ�q����ڲ��A�1_��-�(t%��"Dա`�0e4d��baG�Ո8 �߻W��#/:�[3��~@��#�ړ8�Wnxʁ�rs�Ym�a�lU���:�+}���"�V|�h����:��^q��rQ`l����_���]�j���,{����f���/L6A��܁�|ir�c	^��k����,��,�<N�� �2��7��D8����ķ�BQEu�ȷ��ѫ��Ʉ��|��a�/{�M2���rB�\4�Y͒cajG���6��2w:)�_G3qy���+���ه�G���q}�&�cYs`F��Ť���.*Y���S�W�u�4����HY�&�\U�'�q��79��x��jW(��w��ن�?8Zǲ�)}Sy��P���xQ8NS6/5FB>�̖O���1�m��{d�oϲ����Ǟf���5��)$��r���%|H�hn��e��>�X�?��a��l0m�l�8$"`8��O���7�I��:���)�/�]�bgٝuk��f����bC�ڗ�e�g2��jk���
H�_wqI�a��~%
��#��5b�=��H���A��\�����m�|H[-?����vL��݆�w������A�m�Jq0@	A���k��p6�jmfv�����H4'�Q��,3�������e��ؓ�8��T�:S���{I@�"|R�P�ؕ
R:��C���ҳ��!7��k�٪Jf������R��8��@٘�EY\GS!
ڷ��#G�/��E�{��J�9B?��4T��� �V'C�Jd�4LX����HB�Թ0ENW�2
T���#rWa�G�<}�<�w�}��-�e� �F������$c8��%��ѻ����IlhV�{^�\�;��n�a^�N5����ö�dXB�%
�7�.O!@��1��R�c��������XQp>�T�5D�W����t�o�'�$�'bv��S��N¿*���ð�/��1h���0t����&���[{m|�����R��U�X}�Pag�U�_�=���Њ�*k��ժ��,����u���͘�1�^���s���Z
ڼ9:.����Y0�"�������B2C�}�5�����9�P�z��YHA�Z�#3���x�S6����5~c�<ڜ�3�{��~��'N4�aЛ)��z�[��S���*�YF�c�����fwN\?E�����'b�-Ź��[a�\��wkƌ>�R�oRI�Y	���=brD��-e������8��jm�%��W�h�J^�`�Q�`Q�g3�H�\9�3p�
U�2`���I�i�v2����Ԟ�>�����4�C��6�?��%�|�Mڶ�gy�֌eC��xY�-���7{�V�IΘH
�e^�dt\h��vS u3 ���:���@, l�`��J�=G��r�K�E���S<Z:,T,$�*yT
�G���G��}s�DO�.@�NH5d�e� �#"��D��fn�O2sU@V{]l�_C<ҧ8=�9��+Ǜ�ޗsw.�rƯgW�΃bBQ΂u�y��M<(`��Y�U5F�̔S��g �f�7��YWmt�
a���|��<�`p���'����G,�/�8����ȃ@�D��^�����8�@�?(ĸk�A��c�ݥ}r�[�]�t�J]��nA y��ß�F�*��y��R?]xL1޴wAfE�#�́
|@k��l=m���+,��]�3�ْ���=cR�Wj
F�8���Q�����#.W��ދ�Ϫ#aTQRBw��^T�s�(o��u�X��$�̿�\u�a���K�1���ml��:�{
7�p8�=A0�풱�z�A��p��):��ޕ�������x%ִ�=�CU2�on6(����k�*y� [��"]���y�y)�i /�Ǟ�6��IKW�1'|��Y���$/������.O��
O�0Rw�iD�Ǥ��F��)ʠ��Ȑ	8ˆ�}��[��ۘ�F��l+0�ڝ>?'�6�i�� ��߻�ۇ�T�`���3�>���.�,cU�f�h*K��ۨ���� 'I%x��ك�8�#��yo��<���.�t��3e�v�u:�v���$q>c���&��L�
�[ؽ[]k�0Y�oܕb�^�a�DQۆ��`�K��"�����<&�'1M1#R�}'�&ѡbY�1$�v	��wGHe?C��'��E�ȡ4^A�xz�~���/y��3 �+�3��+�����C;�����
�}�����jE+h;�v7'(��8�V���v�=ɒv=ԣ�q��<�5�<� 2;���n����K�w	a[JiɥX��
�(]�V�G�3�fܐJz��C��Z�i]$����*Φ�Y�)�v5�ϰ�M���$��99�	l%��ޤ���1�.�@���C���B�ʑ`|���Mg������}���8���h���^��3����^�v7l,_�6�������ޖ ϧ=�1��R<w���O� �F�����Sg�]�S�����d�?��g�_�	Q�@%���r^���kxV&]	��GO�*��H��9��>ά��o��u
����j��Y"�I �-��-���� A��p����Eu���E�y츚�%��~:@�6Hy^��.�i��;�Aͨ�u��Qt=m�s,��!+F��!-��C��za
�Q��&	����DQ&�~h�%`Ty:Cqǧp�R��G\��m�Y��������bڄn@}�?�0h��Bh�Ö��
�u�l*Wp�G*�o}�%���>�(����7�l�8�KK�p�H	*���<��0�UC��
U+���8߄��ִ�(�H� I��D�W�N��_�ѥ$��j�V�0�7����eI���O�
�IJ�ͤ���>�X�P�|�U��ב��(fd�wa�G�ү��@Z��6���V�*�D��Uf�L2<�y�v��o�0��߯��͉��M�XeÓ�d| &��pޘ��O��k��_R�^*ڲ���t`Wz
��mRz)��4�����D��wS�AA���%���Ǯ�SӪΚo�G[IE�[�|[���Ll3�^6:��Do�,Z0���˱�'z���YA����)L
�,Ѐ������Yo���ov�:��TL m
�D��4�#�Y�__�̫�T���fс?"�#�#�ݓ��x�;E��pi�'�ͩ�%��}F"���Ō�bm��hh? ?���.V>��"2>��������M�i�O�!��:فh�b+�ܻe�E}S��K��J�$	[e�rȫ���E���W�Yc���暲�W��o���a�v�����'����6��Ԁ�0#ьf��U�1g��KҖ��;���z�����z�����Zэ�^f�dq���߾��i�����T>l�}
��pA�dm�)�%yXf�S�BW	��	v��'��8����WX4���֫��REВ�L+PhK�n�dE�>��E�$ߝ���� ��ʿ�5���LsLZU�6�am��=:µ�6ku��v)�|
�B6[Xc;xI��P��B�N3���
[���e@u���a_�h���J'pe��:�i����J��\�o+�%�̯�H7��|F�C�y*�	+�.O���+F��_�]mζ��gMF�����wNS(�$�8��BL�Kz�ѽ����J��"�Hq'�%��Z��p���6����BŁ�	�ɣ?�su���8�6Z)�lL��x�"n����UhN�V9�˴�(L���C�@\�gr���wM��f|@#6N�;&��>�!Gy���6�L�c�^Pm�F¢��]�_{�?�V�#Jsvyb���0�Y��u�r�[�&3���U��Eo��k�,�4�d&)�_�l�$�D@�߇?
[���q���.J�aX*-8�+��g'u��L�Y��K�*�n�m�p�V�f�_���-�
�r[	��8���/�ۂۿs�6O�(c�dC v���a9ĉ��C������*�ե{��@
�XN3�P�y �-f��U���bߏ��Q� �w�*j;�;�L3T^cō�KX-E[��v����������}BId���@�M��-�Jj����a�3�>|gݺ9.��l��	/��o��7n��b���M1'���s�i/Ƕ��6���m.�X��~D���0��(��Ȝ��yf�!2GӱolWM��'�pʎ��
7K���L�*�˃(5*�0�qeC�yJ�&gH�����-hO��jN}��\�0���u�S㡽*�<`�8	]�= C[w��*�0l���?��~h«9.�y�ȍ�x[t������l�\) c��Au��9�S���@�i�T���`T_r��l���,��MV�+��j�X1��/�`��e��_"e�^�ݛ�)&�w�1'â3�N�= 9lw.`B��L�����T� �E�I�"kXڳY-olI4ܤ:�vM����@�%�5��%���Y#�����Nd}���鷃'��X���@�����_�Ġ�'�$'ȇ읤n�X�������!��i{������KA����J��� �����!$#��G�$��%���P����A��7�`������lEx�;D9��$,���"����nͲ��i�5��A>����c1�Y���_�t�I�xn�4��W�x����i����d��1�%$��ߍ*��N�j��yK��no�M��(FSk�@_VK�|{���G|i�f�/���,�z�kk�?dj,�P `@�H�)�]����rV�<�u��� ��I�^��Q�_�wp�n�h�i"稼�D=:�$H[���MT���=�|?t.�^Ob�����nd
3�N��*�4�V����a'�[�1Ŝ�O��ɂ��)5�G�j���UN��ό=��;E�,w�S,%7By4ܩ ��bX�#P��|3�B˅�9�E��Aj�e�_�×��Y��8��9�(xN2I4��ihu�Y�&�pi^.q�+JMO �1e���T��N%�j��L���%Q���|����t�({��4������	b���˧�˓��o3�G��Z��d��X�MV�5K���W�w!0w@��� S��f��2�]�àʷ����#/�J�X�,�1��3]f���|T�.������a�ǵu�.z��{�GP�,*�"vkzY��m-�߃F���k��{F�|�QB��<�=��� ?*Ý-���/��a >w�b���q�^ȧ��������s3��L~���7���UN�
k���� �,�ƢAx��۽��;٨���s��i5�스�V��y޶3Ή4q����gCM5�ّ�*�ldz�ݨ��G�v������'(�=l[]��y��@B��"�O2bR5�P6����HԝG��>CKC:\��`�ۤ%S���ojj��GJc�!���G���`�m��t9_���q&L��
Q���BRʆ����p�sIV��|�+4��N�D��s%�0���ڛv�/o���Y��G5�ABžaW#�0m�\��A����f�b��Q��z�X�������������&���;���͞����3:߬�"��W�ԫ��NC[mg�i��Q�E@I~3�ݸ�Cu6�S�k(���F9۩B:秭+؀7q�Xs�ȬRD��3/��w^�sTi��]v�'���(�0�%r��ɼ��J6���JIF"�c�������ġ�_)uG�P�sѷ��2��r�n	����`�e�1*4��ޖ,�kE�\�)����1��	!c��/a���A���χ��+>Jx�J�
=�vs�m�]�9��z9]��m@��2l�����n��~Be���r0�7�SZO�Q�� �'SQpXHW4l*���'�G�|����*�P��u��;˺G�뻌����=�ba�tCɲ��x�C�J�
�b��X|�Ł�A�S�;�hY@�%hڙ�81��Q@ϱ��Kٙ��k)���z�������h�r,�GB:�Ï��ñ��T����cVr�\q�RwV0�ې������s�b�B�o�C���VÊ�l2f�v��%މ���R��Wi(kfW�I�G���Ե���};Q:�R�6����6�J�L�%K�O��2I=ZX04� ���d�P����*ۡ�^yz����_�f�C��9��	+�� ��e��{|$Y��Z��g�62Pz�ϥG.���
�5􍜾)��s �_��Aj>U ������uMb�;�Mm Ur�ј�o3Z8��g3Ho{I��a/5���9$�6�+¶�A�*��
�k�2�篌�|��H�W�S���e��
��É�`���{�q�ӉF���_<Z,^{8ZWs+ru�/i��Qw���p_L�[��q�^o��K�(h$P�q����$6M�F��XyT��T�p���O�ح��<$C�yl��1��Y��)o��=+T���N��k�W�3Ddn�g.���䛱҅l�O,h����n�u��G.L5)�Λ�GD���
O��U��YM�~�b�����)3$�Q�h�+_�2+���z���dL�+��G��0��P��� �D�c�k�L��&����/��na���И-�}ǂ���@��L�yNР��������ȼ�`�\��K� 
�K���c=��T���f��SG�q�m�t7C��Hw���Ա��F����%$������֯����m��ͬ���o�a{G� Rw^5]O%�sq1 ��*Ӷ-�!�c�Tg�}ENnEpf-;��hK�c�VX[��/yg�7�����N˔�kDP��Ц�;\�k����D��)�[X�m;������(�&��}g7��'�J��2���p΂]�n�4b�_<#������B���N��6�ڣѺeN�	c%2��&J������idڔd`�9#@[?�{E�Vo�D�Z��I�s��� @]�Gfs9GP�}tIE�:t7TK�Į�����*=?蒢�0u�ʭG`�֢k<zQ���cf{�L]H�=�B�Y�^W��m\l�`��7)��^�]ո!2b���Q��gJ�;��j�Dz�T�؍��(�Zp�f�.܇q��jO6�%Ɍ�,�P�X�������1����.�$�F�<�h��-�Rْ�ʷ�`��!JdhR�)o���*��� ��A>�koNT1��2�v�%��9/��(��G)tKUF�W9{	}'Y�i6�O��?xp��QW��a�?�m1H��)���d�_W�B�������ܕ(�RT�'Ҳ�߫��Y�n�*=#�f���=��ʯO:Vμz����S)2VN#
3G�F^n���PF������Dt��G�Ђ�Mw�Ǩ�Pw���������Vbz4
.^�ZAY�\�7��6���4�ֿm&C���"F�͔-��:%�����3�La�T&�9��sY�&��U�Dg��� =:����z����Gf�U����Hs	���n}r��#��(�+��^�����0�y�*f���l�0We&��;o��Q͍Yu����a=�:q��+�8�-lM���fr�$P�ZY�}GW(��J!�'�F/���K~
0��S���g�Z��d';�Y����l�p���b�F�$�`%Θ�6��}׽VOųI���3��ϴr�����䀻lօE9]n`�}��d�3KČ|���^E�D��LK5�t�,kaS 0µ<���Q̆�B�(`jdm=_��U��>��t�P��/w_� VZ��=��j�,��+a���1���`�~}�\y�m���"va3x��Rͽ���3,�G���ER,?wߠ�Bo=jm���X6^��U�O�%�"��x��>O�n�����JU��
r��
dBTԇ���3a�`�+O
u%rs��t1����0_�.��qL��g�s>���Z9D�-�|�����s[<�����+���+���m��7�˳�����d )xz@
78�]�S�!��D���o?&�.f�d$�"�z���N;{��ج��39��o��s�L��P�":�ԇ8$����'#����;}�m�U�f���V�v�H�\+L's-<_�V�宀i9��W��I�$�t���NK>��W�X�dZ�AB��l��
x#u��� &x� ��,�����A�oI	" ^�f�K��Ep��y ����8���A#N� U�-B�b�EL��{V�TpF�Y���=ʆZBE{��6�:�%���ʮ��i�
��	��L�J(��;�N��%������; �-.�o]�w?:�b��H݀�{�m>g͛Ɍ$����/�\�ʼ����*���_F�u���%�S&5g ��	����;/��Ӆ�@ґl/gA�{�)��2����!z5� C/�ߤ�Xr[�g�?�c�*��ș҂�lR�[���p��7��A�^h����l��ewV�v�~N"S995��l�3C����u.�h�����ko��Ɛ&��@�g`PR��� �ߋ�\�����0�����c)��.o3V�q�7�}��Q��������E�|3*��hX��H��cO���#�Wfj�T���!1 �-y?E���iMP�L���u��5�{����ɮu���9lC����]��ъ_�-��ř��2(�n��l/�$q�"(�*|�w��	hB�XgC՞��H��z��_�{� �C��F ��,�i��b��;u��k��Bp�#l~�#��.����`������p��p�6����`'�o���i��Ѱ���s�ׅ0d�G�:�p|��4=�� �!�!���K�����!�0�R��j�I�U�S��&L���lI���X*|��-��9�'��<�c�'ؓ�]�8�5���:Js��/��J��L���n�uJמ�[����0�Y�S��STF�9!���se6�ʶ�;�]/�rRA�vZ�'9����7 :���b��'��5�/LU���8��|���A� ��
}��J�d��j��q;�9���pC����O⾴� ���pl�C�HFe��*/Km7���Z��rkΚ��nCcd���zW�ĵ'7Og��(�	6�Bר^����q��EC��4�V��\��Szb���>�C���f��iߔ�QQ��|�I�'8�w�S��P�M�e�	��Ӷ��1#΀�����6��]'�AL��p� ��ņr�[`
��(�W,Cѳ�
�k�����&kp����2(���kd��l��[�����n^�Iz�0\�2ܬ�����:����`ن]�pN�p���!��r���_�^�� �>Y���њ��l�����I�,�vZu�=#=_Ñ��@� z*v��Gg[�[_p������>��@[��z�u�R9�n>�9����-�4wg��29y��l+0�+]��JŒ���/5��(|�=�=B$g�ҩ��卆�.$��O�P��f�^;>�<l�{6@/�*}�?�S�:��4��L���\6#�<��œ/�Wá��z�rDf���)�p���-�i�lD��/�$9��2�m!b_�6������VF�c��|��r"��Q�ڦ�^�D6 o1���"ۗ	-޳�l
�o�n:kS3E`���Nfp˷�4��\�L�LƿIx2� y�����FK
]S���y>X�̡W�S��G�F7�{�g�6���P�`�2Id��榲hT�[b�7ɱ�����3#J0�fGaֿ�6ڶ�`0r�<�Y1��8>��!FmIRiF2����&��y"?� � �kv៹ٞ��(���Ov�7b2��T��J��,w���p<��K��,������J��pFk=�r�/f�ً��-A�&zDy��� x/`���n�mMYR �3Nu6�:{�:Bu��P��3�ų���
��i!nz>��+bN"�ZceY�7�~=L������ȹ���k�zv�!�IO�e'�A"J�L�����HO譠���ͼF��Qʜ�e�KMj��f���8:'�^K��,�V?����Zú��7Ɂ���r��g+�3�.�vJl��*v������!�C�������t�i~��y�Lר�N�ə�π�����j\��F�\2����8����=�,bBH>�cN������')�T����J5R�ʌ����J	6�O\o��Lm$3`�;VH�Pζ>�]�(w�?�H�$�`<���J�� Zw�3& ���@TD^�x�7Մ\��N��Ɓ�0��'��&�Q�H]N?�XM�J�6�_ՙ�q�c]FL�A�� 8m��^�؆��}�=9�%[Y>�����IW<%K��tӘ�
>�Ǩ�ȃ�Ù���f�Bj}�ַ��Gt�1��J�&�{�c�{Ԇh��Zj�4U��"�X��|��y�?>	��I��W���	�yX��X�Ӏ�Ele��)�Ȥ6�	V����� �X���uKj/Y�+���S�r�xj���ꁾ����xuj}��|W<}8���$�q+�j9M���`2E1t4�"��'�<��Fj���IA��B��51,`A���X[�������>��_�L�拧]k�~&d�����9�7�]NEsZ*i�K�ed�?ͺ����?���cW��׻��zy������SY T{�)Ԗ���;H^H��ϓ�x哫�ٚ�*E�#a��+��7[����b��bi�A��E�I�]�#�\�dv�j	�ܰx�!Y��@�chk��5��!��kNb�h?�1�����j�e���ù���J�*�|96}1�ʭACv��q���7�����?�0mdP����U�E\��a�%]ՒS_J��_?`�=w5�"MHҮ��W`��AD�=x�>���z�Sa6^��V��+I��3�[��NT���_�٭�"�}A[jn���ˎ�,�!�
u��PDǭ�ؔR{��|��������TZ�U�g��������d~0:�>���:t��OI�!E[����?�tl���WV�Na0(��WQ^�䜠�I�Jב��f?�}�����-��5�D�Q^"3Hrb�����j8g�Q�0A}$��1?�OXJԶ{��拖�"��+a.����pˡ|��Ry0~7�p6�Rzd���գ	�<�{OL)нn_�@ZC
�PH�x�l����y2�e��H~�d�o�FQ@����a���Um&I�����h	�
�1�3���'2f]Ws���	1vw(}b�♠ᅞ�d!Oڲ;˂�k��@��"��b;�$���Yv"��o[ /K�8ޣE�ޞ�Pu��U�ڃ��nΠ ^B��5��o�1:Ã��û��0c�/j�G
V�w��K����v�͂��Vُ�Nh�O���SX@���-W*I~�CS�׹lu͜�Gc�����>G���&�E�X�[l��ͻ��?b�y[Z�P�;@R��hu�?-Y���4�h��"/ۼ����j��ლ��$�np�iN��X�svR������_T� �@Lp����3kZ5�W���=73�͔߉��N���38�j�h�y�������4|)��N���Ր��w'�!C������50aU��@�U�l"�9���7�7������Ԥ}�5�_v⹦��~6�����Q���z��=��3u�I�B�S�R^u�Mj�P<{o5���tɏj���fkH���rh��I������]�-O~�kp���ˡǽ�a;�I*5�:����"�/�anBC�b�E�a��R����O���H���"]����(�J�O��輛}۷�>��W53�L��4ˆ�j��0V�Ц���Cƺ���+����*��kEk6���L�A{9^19�Q+������\�8!�%%�����Μ�n�� �5D�?�|d�͔\_�2#D����VWƲ������9f��g��$�ሞ��[ [R0�釰>��5J�,�'b���k���sAEwA2Y4��f�O����z�|���MG��Α�g"(�[���~�	����ؚ��[�Z=>A�& m���Z؅�_��-�bE���No�hg�AV��W�A���)ul5E���D�폼Î�M�-;�θgbI�<m�F���#b��Ӣ��h1�7��wX���ݙ��G�H�m������JZvBa=�e���i��f3e<���0�j�Է�����/�����ԭ����(\��k��8�9-�%{,k͑~U��q�9�c?�ͭ#��ճ4���v�M�v/�Y��z0$�`��`�r:�X��F0�Ն��p���И�Tk������&_�u���ܳ��1W1_�9�@��rG^ ��./����	�����}㆛{x2���x>)0��
�lN!�6ϋ���6�}�;Zi*I�&�"
�'{�U�7vlN�n���wE���)� `8�a�i�4gz�d�����FOY�#�S��0��Kg��kq�<���E���0wA��qJ�n�6:=w�>��O���ϙlW*�p��a�2����Q%~��`��F�!��(�����Ps������G�أl{��ZiU
��gM �:��H�|�f
��J/M�c��6�>M�}Xā��96�S�Z����^d���ux�&$Wb�4�|�H���A'�y�7�]+���`=P������K��C�9l�9ܶZ[5#u���h
ȿ_�A��ѱ��ih�*�_W��W|���7�ӡ���o�`���AH�o�'�����i0-XO���C#�����ҾP��B�Ęk�Ѿh���oY�9�ovT,�І)�8	g�|NryLc�����]�t��%MѩR��)nTwY������Bj#)d�}���
�XA[웂��y�*VyRDIOL�'!�ÏE��{4\��a��SЛ�v�@(��8	RIj'��BfZ'��� ��.�K�@���y	�K��۩�O34��������ݴ�Z��a �v�4���IfE�U�P�!W]��l�Fݍ����ZTW?��K_J�%$B�[$�'܎�$;�b�N�ڟ/�F�_+O����������dO�.NG��@�tu�&��x�0� �5G�kM���A�W�'�@/f�^DdyT�K�	Z��f��)ǉ�,v��1JۧŽ�cN�UM�?0���j��v����%(���#���`���E	�Ԗ쭋��t�;$0<��3�CH.1���~��(���)��6� �"R�/Z�˂��T�$t|�yFG,i�aҭ���'uN ��#'ǽ�����n�j�,+�����d��'Q�����+nc3��D`��ZQ#n���W��VJ��%L x��W�2A��+B0}	إ��>�l6�SFz��� Y�V���״%�@~P�\].���e�=Yq�W��Bgmw�����Z�8Ȟ@������h�P�-�e	Rv����׫���O�$�v8��J{1`��& w���,-^�? YLF�RJ���V��$eD�A�)9v򒥫3�R�����F��� �b��7C9�hD~��F����u�H
��]������!aU�ʧ�ֺ=���48�LXh�-i}��I�=B��]�&&�H���ቋҼh&��_�3�Ӓ|��F�I�W	99������Г�'
inl}��hD���T���C�o��5ml֡d4릉���RA1p\)M.\��B82�Q"�T��x��cPù��D�}���ޔ�D�r�_�k�F�%��|�8�J�}8��1��I��mj���G����9�b���.!�~`x|]i����sf�I6�ڍ���
I7̎��ֶĠu�k>z��d��A Y!h�<m��]&N��� �H|� ]U\6C�D��oM-��W>����ߎ����li�:f>oC'���K6|1���!+๚:�m���	Ԧ<�[���۸z����{��4�8�-�P+�0�QG�:�Xc��_I�wqo=���o*$�.f~���GLV��]�R�%P׎�)�`�����2[�6�^���іz}�Z1E���S!��,jd�΂"���S���3[vl��O�x���D_�|�ʽ�2qg�p��{�g����C3`ɚ�u�;
ۭݒ��1 2ҵ��mYc�+|8���6����#�R���ٳ�¶�HW07й��
����ֻ'o����uZ��ʜJ��)�-�ᆬ���O�6��ϗ��>,��p��xWr�ҕG\��4�a�Xj���'l+[���-c\��
1�������_�T&\q9 �y��r�^��yݼ���HײtF�j�0�ub��ENH�22�������M;d8���Jx�Pn+6���:v��!B�,�Q��\
|=d��N�F�X��)Q�o1�W/q�-T�ף[�Z��6b�y��j.R9��f�o$O��xݗ���ש�w����뇲�D��:;&��?��9���c�R�M`��l�����������(5���;����c�Fu��ȅa��9��ř+4�]�.}����9ܳ��y�G��K��7ޣp�'/; '��%6�G�WD^�k]!d�A!�6-��6��~f�����G7CP��')��#�����j�9-�0~1�_��gw�RI����[jۈ:�7�9f��ŏ+fQ�0}j���f������'�,�������+�{2mA
߄�i���������e���l96[�p��K?��B�\ �%�������h�`�#��I#�tf�F)nr6]:��Rk x��_�.�ǃ��{#��g5��"M��X�Q��$'�]My�e$���-p4��&����S���ԅ��)��!�`�d��6�0�8�R}��۳Yݪ�}XO��ö�O0�	�l%��u�|r���CeO�A�elŅ��yq�EX#�@��~�L|>C��X�XJ�����0��G	�Iҏ ]�,$*A�tC�&�u��&(ͬ9��P�e�+dЇ���Lu�(�S��P�ׂ�$5@g+R�z�KT-H��JW��ON�������/,�d��D7�>�YC������وS��J�k���J�7w�Ny�.���7K���3Bn	.��v�lu��>�>�D� ��>xe�:�~3��U�`��c��OD0a�Z�rF뎲)�&ܷ�{�z-l�0��Wӈ�	���Y��o
M+� �,�d35aM�'�d/��|QLBKދ��3p�l(�[>T�(u�Â9�nl�?Z�+�#U�erGx;v���n��b�ћ�-Cz���? .\�|]�ؒ�uk���o��Q�Q���╅��lڍ�,��̙�3+QBx�ؖ!�֜�D�qe�*@r.[H�H��H�G�O>e�,񸽁�VXE�c�N�I����f���x���}��5eY�)h�<)��eY�F'\p��wK�r��	�拾WW�u*b���l��,N]0��������Hp6�'L��`�E�"u�!���)��oK�a'��g(q���1��c��u{���Y�֞�� ژ�p�ڴNo�A1ro�s���+�����j��V���B�*{�:���)�S�RD�d�]b�k�z��$�v�)�\�\� q��� �a|+}ޡtY�.��:~��l��&�t��~'�aqH�y%�����b��p�/�@��T�'_��97~�>t�������2FG91��!$)������D.�o�;���9tZ��qp�?��a��TG4A5K�5���o�'�F\�l�,�-�
��Ş3��-���+��h�A�&�8�,Y�&���J���g{a��;�F��߿�.wk�z���}��Px��*:1#_G�����!�]���O�ViŹ9�v,D|�m�$y�sm�/Rba�ì�gNJ=Y���P�n��#�15���3���������Ä:�_�q�j O����6gݐ�_eLY�.Ǵ�x�"�{f�UhX���Ĺ�.�^��y0њ;�|��$���j���Q�r���#�=G���}S��µ�Hύ��&�6�S2漺 芚�dZ��R��6���U�`T4YCb�c9.����{��ϮV}�x�0M�z��8�w�K��D�;2���.�Yy"K4=��js��|�-��[��)3מTi��k���I�@7�hi�ڞ��
�a�/J��a��_�Y"y�t�g4b0pձF��k�lzn4���Ѽj�0�>a�z�Xp���Z]�i.) F�FI"󈀩����)�/�2@--u�D�@�������H[X_��R��[(i_�|&1�f�rހ�����u)���\�#d8���y{ː!P�/�H�4���g�h���ޛ�+���Juk�!����@�����^��v������:,�jv�Pd��󃔃-�_�a�4�z!�����<��2Jv����R!E�����`'�.���E�"�{��d9�i�ϩ�a�r���\^�t'���<�
����j���!Q�C�! �~x��m����鬘�Lh�0���=9~t�oA�1>���G��aU)����D4��cl��d�]HO<E]�RRJ�����/�^�M᰻h׸i�B��9R�puv٨�e;d�qv����dFeq�wr-�������U��S�g�Z6��n���p"��2кPN6�6HG?� @[>W�X� (������J��~ut6L��K%l���|�E�AGkv�rR��䴢2�OE<�o���.W-|�r��O�q���*�l����8�S�v}���H@�6M$��[��nD��V:sG��lZ�K�;#�d.�X�v���;6'֤���ע~�1�H�p�5�*5�m6�BY���iTx]@���٬��u��2����\��Q
m�A�7LL*�wK�d���#��S� �Q�I��m�ݘ�����Q�6O�"O�۾}k��%���4�PU_�<W��H~�-����#���F�f3}�7�Ġ�eV@�ϊ����UT�-h�0>�w,�ڎ��]�G$��m�wSį�U}F4�M�
�流Z��ܮ�Y���L�+�$d�vm�,��)A`���j�l��C��m���V,�SNOo�ȁ*�u���-�HP=�����+u��'Ƭ.%%H��4���Nؼ�^Q%�C��:1bè��)]o�!7��9 B��U�q�xP����:f�3q�Чe-�,	�HO�HL̫�� ��Sb꽱nr�~%��<�O�v��������:����gHB���L���I�mF�m��^!��ի:% G4����*��a�"�8+ߵ_*DL��}`JW�����ܹ7/�{]6�X�81^;��h=�v���g�jm��Y�f�E�	��=S�+��\,�C�� ��q�Ta�^��&�> N|^W�+ҎR��ح*=��L� �c�j��:My����c���#��õ�/GǫXї�8��<##q��['����,{����� \�Wh�@��Α۲�Iu��*U󖤦��og�!���,:�:"7�����Ӊ=�0���_�T�x`��SM�湲��t����i]�>0�~���\\&t�]��%�N�Mk�d?!HԳ�-p8<v�Γ����}Y���y3Y4Na��]��;��=�K��qn�����A-���G�rp����=IV�U�[�������ΆLy�
Z�iM���bC�+hT�MC+j4Sj��h�K��(��D��󭈊�(��.]�>�fy�R����؄u�iIɴ����|Q�]���Z.zqV|0 �Z:@�ܢ��A��b�؜ݒ�� �N8j��6�����.�~<7�ZX�Ĝ����4������oxn�K���(3����±r��C�e?�ө�k���l����)�UI(��B�|ŉ��J41�eB��x��IE\�rh�i�c�M|KV��ߩ��j<�za��`!1��봞ӫ�"�gp�()�~֓��N��&�7ſzkL'�3Lg���'�A�$�=�Y;��c�ן�G���{�1�����|ms��XB�i�e�M@C?^���-����$�����7��V��,q�<���k��
�"��y?��ٽ02U��:��zI�����:����4U]Se�B�Ҫͨ��0���d�
ߖ�M8�U;����"�.�[=�b �����v=R=t\�װ.�0Q��-�r�P�Zdr��w��^a��2A���S�)����wf�R�{�&��O�8���'���+`͹�3!S��䇛%4rx���og�D�l�X����g@���9#��YRF�������Z�IH���U��A���(�܏����Ջ"�-�wp�DB]���W�Ӭ������o�{u�����:��R7�l���JŪ�ﶞm���f��5�g�HB Kz8��W2k�855_r��},n�QN��>d=Q�w�?�[�({�ڂ[hu�m\nO��2�Ŝw������&MG'F�����݃W3�������Ð��5Me�`��R*M����5��R_]�/�lU{d>���pbr*��t�\��Ξ5y���EmK��� ��\6�ҙ���2�f���m%HzA�rm
n٤'�w�,�U��:�j��o"u�[��Qs�N=A�<�P�a?���k�L�t�Ϛ/8�K����h���B�l���u'���ꭾ�x)ķ�_�K�~�%���k���p�����)�Ȟ�����z+6�I
�J������b�E�`�h��$�V�����x��f���+�vzSP�['��e���E
QL|n!�w�V�59uM@��M�/��u_m,����mG���х�F�	8��fnH:�Y�H��.Z���q�.za��I�'1n�q[t�c�b����oJ�=�Qc7jCZ�(L&�k�M��^�����)��r�����$<:���b>�4\< x)�'�>ޗ��^A&���I�d�������fv���rx�"�KL��8ޣ�s!��Ƶ����K�k��Ce-C��ʵ���?����r�$��UNq>`8 ���8�t\�P��ߛ��ȢҮ�'
�� .�4���}2��'�=_�!���qki1�%��[k�_�2ț�P���L�C)1lw�%4ӻ� �����'=H�.z�4|��̹�VqL7u�A�j�7\B9qm�FT�`y�����<�@�Cs?�ϛ�qa?*��F`�e��W'㊧�D��̄�����{�B���5!1j���+��ۣT���^_�"��?Z�ޗa]o�,3�����U��ᮜ�*H�k`��)�+���7&�eU��1�7Ϯ(C{D�C4�2Un������ȧ�@/>�����v�t�\\�g�aJo���f�#O{	8�}T�/������HI��/�@�6Z��Z壱.�c@��^	]��C�2bn���02T@G�;��,6��l��M�����,����O#`y 2�= ��vE���*&s�d�1�ҿ�K8� �D�p�~���ύ��3c�|��L
~��4�N>�.�ylK�xw� ��	鉪�("RLc������}V���Y.��1�՘�}���7p����Rm��ה*o]�hr��K�:�+f۾"L9�ӗ�R�o<9�h,�|�����5f���oOĠ�-2��%��Gh����F�ڀ�О!��R��$���ȋ�J�ľX��/���������sV�����*���bPiI��O��EQ �MdV�~ -���"0ڶuR1�ģ[dܮ�Z�;Z�T�s�}��"��#-v��^�<�{�B�׵�x��.�q�Hpd��\���t��'H|�E�n�6}�̎�_-���'�0c�dT���n4�8u_J�R��1O�wنk�6�)�Պ��?��	��m���kO���?Wdp��Z���Ϡ���ђ��73_4۔�AY����-�X�IHv�*�Z��
���>ه�it��R;�\ԮO��AJE�zĀ�T�������65_zE��z�@���t����,�W�v�|g.2/��ew�fJW{�߄N���\�C�Gv�|� :�l'��<'
 ����ȧ���e/�W�BӸ��n�VSwtF�!�E�[�<w���?��/#U^����G��ҝSEi�������i�<��=<�,M_�[������@�p��D����v>�wo�F�s{׋��͔F;�R�&���%r�à��e����d��P��͔Z�ToQ�"��l@���}[�~�n��]��63C�H�{L��@�KK��`�	����Z]�I�����p��78�'ٹ�T�n�벶�%��x,�פ�Ͳ�le�;�$%
j�����2-�iD76;їTWM�F%�*�w`9|h,B�ic��qX�D8�đ�m�~�-2�m���1��}����6�d֚�����B���k��"{ NP�)�M.����X�ʺf:��<�ü�Igӵ��Zk��Nt�#��H\��h;�^5)�g'��_Q��� ���إ�x�g����Œ��^�����Nw���V#xH���O��˗.6�QB����P�T#5����mH�͌����p4�O4P��TZR44�&���tA6���zRB*Cn�W���3�:W��O
M#7�;���Y�;�e��M<( ��2�N�j�#%�`?�vHY(гX�$]X(o�� #���v��Sftp"��<�?��0f��9^�~~�O{���v�(�a�&�W1qZ�҆�	�~��í��B6��n�����h�h$9�˞���9ß�V�d�t�����OK~ː���m���PR�)�Nѹ��D��sIN�|S�),`�O�=b+n�С!}�L�74��L�����ֆ8���Ǽ�� L_�@�	,��%ZU�Pt�?�f��f��-��$��;W�ZE�j�ҷ�-�{����2֒1�3�len��d�X^�d�_
�;в��<����<�P.�mh�>g�e��g�J$P6!�lWJ�?���v�̇��9��5�ڟ����x��P�Ў�)��Q���������f����;�R���k��{�a��C!}��@����Z��_5@6�hz�W)�E΍U�o��P�U����)y��U�K$� %�No"&���A��2��6�ˌ�2��C Oj�ǆ�nF��y���tr��J-;�|����V�9��1 g4V��U�á���<01K�߮�i�t��͌)��4�bŎ5��f����bAu��%���T<�l��q�O ���đ�i��ܔ�J#0�����E��V��Q�~���b�6�A)+��#��J�FKޟ�-�t�`��!4�b�����e�A���fҹ���c���a:�V�A4�5;�k�q�W4�-+����~]�`P ;n���Q�a�$�Y�g��9����� ���e����.�h���J�cm?g �Y�Q;�H��m���M𮙛&
����آ��-�'#���^u���ěٕ��Y�Ϣ�
���<U#��,����-� fE��/+g@!�������Bŭl�O|�38i7��U�!�p!�	�������{*�Ef��'�r����p}�s��N��3-�/�z�����|"��Һ��MMA��PY3?��f��CU�f���#�J���h�Z�?�̜>P�XA���MlX�����^��$��g�5x���X����.��o8~[ԃ&P[�e�%V����j�U�$y#����B��k�Dk�R����&_U}����iK���=D���L���Τ˗k�;�������BDK�ۋ̻��n�$��<:
V�oH�Ⴐ��T�99<�>Q+	�#��r�:����iY�	v#<��7��5}���('�!���ᓲ��Ȥ���M�s���.��T7�mh|���_��]o�xr�t���O�P�A� ��U/Gݻ{�0	ڛ�\!^"j��
 A?w
�[9�QmQ���-�e"��;$=��=�>�˖�-��FR�`�����׻Шh�J'����"���J��i,~)MP*K�� ���2J�l���\� �՛�{��{����.�ұ�����%�������V�2	P�e�Dy���~W��SwK��}b���v-ا��k)[>0�1�s%Fy��𿯼��G�#p�i����Y����[ �ܹ�U�LA�9G"f�a�9��U/���RPU�R[�-�n���&sG΍S,B�'n{ƌ�ͿW�͏5�.��`�����������#�v�5����-�FQ���0�@��<�k�L3`�<E�y�o�ƙ$ǁ�_I��v�E��u�lk�,����eA�!ԡO�F4^���V� &�>���1�>�� ۦɞכt���̢1z�z�ް�����tc���N	���Fz_͙>̂�9���o����~��6��C��T�l.��X���6��W�:.0�a�	��8d�h��7�ul�,݃L��G�`�#��gޏ���d�ii���\���۰�-P-:�l����7��ҳ:K�ǝ1ppe����S���`FG*�Dz=��^Q���̯[�N-ћn$���ss�i�X�6O&q�n�O��P�ѐ����J���T��,@XT�Z�T�c�