��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ���������-���8��o1�+&qy���1��=�%bا����%IҬ��Xh�.O�۾���0�]I�yeIR���k���K6��	T�����z��#�?�)�Ka����Y0Z�r1����U̻yF�ՄД������s�z�#1�FS��H��s_�S�*��;��^�>Y{+����� �t؝&���M���i�b�N�!��`�ջ���W���s<�غ	�xy4�I��Fa-�p���DJ��J�5�鄜�;�S3�R:��5;!�Bu���"�]�0��1p-=��:��Y��rf�����?�n�T�6����9��7�l���6w6`i_�8!�at+0�G��f&;N��!�����HRsl�>�5��Jm=�
����O��?YJ���uU�	�}D
��x�����gK���+o��ͣ�L���<�	��x�Ok�3"�D����^/^YR헁����k������	Wp����2�#�߬_K2>. �]�\�䛌��7�O3h�-֌�W�.� yX�ő&�~>���Rz��Ԡܮ�Vش���}��h٫+�x{��qŮQ�+�c&�`�8{��Z�lH��q� �F$QN�5��<��䇐Wa�U���$�F�M�<�F+ɸL�X�ߟ�(n660 �%�1y���?��P���� ̷��/b�vQ��(wv|����c�_�2Q#�%�eO8T)����3(�<��B5D����D!3Kd:|]Ct+�u�2NG�1�,���	����`�}G×�'���O���7���s�=نC?ii�F4�s-%1��9r���=�mHĦ�u��lю7��vؓw�s'y����t�Ւ�J�C F|o����8,%&����Չ��K�%���|b�'��'��~�f5g �P�@酳����ӆ��AVG�݊ԧ@����ˏ�{�35@xi5��`IY/�S�iB�G�;=�"�H$�����)��Ŧ���?�j���ŕ!P�Q�@�o���q�� 
yě,��7匬�8bG,+�2�������@���%��>���C� 8�ڀ3�����=�=!I�([���-u�K�Zz����T��g	����,N�Je��ï]�����/�_���B����������=�L�r`����ʘh=���;6ݖd�7��.��\�55�#Y��M��sUM@O6_�Pe��v�p� �ey˷q��+��ˎ7-z/3Ԡvm�����Of~�w�Y��v� �{���@�ڿy�z��M4�>�!cA�٦q5�S�"�Ǣ�H���9��e�r�@���������ād^`�6s�;[o��~���/Ѿx��x�˖K$Wg�wE��\y"�XVĿcY>�1if�ȑ����Nx)�E�Ts��_�6��t��4��!���>��m�e֡=�s����Wx�t�g�Y!4�y�+���9k�_��,7��(��Ԏ����`=�����̃Y�,���PW?�q"����X��̋�t�'/	LD$I�=��>�\Jh��?	Ꞅ0&��3 �Lٳl��))����ֹ;0��8=~�hF��V�%�������)
�p@�B��)MHU�ae����ap�J>���H�cC�8��������5���v0b�1���V��L7�8t�4TZM�4�,/�'��<"w����O��P?�����"��v}���qQ^��O�W�j��q�z87�\.//�S̮�9
a 
`"䭎�\iNGd�˷ռ�S�-��������U�ƪ
��+V�Ϫ9x��M�FG~vi�/%�"b
*�&�vQ��g�_&���q���#X4Y�� ���N��Ln��܍�P���~+�T;E7C�
���ӤK�L�g��(D����Ԇ�ؘ���q\cỢ�����uRg��(���w�_Z_���0�K�q�>��6�W:g�l�j�"َ��ތ�j�g�N-����`$'�m��:I�^R�-j��L��x�J�`NG����z����*r�v������ГX������>5�S�eҷ�ś��;�=�t� L,��m�\<�2��,�޾yr���y��zA���hM7����X���D�4�3��X�m�|���m�gPpf欞�+=�	����0�)()JM�n(��&bW�7b���rCL�9(���p#�y�W�T���<�c�z���/�|e/��\��o;+X��m��ͼ�ի�\S�Y�Q����@�,�&�2η�x�`"I�$��:��h$ƪP@�z)al�V7,盔ֱ�hE�:�E\x��l��X�����}�q1�[b��)D��.)Nn��Tx�H����%A	wЪJ@K6*��XO?��_��v��U@��	=@)+:����s>�:}Ǟk��j�,k����"=Ι��͸?�&�Q�yU,w��E7��hX�.�u�/�PZ�vl��H-��1Df��Q������-�3���R�N"� ������l@Д �x ��9W2T����Phr�ڕ6�0��Cf��I��m)�FLa�^L�-�je�E�tǎM�V�4�h�.U�?�V�T5�H*@m>٘�D6���/��I_e�K����d��C0I�Tec�t��z��ً��F{��IߦR���ڑ�]?�f��7���[�uv䝚�L��#���B����K!+8;�4��{v��O�nx�dC�8[4�MUY�W�ndT@Q��ZlV���BC�͔�;�=ҋ��r��8����$�:�X�W`�"L���7{��8�_�KBF��@��X������d������fD{L��I����l��"�F}��ѿ�,�	v7*|I���7c�p{:X�=�f�3s!���u3Ւ.����i��,�����^��bڼe[��<Z�m�Az"I��#�����bۂ`�Ĺ�4��9���Ă@U�6�\��o��=�\D�������e7��Ҿ�V&����)ў�ͶN#b�H@�{�1�	Z�ˢ�k�@TUK�DjK�����)�ۺm{OU+�ُ[d�.�7L��v�Nŭ{���M,�:a��g`x�a�% `.�|�[Š�_�|i�{�f��y�rV�#?�,���βAqik���Y�
�?L����% en�|ݳЗX�e�b���Jn��j&4�P�v�rPk	a�{��h������q��z��/׊���?�\m��p��;�^n��>c;'4��b�@ƅ�Pt	�>%�o�B��p�S���aCZ���\B}L_E��C0#�w{�C��/����\���ƽ����o�"rj��߯�s��Zq 4m<�hŃ���$� !8"U�����Z�?�u�$�-s2t���M�^	����F�3���uD�P����;_�}�2�E3A�8Q3�&�JD�:%g���?���eT2w+��+m�^���Ӄ�A��	2PA���f]z�xa��V�9�W���<��x��������[�PIetF���pj�A�7���y59��U 蛥�W��:Ҡ���u{��;e��!*L���(׉�p�q�c�.{8�u�^^�"$�C�i�j�c�
�� �&�@�����Q�<��:O����` ��ob��B��Î��:X�h�������a�S�̻��F%���´�}��ӂl���w�ˈJ��hy:6瀤Ed���Ť\m��/0�q�B-wVcۢ�굫�Л��M2z#��:DNK6��R�I���'�dd��1�SN�&k�w������ui$��
�<܏N6�k�����.�c����:8�Q]ǚ1�����>�z���#�'P����Re��SܥƵ���킠%�,7��%HT�m�&h���pZ�h��W@�"-/5����f}3H<�i4Y�,J��aJ��������i�b$H���,7-��$c�]� B��lr�]�l�7��������8$f��v�_�"vPE ^^!���1hk�+��Nf�&�o��A��X�r6����;̷%�*�wƽ+�CEe�:{�¯v@���/�`�VR��a�Z֊=L��D����-t3
�n~��ǂjrop+w�R0 ����k����P���;��ˍ�������s��_�rd�"�k-Sm���7����A�����v�;L��kZ�/��4��PeOTek����p�{ ��M�h�4�l�8���6U�:/;S�����GEf�Z�g���ȽI_ �^��p�f�/���-�;V�/��`�R]����w�~���O�)��8j�^N�6�k�)�柡�]g � qǆM�4+O[$�QY���.b����@��0u1d��� ����5��;>�e[;��-�o��a�	V�d�cUP��4���/�F^y����I6)��u��Ekw���x�
e�Vo��Wg��vm���U��?��m��D�݂�풥��A�駉���=�&��|��7�o��bˀ��xC���}���A�2^H0���c��Q�ZE݈�u��к�E���sʓ�����v���b���:�h��^C; �]X=�C��$�@��f�&���(�-�GkW#R-���}�]s��N>_g�Iy�-~� c��i\2|6������'*���� �R}Q��ch��fe��\5���]�D�7�@|�!�v�+���r�� PGۗ�w�{��B��I���N`ϡ��f�;��3K#�**�F�� ���j�� �_�����	Zx�D\�Pr�P"�&���j<�m ��������/̉V��d����7[�vt�(w�JB�գ�]�x��c� 0	b�m���3�b�[*?gZ���_5�$^������������CL՛F�~��'EJ��ʙ�P	��P�Cc��� ~y���3M]T�Lx�c(z"�[*@p��H_}�*g�<H���8�l�o} ����V#Kb̈́<g�G�b�&�HP���vyX�����+����\W�u&�V5B�a�D���`���A��	�}5�����sGƹ�[&Waw:I�p��}��#���2�1A	�~C$��2a.����b*�n]�'��7�\d�)�r&�����\�9�N���4ݐ�XH>�S��}s�O�H/އ�a�nۖ�}��+�?rZjK�>�Y~������~M
ԑ�0@�{?�m�%4���>a����^!w{��Ԝ�����#�pj��k$��R�R�eX���.1k*}���ea(���ą����.�\uQ��j�q>�J��8��i�\��I�U&q���|o��O�"�5d��Dy@=a�l��d���֔�'����0�"��GU��s8�����%;6�ZH&F\���h�-�FH�k�ܯ���'���ئ\K ����&>�8����\���JG�Q[�w�*X=RX|�0�������;�Ieya4�3����{g��b���g��V ����a�V��_ाץ��4�iG|��>��,H��lp����\�xWK;��/_��i

z��Q)�Q��H4/�˄p�R��5!>'�x�[�Z��_l�
��,K�=1�N������bk��u��-j�Ȩ��%��%3A!��8m*�w�\&�	W��`�wX�(��o��t��oJc:H���>&}�a��2M��l���[�GC�A.��O/J�FI����/I�����.Y?1kC;?�倁@��ў��s������d.�i�3�g�g�2���ڷ��I����*K��� ��d沚/�X�|�?G����>+�EƶD�K�{�� �(�0Z��@��p��|�BF�J�9�y%�竁��+��"��]ψ?k���6�-w���O4��Uu��O�1��g�Z	�1��%F��tv]Q����)�t�^���8��n\V��Ü#�lZ��"�ȗ"�T�_��{�nF���{��\0<C�'U#�tC�O��]�s#Z�;��1~-V�t"?�AA�6Um�I���5P��m-�&�j$���֋����rD�*�v����Q)��͡�Ճ(i�K��N�Ng4*������m�������N2b�I��:T�1�A�+o�MА�LN���LQ���cгF����ߢ~L���ݳ�@Դ��ú�6:���6�y$�wSu(��.5F���	���
�J̌��_���r��º�n�ך��9�<�E^s�2զ/3�e&�,���)��*
���fG��y,��5N/5%T{���ߥ^HcN����e��wGO\��zb̜w��;2�(0tUfN�?��W����-�<�˖Q)s��!�T�&�4�D
F�'בּqM�.=�qz�����_����곮��wY##�ף9��E��Em��fW	�fΟ�x����4T��$�XC�X@
�~%�?_O�g���#<~�(��b����jpq-�F�r�CWu�JQf�<��4��6S�u���,�A���r�����"G:ϭ"�p��'G{��d���c��	���N[$�#Ĝ��}U��	�2�]�4)�FT/�N����ͣTPQ)u`�A�S:#��I�P�7�E��W��+�R���Q=�P6X}�l$����F���UD(���*�'�Q�������6.�?���fN�?$J�)(�ê)1���\����Z<�7�'t65:��`�>�L��/�l�:�vq�D�WLe�g�$3F��e�߄ �h51�PrI���5����k���Ed�E#�Rz4T��%�]:�1yё�g=C"}����ن>u����0b��ߣm�_�E5b���_G�K��� ��z`AB(�͋�8 �3j�y��㖑kB��<�*i�M��]\��Z[�e�.�i-�S����V�g�"\�dL�4��3�������	7%�.�߀��o=��(�K���P�x�xG1Ԙ��|c�����Pt�@㸭֘����+���9��K�wК������B0�,:r���VCLU�d`ܜ�L6�xsS$�ӏ�[{�Qˡl����~0*Hv�`ղ�����}O��\�ՊS��@b�ߔ	� ���O���"��j�������HV�����؄���Q�#����l��%ݫ����'ѳ��aK�kH��q�3�y���g��zc�谪]���K�֔C�l��,ܐ�p,T@u��gFC�dMZ��f�����@�h�#���?��-��qf��:NJHƵ[��@Fc{���m�}i��)ŕo( ��+�Q��z�w�߯��ALQ�t\��G-�x�'�.[���[N��XI�{�u���}kέ�(|���W֥���E���0�ʫ�ʤ�a�&�S�8ӣ'���;��L�����^�ÜFR�G���*��9Gɍ��K�3�+A��1�=)|��:An�Ŝ<p������e�"츧H?w��xq\�	������[����'�G�pP3���V"-�D�j]T ���3�U�2(���J�����зנxY�&Ѹ�$�b�lƘdR6���pI��k�1j�� �s��I�Ú'�����A\=�ph~?�Y�����45O�ݽ8kֶ2NF���E�g36��ݽD�@2�{ѤW�	/����.�%s?�4��jR�c�GY^��?�al���V+�,��j�\�U����w���ʈ}>�Y����Iv�8�{�,�igf��p~9���oSԑt���>1�AR ��+R�Bn��ч��)�qG�*	�����E>�̌����������C���V�G%��d%uS���p��N,�)!�ܻ�Ɉ�zq�+�(�N����W9�_�w�{����.�Y���a������lc�r��u�U���B~OŅs[?N�������Ry�?[F�E&쏋��?#�Ԩ���eM���LnD\���[��5d����4��3�w������L�N4���0�9x�&F�&��zSU0SE�Y@tɴP�50+N��=C�7�'ߙ5���&�S�<�t 	�"-�	��?)GK-XkS�JCb�����J;c7��_ԉ��v*���C��E0l�I�4�25q�$W������.�M��G���7�N!��>��c38�N�t����dfE�v��o�zH���Ѓh,nA:�����@bp%�z� �S��$�sw���z�V��Z*�d8��¶N;CXd[zL�u�Tl�2U��.�Ve}6� !��nL_���:�*�)��0�%d����dṆ�5��t�࿃��ГG	M���5�-��Vdn �U8��6���V�
�Bf�q��|]6�
���.� �d�d
��Y�}�>�̄��-��"$9y�2�ic6^�^�ȋK�	+D�e���K���Irq�4��ԥ6�F<����t���0���{SGg���P0ȧ����U2���xZg�B���h�Q	��9�/�03���gBɫ�ј��RFb���`%�{9~Q���^ R���h|)�Q��g{N͙��;ܖ��_`�U}x��H��l~�-ʹ�D
��qڪ�����"��a�RN�w����|�-���! &QZV`�����C�X��"]��K�� TD�q�la@�7;�LE���i��Ǫy�F���2�Y]� �̘�4BF�j�1~r3	�y� ��)�⏗��������KLkZOz�`��XȄ�Rդg
	�Vu[�^��X	��*�]	s�БO.{��-���I׷�8�|��6T�f>ߏR� ��8�؅�M�����R�x��F����0]�j���L��q��W:���UВ��؄��2���b䄶�|�W�/�rg�4����Gc��o�7z�X笔N�.2�/ ��6�<��2C�%d���N��n�i�T�f�d,�=j�un��=��R�x�a	G��|���8/�;�w��>p�z�~�X��^�'���J�Z��p(tV���F�cp4l8�[WS��X�c9�	�j�<q;+n)'XYaU�c�~���^{�Ŕ���gY`%
�|�y�4W7��5���������V��!h�k