��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ���������y@f�~?A�;���\+P
Q��c���.S���𓴡$I��$�+it٩���.��B���jԁ�=���MMk�P���x��D�\����ڒ�`�p�P�����[�J����şL��6a��y\��2�ޏl�4�&�;�m�N"���d����<����D�EջZ����
,��fv1����ꁮy�Ζ���A�^r4�m8	��S<iDf�5�u��.�PC'|���Xt�6�.Ah��sO��0N^l�m��F}�ﮇ����_N�ɿ��@g���_��x��CE��t�!��y@����X&�jм#B��C� �ۋ1��1 ��X�^���`hk���@����|G�.��K*]3�(z�h[�'~Ru��J��d"�3c>
� cdy��@�Կ.Tbg�(X�I$u�A(������â9	=����~~�Q�4�sL��9�ˤ�QXFU�w��h�٠���;� �F�LԷJ���l���>��8Y�,������}lE����y�Y؍̗pݩ�C�4�&䗜!�Mt���K�[��6n���g�;q�R����T�C�7�e����5t&!���fl 9�a	JJ47�̶������2^t��S"g�nSnCh�TdX����8���=u�p���d��&��u�����b��4*��?u[5�y�.{D9��y�:g��EkۍJ��7LX-F�^y���̹K�o����A�6��_rH�٤�ŶØ�%R;z���b���� \W��N�t�*2��C��W�ܖ��%Y���U���i_3�Le�w�r�I^�$�L��I�?Z8���ᤙ������/�	XA�����Z�Lb��:0��ƌ]VH,QxWM|<'��ݏ�~�������e�ԥѬ��_3d1�<a5����K�Ok�x�'D>l��c �%�1�X�%p�����߬�/FrqD�R��{V1QQE0�Z�9��L�l}VU�K�U�|udJiPO6�G�|S0��2��Y'@����ߒJaM�r4 딓�8כ9�.�0/�m���ʫ�@��a���#�~�^K@v�,��W_4�����Y$*����l�[>���u�ƚO"D���x�̡o�q�[웇�H
,���9Sd8�gf m�Z�4�<{�OA4�;����j-c����f�
���.h1>^�/�4�ɜh�ͮ2��ώ��5:8v�Ϡ�U�I��?�@�$޿)�B�ҶO�@�����_`�ʶC
�^u�Č8��o��19��ұPF�LsƗ ?�맰#Y"K�
��Vu*���hkI*��K��H����ٮ\t�,�.�ҹ6��F!>��m�G���BMr��j���%�ް�-�y"�������a�Mx�>�%��瞰�eB�[.T��˽F?e�\�x��3�A������/ny��|�k���g�#�9��s,�����܀�m&4�^�e�����ߙ�%���"��9�����t>�W�Ym d��f���6x
�kۈKZ_@QRd�Vh�<!\`d����`16ӎ(e~R���t�a�u�ȋ� 	o���}������{F>{f`78T��u=����-��\�� ,b�,��xZ��g|:�;p��&[�V�ۖj���챖u���N�OL�|��G���7H 	"ߩ��>;z��-�nRe�<�����:����ilJ�v�n��3����ʏNw��|�6h��ߨZ���#Bx�Ņ!���A"��?0�g�����r_^�
ɉ-���G���A����v�n�9t�L��C��5խS0�笋36�89�����f�p4>�G �9�V�,�E?y���gg�o�#z�����E�`����?l��l�X���[�����+��I1���)�w\r_[*5[�Q�x1�{�}���x9+ ;GS0�+U�T�=:�ȤV(�|�Ns��t�`�s�R����R�2�d�Cͦ6�J���F�����%�<iY��&�[�����v&��`\�@���M�,������yO��>��H�Ƈ�z�=������8M(c��`Gպ�AgU#�,���%�{�ʳ* J�����n��33~M���f$��� X��Ԑ�h���ޫ6o�8�u�k�pǓ�+���F�$sOnX\��+��П})��+�zr��޶@V�� Y��3nVO;�p�'30�Ӷ��[?��Qa�y.������ǼAo�؁����<�ꮨ���LyJ'E1>������)w�����Z۝^������I	�.	[����V��'��en] �XR��O���������o�9^f��L"�&E�Y���e2��6-D�nI�0��L0v�����2 $S9fQ-���q���9��u�tjh�����A�5L!���X�+��LMldI��k��|A�e>�
��X�t��|��IV�7s��(&�����HZ-�&蹝d��ym�����PM.�đ�`D2��ġ�Vʁ^�A>w�P�fO��A����r�hn����O�<���X*���FOzgH�И�
̖�Ns�O���|?:�3{"ULܵ��-"����"K�̃ʾ�o%�4&]���Yh�j!�8ׅ���^�V4�'X����G��]�k���R��z�9<���8��N����RiZ��-t�	m�����&�qO���h`��Q2s�=��4�3�G��� \p�H���w�E����-\E>	7�D��� �	�8D*	��׎j����Vl2/�u4\���ŝ^c�D~�=8C�E&f��L(��o�Y���u�f���O9���g����W*�CA��k�N�g�;L��;-ߨv���@�rw�%?[KG4���0!x$�Y ����!)�~��f�T�!	�[`���`�R���ڦ˾�=&;���꛶&�F�����R0��-з{f�#�9U�C�a��j�@
5�hk���F�3�� ��۝I�0f@3=��d捅 ������Q����gS�Ԟ�X�d)�^�z>���P��o�dr>M�ע�;8�Z���m���+#���'��~s3�
 �>���_�;q���1��M;d���I���s�X���#��<�;��g�����ᠭ�_�u���9����*u}8���(�l��.i���B)Gp|�Q���}��Nuc�{9-Ͽ��m�+)���6 Ȳ}[�1`�4�[}�F�D��LY%ץ��8XL�+!�8��@S�R�v��4E�͹�p�--��|0�*��C���5���8!���~�W���!nT=��w�.�شB2n~�����?���V����}u��ٛ8���kG�����۴�2"��H����3��=^�ZI���**g�	�=�4�_b;=�yT����{�{�����f�:�����l�$�6ӭ�i_"_�H��[O��0K�8��:Oh�����f�:���:Y)յ�RG�?,�f���0������B;>c	3᫨p�Wޙ>�G�O�T
`i~E�6wS�ľb�*t@a��\p��;U�p�"�TlM�Rt��D�$),�ɘ�j�Nr@��Щ�}sfi6b�d7�'�_	�o��^������s4�H�im�xZ0Э���e�� ���j�I�X0' yjr}{{�����%O��g�m�q�2oT[����h,O��¿R���C��w��Q�;(]ђ �.���!�Kx���q�e��
{��x�6	��ϱM��h% Z_�ݺ��C�ͣd��u��C���;�R��>!�QC�pIr7����T����1�C��AN3k{����0}����^����сH���#n	S���˙�$#K���g�4���o�L�D߯).�U�I|�Y�[މ�d�� �+^I�Tp������V�%5�.����xt�7wˎ�ia�B=���d͆��"|����t��rٮ�(��)m�Ȯz��Ph�P���k�K���Ѧb�~�6�=�[?�
T�qi������`�nT�_�iu���<�$�^a�\݅m'�F{Q�f#:�U�<�Ū��9M޽�sDʙ�`�_ә Kc��v����CQ:����rBd ��=��;@� ���A�׆�FG��U�e�j��=��^����7�92�o�7�[�������T�+�a�`k�`"B�F��𸫤"�\�D�I_���l����-1h��#!h���r���{J5��D?o�7(G�*�խ��y�۠=y��t�,n��� 2��^/��O���1;s΄�(f��+�Pr�
�h��mspӲ)���#T�Bt��[���՗y%���A�8�cv�!9��U���`��[:x��e ,���e��R���ƪ�`�{��r�,!,-��6a��?�:���n�\���em���E?A>X?el���ſ���ǟ����ViE8(�R�^,�X��6��c� �A �� ������'����	 n?×��r�~�f:��=������X��yGX�2����{��7�n6�_ȇg+�!^ޟBC�lہ1�=rC�e��y݂�`� ��W,��(�L�F��W��%'X�T&ɤ�����T�"��^�`'0�R���+  �O-�q~e`TӳT�_Z�r���_��zH� s�)��Ձ�UA�����8�3x�f�;�{�fk�jW��	�#�S^{���/N7|��q��DBs����	���m�N���Z8.��s�l��З8�*8K471�C�?�3w�ψ���W�%�(qK�Cslx������#"��Ο���F.t5�'T<J�B�z���fW�qT��u�0��$�f��OBS�u�$9�fg�?Е��Y���殉�� B�0<"�f+/�;�y�V��1��gfC���	�}��~���!��S�G%͜l��'U*#)�q�p�i�I���Ψ�?�*��&]�ǟqv鐝R��@د�Q �x��
u��0�8&��8�Go7�[�P�su)�x��5�u�7��a�੤B3�G��c�'Ԑ/s�$s��y#Hl���V���WD�ϵ�7����57�@����ܘ ���.Z{��k�@Xr����{oQ�����/K2� Ȏ�mx�Q���E��95�����J�S�!i�/�]E���G�e.(K�A���M5y�	��0a?G��:J@l���d�X� �^O}`���<�B�2S��F5�۲l��!d��B�K��!b�s$�Y3��8A*�i�څ�Q���Ͼ��gUh��,�W,N�(���T; �[ː�����[bK�w�D҉c�/��}�d
��(��o��-N<g �f@��h��y�Gp������#B���칋E	n��@����ϋ� ���l��c�f���z֍v��|/�ݕ)B�yTU�|�I�HA}EQ�T����u�`�_�&����2�.:ٕ��*w'P(�C:�}�9IQ=�.e�+WC�kP�4�/���聦*�몚�^m~�q~/y�5 Q2�n��>�\w@m���CLj4�LI&���e6��kyU��5�ϔ�:ϸv�k�k#>��&?��c��u��wv;ӡ�$]��#�	q�j4r�~�U�(�X�(Ɨ���PE�$��s	O}�����Q��n�^�܈K7��0uG����/�*JK}.m�Q��ͪ��K�^������{0�R̃U��A����0m�J'_N�}\�'�LTT]o�>�n[�g����]H:���$��ᝎ(P?R���,N.j;`���+���U�� ��E�.A���{?H��;|�h�AX4������A������ڊ��$ �&\θ"��s��۳��~�o�f���M� �ܥ�p�7��L��N��ܷ���j�:����*&��{����P�X�
q�l���Z��Z�\js�D�T����p|����$�v���QP�3ZhN�y��� ����/��v2k}���ź����7T��Ϛ&c�(o�s�S@��qҪ�$o�$���\�orOd����ɥm��o�t�Q�dȅ)$����OS�;��"�J<nR|Ƹ�גvgs
R	=CX��^�UQz:�Vߗ��n�x�_�s4 ~����+:�~6#Vi��l,�m��M:�J7|	��H|�[}:'h�D��w��HU�9Bu?@���v��O6�������Ɠ� ���V Qz\>���f�)s��+��pnD�_L�6�L-�+��x���a��Mqd�wc���-*��1�<��`8XZ��+�ѹ������l`� m.��p�W6.�2Au�w���yhps�.
&�R�q��q�1�[�1�[c�ȵ��B�/t���H�a�M�QT���X�a����m���c9���������?�9�l�W����1b�F�B��D�E;�E�.a�a�fe.AD�*@Z./p�O^�ï�OU��h�u���dI��:HIHF�j7 1ǲo�����<]�-D����=Pg7���2�䟹�T��dh`t�ҩ1�S��(e�蜡N�rs<W�e;lqA��P��vj��W�أi(�@�#~�?��C���{���i���U�:�3r�����؛�\2���va8���D;�~s���W�hz�((��W��JF�e��yq���C�?���(P�����.1s ��k柊9A����
s�e��F���:�����ONp;ԁ)�j����D�(��lꜩ�iLN\��j!�*21�qB�h�&mҎ�4��z�DJ�4���=�����G���ϭ��I�r��3���D��3�q,���	J��S�HpL�`�����|E���L_�����e���Xʋ����7��F>���@Xg��`�*}/�����M6�P��8��i9��z|ĸ5����K�n6�(����u� �);�ō�
aJ+��P��0�&6%"��S��g�R!s����)t�\����xCD	���u��<x�q<W��4GV�T��H����QS`dd�ԡ�D�]��h��g��)�:�R(��;w�2^83.l*�\�i&.Cy���uMOH6��C�g#��u5��GR6n�p�D�h>�bS=��P�Cg�,���
�=�!��"�P���h����)��qѠ3���~x�Ո/��  ��>?���`��dw���߀�S�G�{R�68���@�sÒ�=���Ur���y:=5M�����?���A�`���4� ���.�������D�m��=����#Y�_:��)�q���-�Ե�=�u�d}0�a�:e� ��Uq�kXFM���kߎ��X�����I��⑅�e7}G$D�A���OՉi��M(L�m���	y��B�[%S�h*�;��y���˰r�L���J���e�~�ͱ]�+�
�E���H�6�R��E�U�I�y1�d �p�yO�A^""eN�m��'FR��v\�R��a�k���h��W>0#j�qPĺV��X��D�n�z�<n�v$n4A��DJN�����<�2p�PY���=���Q>���Rʻ�Dkh6���@B��wZ4�|��g� ��%.R�\���%Q�����HТ.[�hy�h0?9�t�5-5�y��C9�4�e�]fM�|2
��A7�@����La�ZE>��|2�D3�X��y9)�f	z	 �?�?��H�݋n��-��j�|�6�pv��b[�B��[g��S_���&�_X�6q�h_��J��p-���s9*�݆�gy#~GT��SX0�Z�ZG�2��9n{��Y��%.ymh�����D%k�Z��~�A��-�u'�Զ�׹��d&��k\d��N~&C��2�G�B��_Ef�L�4n���c�Y��t:A�7�E�x����T��	�'.Z�+Ӕ�jt�m�ɒ0M/\`Sx@������&8<Z���=�a�[ouS:z�֣ג�����ў"VHt�<t����|���'K�g?M>@�w��F����NU���Y^�(�YM,M��*��e�k>&�XL���A�q�7|E�~2-8��NӀ4�NZ4P~�_ٗZ�_���+f�=R�q[�^b�R"��	"��Q�Ɲ�=�ca\�q5P����pI��l�O�e�4�$������ϛ�P���[�_,���uh��Ү�r�W�m���� ���7�D
 � ?;���-b�/Z�D�k��C2Ӫ�*F9���!�K�&����4(� =ﶰ�k!H\hv��G�ʅ��8@�d<�
���J{ �aQUX�8[�#�%ʥ�ɗ�����`��#h�wն_�a´֒�:������`��=��e�~3-u<�e��X@r�#�e^_z�������=��	vX��	(�b�u ��)�C$��O��S@gU�赾?�<}|w0�i�,��l�����~L�c�L�-�!N���m!墚Ԩ�*��9��p-ᡩ����uɴ�캌��p�߇�����L��濏k�k�8����#تx�����A]E=t�p����,�PX���9����n�/K�	��r�'��9q�9�KI+-���$��C�tÉA�8�>a�f%E� 9Rҝp>�8���'����7Z�p る5j�����b�I�>Gyi�!*�.���V���G�l�c� P]����W���r�n����RRT����k��	shFa��ZbR����}{(02�*=SŮM���ތfA���G�)r�������>�C�Pݿ*�J�<
8m?�_CB�ZR�r��a���p��y%�{j�_��)f��BW*�n|Aw�q���������g��$���J�L]c?��+퍷��en�ϼ��7�&a�
�_Hʼ qG8W�cx�Iӳuׁ���)��SwXq:����
�s�gm�W\����W5�Z�o+z�qk�6�Gj���M��㑱���)$Ᏺ��6]f:��2O�}cTJ�|*��9{^:��@1׭��Q�P�J�J>���q5y\�~4,��"8=��Uy���з����N�Ea@�+��c�< �E�;��O����'3l�*)Xrۦu�uJX�Ј1��࢈�'�^�CDC�lP(ĩK$p�VM�C�]	����P���[�P�库�׷���p��Hu�x_S���M40�5/d;M�����gX�ks0r�d�+��9�O��!Mw�J���
��'dj7���*/DX��F��I�C�C,}85q�|�r�k�j��8G�A�ybN�[Ȫ��fr�ST'/ez�#>��z&jʺ�O��!n���J��g������f@���x�ìs��!��U����;�-)r�o]?(_	CI�de+3���N��밪�F�U�t�^=t�)I9E�\����h��z��U�N�1:ʾ`�M!s�Ni�-_�n|�G#s9����)_�9�W��v���,M��^~����ȁ~鈕^�� ���c��0�zw�B���gڛ ���0Q��
K]���8���vNP�(��?fr^g*��SD��v.��!t׶�.~��Q���F�s��ve�L��@���#{���u1;B��;��t٥rw���x\$M!F�+���n� P����|~�&�C�����DA�B��p%��F�*W�B{�и��^ث����1�8�YJ��к��f�O\�i=��_������X�Q��b���<ٺV h4�e/E�
$�p����`{����E���7��4��M�~�%Q��+�`fӠR&�y)s����ٓ^'f��N@�ƚ����>PJ}��I�_X�UҖ_��ħ��Nɛ"I���X@��?��w��)$m���`��YE����5?��)����O���q���x��a��nK��7�����3|C�v�(+c4W[�k-E��ǆ@f�T:"|{'yy���6D����*��&�f﫼��c�޹�_�q�*�#:��1g������E[���o{���BS�h}�̳�Q�s��cꖺ��<��ӓ97[	5�t���e����5��Vl�]���!�Ξpg�gq���ߡ�Lh~��z���o��N�Q�h�ɂ�ݴ�H�R[�R!����;��>�(�����5e}?�z`G��%B�x�����>�A�:����v���7��a�|g��;^�"�HWb���űDE�E���\���ُ6��n�PF��v�=2��aQ���i]W/��s� �d�$t`�M���]8��iv����2י������s����� �߲�c�·���i+Q��B�&���
<�[��5$G��%����aq���.�Y}�^z��n���L�T�I7"?�$k�HYU�<цBC�����k��bh&��Ʒ�t)��À���b���n.�"�y��Ί����X�#u�1�cjI� _���g���q���m����%κ�d���W���QbֺΏ�����Ԅ#��;X;��d�7PH��L(��(��le;�W�t@��X[��qy��u�Ԡ��H�V��n��X���b����1��hm��E��_/��@W�zeq�Gg0&!$�l'�V02V�T�D���b�xv@�@"�ڦo�Q��T���%j����9�p�8���c�A	v�n��!��x�	����uܭ�{K�Zz$牱�+1��t����:pg����w�Mv�I3&2���K6���3�s1��W��Q�݄�a��wg�}�@|;Y�&QyL(l�q���oQg����o�����\�Q2K�r�/�*���-�&�|&Lu�d8t�H����H�������w��SD��rր�����9�U��l�I.t��1�
��
�_������BX�KR&�c��o���lw�*�	1-�@ޅ�[�å�zJu��K�2�����\W�.[l~W�xc9D|06�k�y�q���ReG�� ��;2�I����ǖu�������&SNٜ�Q]�NK-5�0n�����~�M��%*e�>~d;7Q��Ѿ��H��Ә�`+Qpt|