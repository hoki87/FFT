��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#���������l��U�~�׏O����j9�PY���`T���x���s����uí������P��"��b%>�1eτy�<�gܰ�N�Y�	� {��I�ɍL�ݫ�G�R�k��Q�!E	�5E��.��:�͂2��y�m�-�.E��i�����YS�
��@�H�ۼ��nD��Y�l"BU�.TԊ�=�-�����q���Ǹ��j��ԋ����tr�a�ٵ�]�b	��%�ɔe�)rYOjX5;V��R�������M\�	D��ҏ����9c=�Vͼu��Ro�P�Jf�tRvsY��c�"n�XO��	3g���Q���^�Bʹ�7gQ+Г���$�-��t�8�����A���<����l-��*�|d7��v|>O) �(i�O&?G��m �oˮq���W& %���ʓF�U-'�����n�E�G�K�}����ߎ;���!�6��h��,]pZ������$���eSqF�%��l�Z�˱ں4�t/�EG�E��\��E�!�ʳz���kVJW6d����'������4��"��ꉐCU��9
�3_w����}�Q�8�����.x�GLA��44�SsNΣ!y��p6
q>s���'!�D�-׫�0�d�M��Ɂ ���sd(�h��r�o{Gp���,Mu�p^�e�Bp̞�(	�E�r�v�ZH��H�8CC������C�_c�H�}�ɬ�Å'�t$h�ӱ�	Ûm%4��3���1a���@�v�*|��K�y�M���4@JD���3Jk������+���*.�����\�h
E���P+�����-�ǉ��A��[���N����3����fk�����`�Ɂ��"�# W6�*g�8�7�o������(Hn�;���絬1���1��-˚#/:?��T�w>��Ol� 3r�&�����	����6��IP9T2¤��f�H���Z�E����OG�C��h�ŉ/�{�6�Y��}�=�<:cN��<	�؆�5�$P����Q�������ƓQ�30������k)6pI�l���h@�a��+E|�����g�TK�@!�c�}6��z�Y/'���n"�T��M�ku�t78�pI�`� װj����:@܇R�ׄ��W�hs[Z�wJ섴��%A x�Ђ�f����p�_�2#����;���ഝ��]��:��S�M�c.�ܞY�P(]�K��Z%ȺP�z�����5�=?
S����P{�\���JLo��K�ž
���9����c�[7�.��;!��]� �ZO��U�Ε������!�)	M��~aIˤ*+A}��gh���z��͛Z��ʃ_�9R%�L�$����E�-�ms"�W\1Z=�v���K%'C��k���ۿ��е�
�J'b�?��?C%����bj�j�W����9g��	0�d�Ǭօ9��W��N�w��K{:q=<)@k���
�?���?��',B�3@��X���8`84O8%��"�hWT:Qܶ���(`*ir�
���#�r{�9��Q�M=�� ����}��s��
��W���Ʊ�`	Ҧ���پ�>+k��2�����q˔	�ر�@*���wZV-�w�N����R�d��Qq$�4\�!k9���v1�;=x�Q�sI��
����;Ht�V���m*3I�j�U#�N/����'Iv�۝tv�R�1)�Z_�\|t��@;-�"1�ݡ(�HDJU-�el@�)/mM6�>�)���_h��4xw�~9���r�I���uls�ne2=���ɑ�>�u���.�@����܈A����N<*l�+y$�i�w����m���� b�N�6䍆��șu��]�ъc�ܤ@e@����v96V3�F�����" d���g_��^�������]CZ!��/	���F�������k���G�K��ש�W�a����ET)(��x}����&��s0ڗ�T�StqW8�Z��y�]��P,�iD�`��hK
��sR\���_ؘ��5���2A�th_Ҿ�E����8oNi�zi��.�x`:�A��@vy��O��G)Qy�hQ�$�}\c J�EŒ���� DѾ҅3xD���A!��؏V�f����d)�7<+�݂wa/&S�+��
�"�^f쪙���sRA�L�״��
3_�&�j�ٝ�:��^���b���B\+��;t�x,�'Ҙ���Y �r�ްo��-�,�X���>��I�����9`�x�D7��p�����<eV,�����Oz杄t��a&.�#ha���?�������3�Z����}�Kw�����V�9���3�</т�uaf���*��r�S,�P��I;�
6E�4��@�5���sX�I[��7%�4M謆F���Qa��Y��g��-&�
?VH�.���Ǫ���jO��-~x��K�6�W��Zvp&���o�=�'[��@���3kF�G��)f���~�A|�>o�,�n[6�x��! �F��	<>Z]&A��]3%�%Do��>Dr�ۄ���IHN�y�._�a��^�WV��@A�YR�6��=�ach�N���E(+9)>И���R��ı͵�Tt:m#(ӄ��b-l�1���顮Ʉh�G�PA)���/�M��VM:���	�x
P���t�T�M$���>{+ϭ�h��lYiX.@Vph������/��h�єp8� ��Qh�"���;ƛ�l�*�҈��$`ja6qξsjT1]H7������M��iS�9=�C߃͒%q��(=�Y�@>��Ez�J��S�5i>Z�e�Q#x0L�*�km!s�8����]�4���M̲�ȳ�/�HN)�,�1��R��l���[y���<q3^�O�H���v�K��+f
�H�a!�m�8)=<}v�v5�;�c�{��3�M�Ұ��"��}7�QV ����N�����=�7�Rɤ�M�[��0����0���9��nD�}��`M��b�@���
cن���-Ԉ������s1��?���aG��A���є�<���/t �y_�@���Ai&�������
κÕ�λ��0�<��A�C�p	V%�  :ne��]1�;�;���!���D�6�ή�1�Ȗ�HD�0��L����G�/�|-�!�x�j{���~�C�S���1!xJ�Ry|��;���$����r���@��bO����CA���Fl�����	�v(E@�UT�|�h���c�}ij�#�;j�ޟ������ Ű�V\U��Ӗ��`��
(�k������w�T��w��f�_>�}�ȉ�U�˻-����5�CǴB<��Uj���HM[�.��1���3�>�:c]&�<*q�+s����Η�\>#��$v���L��L'�S�d�E�!\ޢ����އk�����XT<��jS��_֟OSPnjp9��n�X+��
�?z��v)%1R���3������S0��5Y#^��ͪ7�o�����ln���buMJ�90�u��,���ӻ�Z�唾���sG�u�	A�Qv��E5\�����E�#5,����ݤ_�#mSG=����]�V�����0�{�x�p��a��y&g������&���)��!�	PϪ�{J�I|5��c�o���҇$4��z��m0~&� �Z��ӛ6��s���vA���(�����yh��X�{��ӵFhP���8rи�䨷a�ȱ�(���������/�vz�+�����I�\�ie#p�P�(���=��N+��m�^�z�k_譁�����	����y'9(��B�9S��ٵ��|��r�����h���	�U���1�d{�^�7�]Σ��pa�d��'+�z�Ê�K��\�G6^;����$o��S��iz��oP�9 PK0��Gu�Ǔ�o�	20Q��f;�4wм�r�t�x|�r2��Z�Ɠ]T-a�ԪHA�"r��� �p�7�^�3��ve4oݖ
t�f�o$EN�{�1n?��K��*���]O��\ymyleO�$`bԕRe�-��6	�V���P�ۑ�Ռ�ԧ�\���� �����>/t����]ډ"4U.��]�����$�VJ^��J���g�
�[����g?]�f*#�3(�'���3�i-Zm�P�Zg丷��	"�_37���>.�Ze"�89�ҔaF��K��a�#�A(d��A�٧�=,� ^֧Q��d|�M$݉�������*A��Ԏ�ȴ΄XW�Z�E��t��!��T�e �(�w]ń6�UU�w8&�hD���A�.������3�d{}d;}-q��!o�Ƞ�;Jt纑�ż�� 'F�>K�c�4��~!e�R����e�W����|�;|�\�Y훂��o�y�L��p�Y��(�t�$���|� ~�h6A5�qƸy�)�c�2#�8�2�<n�TP�Z��M����Ű�M1�`�������0���l�vI2ݬ����`?�l����V�=Ad�����H1���(@���OY)��j���z��*;�2�"�~��Xx���gG�^y7\Й�t�B��N���űJ�+^�)�?cG�U��-Q�x	e8WU2Y@Hu\�����4b[��v�v/�_�9_LB����'�S����_��k�x�&~2Ƭ�H�h��*K������#��G<Ͽ۪�
Howm뽬�S���;J����L'��Q����S�&%��#`�|ҠmN���Ê�h��	�م����B3OnҸ����"(	l{̀���u�P���T�(�J�h`7�`��aK�8o;�\�i��8�W��T�e@K^c�D���`�YhM�KpgJ��4��h�91�c*c��Y���m���s#��#��������Q]u�8���6����@f�BA͡?%��6�^q�SB9�;ٍt%��sZ��Z�'�p���ML�ف{���C:�Չ=�A{�"�#5�O[&wX-���b���^IP����2���V��=�����<�Q�V�2�PwʰIc�_����R�*ob� n�l�L�F=4_��X#^�x����B��;#��]�l&6�CIh�[J"�Vگc�/x\i����٨�qz<��ECJ��`�ɝ�jrF���]��gw��bòv�CN�N\��C>O3?����l� ����d��;>D�Y�Z4&&�8��/������+��X�ONt��AS|�r�Д[���'��-�A�o�σ��y�y�P��ȝt3!����8��A E���h�x�p���"-Q�	��h�������&�������c�6>C,!�Qշ�qjwu�W���I�bҀm-�iZ�
�Y�D��[Ns;��X��ּ1Dk��b�o���z*aY�h�9Z瑛~"I�Ed�-�����t�׌��"u��e��_U� s��[!A$hָ�1���#>�~�l)IP��K��btLc�\�f�d�y���,�63��c
��w�)n���s���l?��q�
0o7	�U����]O,���14�xƛ���'ﲛ1�$����'y�w�u��׻�ZD�$%免��ҙ�o��`���f��z�G|��9&�l�I�{����'��	���n/�+@t��{�t����g�+f�q��Yh���O�t�i[�݋f��d��X�S�_:���l	�;(��o��<�O���Қ{�6֎R�i��Dj����Ƌ�?L�2<����\���~��e/�d�jum�`��~-�Z�P� r!H�g�%����V�2�H4����{����A�����A�W\���B+D���2Y ��u}U8�S�"yز*ڵ1# M�FE,�_�XL3�N�R�M�׷���I�p������a�����xh�3�\�m~]���D�v��/q��Vl���q2�-���?4�8H�U̘�y��$�=��{��j���9@�c��^��D��Yyf�g�N�b�����D4�~�V(8.t�a7��*+h��ED���j��eOI���W��s�g ���ơ�ǒ�����S?i��K����a�Ô�T�ޣ�����-CoO��/�y}�FrAA��,^˫��|�	��5��wz/Q������;�����>+�rĠiC�Z���[�:����t�1��nn&k��_� �1n���Fq���1�اݩxU��y���j�ټ �RHOɇ*f�r��&;��g �� ~�2�����0�:S�� �6_s�d��sɌ=T����CÚ*��z�Q%���E�+��*�˙�mŃ/s���[������	�����"e�I��d��ei����)�m�Q/mߩ�=��l��Ey��r�O�dRw������&�V-W[ٓ��`H_�!��3��78�;��"C�)X�#e�zo�t`=y� 2D�h��H��3P�$*