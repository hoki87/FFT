��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ����������h�j����]*uNŝ�.�w+�e��#*
?u��X�`�β�~T�`��Y�R"��;�g�ƅ�r�� �!z�<~fi%y��@ދ��X�N���C�͗f���f�Q9h����Ա�R�^-X�.
D���U���ǡ �\!I�=�^8XS��ҷ��}���ec;�'�m @|{�2�\�%��j�������[��١�Vp���RD��눅p��R�u	̥��e�5Q��Pr>��'�B>�k��Z'Q��m�6�^��Z�}I�m�SJ��y:9�6{���sF�h���=��jN�(���'�M������+�v�k����?r����\?@���.:ǲA�<O����m-}YT�U:��ϤM;����i�r!�z��}z�
(2�1vǻ[@��:����,�	���5ى^�$���9����
	�n�2���ߙ0�.��8jŭy��O"��t�2��'�,~˜gD�%q�Y��3i�}s[��C��Dm�~�/��(�RY�#0yEQ�qs�����uɨʞ\�61oAI�9�Ic��}��h.���f3䥸wT5�em����e��d���x�����X��GV:)�6Y(N���6_I��ח;�I1�,�����!#�鍥��˭��:��f7��uԅT?�q*h'֧��A�z̔��/�ǡu(4�*��V8����Ɉ06" �8x<+�V��Hm 3\�23HlaQ��7t��uQ��f�C)��eU�PDN�]L��$�He6�L�1 �C��	��e݄b��iX3�kCɡ񡸦�U^��}(򸖹�̜40JZ�Z�i)Nw�b�-İ��TK�}y}��m�S��>q��Y�RK�e�")�pN�Up����:ˁ����ȎG�ބ�,FQ-Û�!��XL������i�5�X)ftbN� {����+�h�N��,���t?.�Q�k��ÜPo`�"z�&'1�阈�+�4��9*n��Q�|5��_��#���Hγ}C�Q�
��T3w7������s�w�ك9��[+���I�jIE�TC�Yu�r�&���H��a��z�a7g�1�ɉkv+��XT�7�Ow:��9~ �b�0��WҘ����NO=2�s�����?�� j^�����@���d���q����T���ZyK�Yl�Үa�
�s��gj2bEO��/]PS��\�9�*�s����8d�"�����y�Ђ<�ĭK��<d�HW��[�T�P\�pb\�o��L�`����o@I��c��3�$/v֤$�{u���J���Q��
&�薙V"ZzW�b���
T���,�G�~��( �`+���'��qbmO�W��1��Z�P~�7���pqO�ru��ҁ�Z�o���:�l���T�	Va�,�W�>h�f����L��tIP�nq����p����G�Cz�]R�F�V+�\_/��������P}z�D/���u�Sr�"ʎ1�OY42�d�G�L-�����-����g�7������@M�!�����͚�%'�I����kvGW�qނ�+E+�{$�+ղ��s��΢%Č\6��M1y�U@m�Pۯ.��r�����}��q4��̜.��T��"��O/H�iG{���:I9sh�o�LN&���U��Al���4�ƃS@9�=�K^� �?d_i>��4ӈ��hkM\��^,BTZ�lm��_跂4��A�7#�f	B�
7��L��S�E�љ@���C��BD2y�N?�^�y�;eۚ�͍�N?�q≆��K�؊�1g\�r�5ZƟ��}��x9�`v�2.S8K)L�9�z�|�M&a��q�p����3.���=��#�I���a�#���� ]iV��կ@b�F�j�ֱ�����������3�U|��C���Cr�$�5F��E|������]B4`�������t�.w����|�ָiH�xS꿿H��Ts���(���4�<�
'uq�?�aʼ��&�>d��vi�a-�Y7A/�� {/�DM��ɍ1(�ͼ����ݏ
�E%(��9��	���1ņ�گ����I��ΌN��z�_Wz�����Bl��?�W��)�y����*\�=���b�mb�ܢ)l�7�C����V;�{��(��M<�	A���J�6VV��{�1{�g��l� 3N-�=������Q}�V����YV {��^L^�[��h����H�om��O���(�|�"_~�k[�'*��#�+���P�g�9������6y.n"<���[�c{��J.��W�tQ�Ks}1���F�^w�m�� �TM�!�es@���UۚYx~�}Qz�q5đ��|P���k <l><RvSiPQ8AU�%_p#�o-�\Q�A��?���7���gv�e���f�7? "�=�~;<��c����
�T�x�GPTV����	^�U��'����Y��Q�p	{�c8�y�B��o�)l��P��I�պf��������r��
[��s%"�1��52	Q����B~����~��ʀ�
�I�
;���	G=�p,�J�)b�C�v�-��w�x �,1q�茖��
õvR�`B�ה߯B���`Ma>Pε̿�Y\q� k�9}�څ>C�|�&��S����|f+-s6I�%{`�
�k/Rٓ��w���Fj���g��88�g��(�YGU_��n-�T��k<bq�Y��r�:�{���9�%_J�Sg���*�T��@�����/�m,R��D&5��O4X��I��Fp�7�{pNX�����#�J~��nf���UӾ���:�y�D��.��IJr�찏q������D���Vb{����8{���i�X���<�l>*n�P��)�u�$���M�fX^�|�����l�U@5	8����$��?Ϋ�u��ƭ}�{<��v�ѺpEn@���i< uxIz��ջ�7F[��`[Dm��Cb��f��ަ�k�Q���{�OQv%J"�4�ы�}F���X���B\@�$�T��b��*Ñ��[����4��:�d!Fa�����l���"y��3�k#��k��SR�Rţ�.���1;<DfҀ!� ���`�`�V�Ƙߏ��4�+ҵ�[��Sw�2�DW�6A�	�2�D@� ����0ô�dI�{��W�]_a�,.��z��;ؗ��-[��c=1x�=O�� #��:h�;��˺E����",y�T%worw�.�,�4���BGig�0?q���24���������#�iG�:.�� ��W�e�m�✱}%���BL��%-����C%���������N$s��`l����5�L��MDi���-�zG�������ͤ��Ϻ��qr�]!@	Y����a��߉�6u���˅�`ގ,�B$��� Sg�nT8��7��b����*Ǆ3�����O3�/�0]����@ ���7�����P�mYA�2R"��w��o6.�=���]7�<S�@�X��m|�~��4U��U^��̅g�ۗ{��3�D=��l����:��J����J;�����2?���*my�.+�Z��6"�)hX%?�4��ļ2�
�X6��m4!�>�'!v5Y������S�Ʌ�`��T3�ay&�/�~W�����v��_e�LZ��W�V�S?5d &��0R�v/�?
���xg��ez�&��/���ye3�����@su�qcv\m2�G�ע�\���-H�%��Ý���l6t�q����|��}a����F_��0���֣?\f�\8�p�Ҩ���8`�d�n$�68>��,���$�<�c�`=SBZ[����\f�oeB�U�.j�n؃a�GK��Sq&$=e���ӵ���R������C��Y��"ګҡ;���"khi��U���TV�OV^vN�J~����{5����L(Ct�Ml!��01�Im���Ů�\�Y�|?��6����a��Z�A����t�Vf�Ӛ>�Y�p�F]+k���Ȇң�)���SU��>����y2|0�>�ޓ�v�6�� I���~M菅�Փ§q=�FޣY�A8���X�*��K�����H�'�E+�6�Jo��;�$#3T⚡��` ����?>�e�O�c\�?���/f��^��w�lw�I&~�|����/������l[�ǄA#��p?�)� Ā�l��n*S����k�l���p���,��?�t@V���C91ŋ���րUq���Ty���݅�����+�So���7��"�mn]�"�Xb��R��D]n�\�E��m������h�� ��]F/�j�Z˯?����?��������Ë�c��j���{2��YT��z���ņħ7���b$�6�1A��{� "v��Uy�l>�j���Eaz�?�_õ[?f�m�-B�I	���<��(��ٞ ����/BZ����DC�����TLqI5����f�hcA����֖����{tW�l��x��x�U��P�͛?]�z��H�BZ[qWt�lmK���n���4�Sn��<Od�
ެ6���g�u�G����5l�����\�C%�TF���e��ڗ\:fl�lt�	q�d��8��`�7�C4|X<�4��Z���.�t����qv�����qfA��/�