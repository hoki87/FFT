��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ���������|���sAՑ�0}V��a��[�#�r�LՑ�s����C�Zp�-F/5Mp�_��͑��pz��"����^Ĳ(�}mW�݂"~����y�Y�~�-
@M��Y��P?�����-�9z��x�|E�VUݻ��6eY�v��֯ބQ�h���&m���������:��h��Ǒ(V����Y-Nd4�ܝAV���*��lz�Gu,�i#!�O"y��?Z!y���P@��mӸ�f������;1�H�֠#��c�5J�\e!uJ�SE�G9�Ӣ��vV���"h�,�X��я��+G��C�����K�Oj���t|�̓_��-($g�Y�=��0�6���O�� GR#�vC�oL3R[���N���7���& e�v�Z�4�	�Ys,��S�%���qm�X»O(M�(7y
L���/�W�M���s��b���� ��=e���d+ջ�+'��Kc>Ƒ����[j��r���u#;�8Ny�,R�|sD� Mr�
ZN���Q�ϵ��d�F�����
?�ZzY�F��N������`��;nԱ�@] L�"����?&_r�G۪m��xA�^~��ƿH�zSr����s�;~l�D@�^ ���%١
�}�	%zE��N�����,C��?��o���}�����S�&��*��WUg'�|����넺��"�K�a�\���������D���&�XeU#��Ka��!4�����z���J���S"2ڼ8p��@�0��D�R4�?����vi��<�{
���N�p�����׈o�6�^֊{��ʌt:gƧC�]%�[gS�)��	��|~Ǧ�sy����ܩS�1�RP5�Q_�d�j�:�Y_�F�F:�:���tt�p�Ka��v����T#��ijd{�@Uu@�t��!b�<�w9��tkD���"�_j.���Z۱�8bZg���O�ݭH��P�����:��n];.�
u����"z���+����y�\(ic�#¦!I�ERM�:\���Utolw\�T#kx�t�D�r�g�����}�Ůf���4�����C�Z��	��F}��1	���d:�s�n��YdP,!c�-�e�>ڒ�>������
Iv������ߐ�ܹԭ�"�ƺc�/9+����"�%���2:_�a�g�| -��FaoF}��f����Y$�}
��ޒ6V6.D����|��(c�>#�$_J	G����d[ϒ^����$\�����Pr�/?��09�O�X/�����}��