��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ����������QF�4��p)Od�,��kBxZ|u@���:I����Oi)yȹ�������_D�����'�qS����\D^a㰥��\��_��6��	/.�t���{E�~D�R�5F�_�p`����V �@}��'���VVŘ����6ƥէ���6��T�ä���4�w�i��2jZ/�FT��*V���}1�.�a��x�9�
ɶ�UI�w�]�����\��/+id��q�|&�(���:@�8}]�	�	�>�x�v(&�R����Jkk��Pf/Mg��9�L3e��H��m����5;ٖ.L%?]8�&x:��D�EQ �<6�ކ=��]���#,���{;N��Ҽ��Gǅ=O�L
���F��l�+H"�Q_I�,����r2$��c7ꈀ�7j[p��p7"`���9��Z�u�j.G�Z��;'_3�^7�&9��F�\�1$����>�C���:�y^��ς��3�LZB���:�c5Q�;�׮�ܓ ��vo#ؘ�o�Aj4�O�|؊{qq�㭠�
��5��� ,d�Y��hh6(�_B�o�0�S�����PJ�.m�Bk���/�i� ��j��K�:tI�b�u��WC�պ�IA����KS*��:r��I-�9���} 2�ǖ�M�X�!2I^�f�q�(;�J�D�aYVm���W2J=%�S����G��1Ӟ�<O�	ev�¤���Y���z3���D�U���$�ճ�Y*l��ɑI�M��,�L�����܈\&=Ϧo���t�߶A�zňl�X��EB,���Bƽ�����E�3�����J����sfC'���@��l��ۚ��[�Lx�71C�rp4z9S�
�*c��mӽ��\7�_o�M�V[�-��bռ�#�k��7Y�mB�1�F� 0T���b_6��=�U]�t����U$�_��2*g���l�Lp*ʲ�VH�w��S�05�Z���nr�ޘ���q�7�S�n���#�t����)�}�u��'��ޫ�أ�E�ÿ��\������Y� ��"��������dԱ`9��7P�T�ܥ�R�{{{5��:D�3�f�**bw��=��<8�0�A�7�)c�$��џ��!����H�j��2>Fu��,���:9��#���j#�f��Mq�^���AY}Y����8�$['�&���5��c��IO^*���L'�9F2�(��9���<�9��+�dYmxW(�r��)<������������	�kwR����q�mS��L~b�U`��x3\9R̽�M���
${]g����04'=�ڻ�@�٫5SZ��	6elA�*�r��*y����޳���/�
�?蛎^]#w�?̤-u��؝aΝ�#x]2j/F���a���y9�x9��̅�Ь<���&��޴�vC&q8����kz�6�r��
�)��G���2�+�VZ(0���ܞ�T�K% 0�X���