��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#���������l��U�~�׏O����j9�PY���`T���x���s����uí������P��"��b%>�1eτy�<�gܰ�N�Y�	� {��I�ɍL�ݫ�G�R�k��Q�!E	�5E��.��:�͂2��y�m�-�.E��i�����YS�
��@�H�ۼ��nD��Y�l"BU�.TԊ�=�-�����q���Ǹ��j��ԋ����tr�a�ٵ�]�b	��%�ɔe�)rYOjX5;V��R�������M\�	D��ҏ����9c=�Vͼu��Ro�P�Jf�tRvsY��c�"n�XO��	3g���Q���^�Bʹ�7gQ+Г���$�-��t�8�����A���<����l-��*�|d7�庑˓���[�8~I����C��k{P�R��W�ġߚ��F=�3�DU�{���G���<��XgXӥë����!c��o�#Z�dz"�T�"g)Z��g��&-�ܮ�� �fv<z�o�X�vIIX�
9�G#�i��U��.�T,n��%<M����ƚ�u�!-���� �,�y+��^b5��{t����1���1��M*�b�W�հ��<P��*��3��,M��>�י��38�pQ�ZC��Z!#Ch	��d�<�M9��0
�=�A��V��ω���YO ��Z��� ?\(��wHl4\X2�$���Ǡ<�7DxoG���b�]�1%��~#��q�W��o�Oۼ
��%r;jh1n��w.ۥ������5QI�hb넷�����]�ƭd��*���&|�] �y�����m���0� kcG��r��h�P`l�|���������c~��	�J��׵�z��Bk� �֟"�V�f��hM��3A���N^Q��Z��l�:�I���3������Y\>x��q������K�����t��$w�%?���?�Х*d�}u��� q�.��<Vk�c]����,�Y\�O��XK$����YT%
���:�RW�ZxN�h���v�vp������/��ƀ*�hn��������,�:�#���\f/���#��-AL:M����<	u�"���r�G^uz8�;��������1,=��1+=`z��KPà�w<xeќ�d� �le�Z7��DIr<��3x9��p�tǺ�����2U���*NA�1,�w��o:��t(��rQIR�ޮ� �T7��Q�%N�7H-����zu_�c>�fc7��)F�Oz0.a��N�Tz�+�30��2���MVA%�u��}�.��^��"�^*+��b�"۵����^��=Ӊ�d�
�֝QP��=�Ɯ�Ի�g��$��a�_���U�hع������_iNp#w�ru��]O_h��-�����<�L�\�J�6�Ӽ���I1��T��������Ω��cZU��Rk�ݳk��#k��b�B�`�9��a��[
f=o�b��
0zƽ�l��5*׀���7d�˄���=�2Y��z�ӟ����ގ�@ՙQ�Ix��r��6�&V���U�i�������Ib�P��
�d ����0�?�j� zԬEӨ�T)5���-`��V0UI���/�f3gƄ�[�w�ծ�����N�~?^1�bN��)7��'��c��)�, � ��\�N]�p�=刦1e.���J��*֜�\��:��*Vi*_��G.�H�N�a�b�49¯�Z�ݟH�x�猛�GO*�� ����$��<֞�����6��ҡ��k��t3��:��Ь����!~������`D愲Z���&�j�/����as��m9��}3�^��c�aiPyn�4��`;�4kP�Z�]�f3�'6����c����e��º����� �ok4�ܬ�9
�:XظvWksǄ�k�+��;�¶�~�@��*�hg����{�4�i��(�yyv��sX
f�5 �+ȋ�\��ST�ʁ%���D� 
�X<v��>6����d������B�̒�����\����M�.Z]���2���S����V�1;�u�u�ų�W|�hs� �B��+�#�����S߰�h�*����1At�Ӝ��)����|^yJ.R=Ms��|>�B��=���!�SU.r����uޅ����&�F��odE�[�?Tj2&�y 
~�8��1�Sʠ��M�ݯ�3&I��yV��
D~��T!Ǧ����3��I��،���}r��Pz�۲�(�r�:���{��#{#�M���v�EP�d��]��d���g����8�r��4��^�;���
�� bO$4{y���9�c�$\��i��d�ɦE�T�z�MAv_�V�A���3b5n�(�Y�2��J7�"��DdMz!l��P%8#tN���6n��鱀�˝���0�c��/l3�~��ߺ,K�U&څ�;Ǭ���S�����;N��:�ɛ,W���;�ԭ����I=�~K�C{��3�)5�ΌSXq~+E�<&��l`�tn�����
���P��V���cr���zO��ȍ@�ޤz�JAM1�~�j�Y�>��r�G��}��7Yũ�6ޑ�P�G�Z�|R���|&�5�Q������ė�z�0��>"�����}�8�q;�@��ˮ�����2��ϭs���A`�2 0��8I���jS)y�yf�z��b��;�f�Q�`�Xظ~y<�s�*Y\�Oh�,�K�f�+)<=x��0���{N�[�_��ZE�,A�5 \��M�7�6�_�a|�|������#���E�󢰵p}����|HV��t��3qW~�[h�h��z|C�����Z��Ĥ�QDr��ƛ����]1;�(QJ�#!Y���v�J��ʞ�i�0~����a��|5�9��͸T���ᴉf� �6�鶱�oƹN�����h[u� �"+X�V�͢��vEm�?7:0�xk��o�k|`3�ە؁��5�i.���+
G>��S<_�OI!�(�R�F2��zۋ�������tc�
D�yx���i��=��lQ�7�ȝO��E|g=I����w6�Jr'A�V!`�j�~�ytLܪ��_�:X���v8�e�~�z̜㼾��g��pYq ��C���B���夞PVi�Ǚ��m��T&)�sB�L�����Y9$�<�<��2�Ā��%Q���%Uj4xp5��U?�ְC��,SL�tq���B�6���N
�ի�����-?��nn��u:쁝
/J��|�Z(8^e;��h��66��a5Ǝl�U�b��p���$X��F�H9�.�W�J�L�����g�# #C�@��ѽ�+��GEK��j��sb�,��޲��ҝ`���Dm����������N��je��+qV��8#�ӵ>�z���K�1�0�� �4��u�)�~��δXs]BVh8��XD��'r���<֞r㲶��8ʒS�Q�)�w�H�Q;G��)�?�������H�v��"���P�cP�z���!��j��Q+�5YYd�p^a�P̎�a��xJ㫗���P�ӑ���~4hM��oa7R����{���O�$�_+�H�I�W����W�0�A(��S�������,����ŭ6��JrF�swUX�E`��@��a��% �6�;!bg�'�Q�C�DhU��
\\���b����o�[�ńr<)D�%f��V���\���{R�%κ8�.��=����	ur#`Q��:b��k�Q���lw�7@���y����O 
�W�Ȋ4uV��lhy��� ��2�u�
UsJ5gl8���d纽�%>�	B@h�9=�?����,wA8��Ґ��0y�����ě������AI/�\�±|,�y�.���������.�k&��j�-KI��]���<�E�f��fgk������Z� aʉ�xV�2�F�Z��R_֜3N[����⮐��&���HّL���e�K��T0�h<^��9��˝w���B4W*�ϰ!5jt�s���q0a����X�Q�vSj��*P��q����p=��+�	
@�Lg_�r�h38+�:<����c���:E��W=���o&,���B��O6�@�V�Bh=<m���y�X���[&0|0{�T|W&�m�����')jA�+˕����H�"o\�d��N�s��:��s1e)X9m���k~x��Α;�*Wd�2��I{��rg��4�c.��.��P�P �SW> +o�2�����1�~(�s<����N2�AP�
�f�s#S�]�H��E�z?��Z�.W`(�0#`5�G�Yg�|�ձ(���~���cd�^��:a�Ks�ނ@��Jk����$��z�U���_ ����pc�ݢ7�T����Tl�@:�s?Ls�f<q��(��QQN�m"7����l�>z��$t *z�Tt�� ��4#	�Ҭ�~�pT�^�s��8;�9a�.CdA�z���f�����I�TLۜ�'�8��,P��Dp_S�G[������9�N�����aO��¹��Kq.�p<�҅Q�u�}݌�yjnhR���$$њ�§�8JFˁ�����j��y�c��g�&u\���$��݄�����l�Q�~���*���y^�Cg�D���Hn/)�H�܈�{�;K"�g�bIX�SJH�`RG�?2�f�^�����5O ̍Bȍ0�垱,�
�_L�ǚ鿦��}<s�]E/j�7�Ƶ��.��^e�S�'�#��1;�Qi�Y�AΉ�H�I#K����2�n����'/���r9� �-�u�9�
Wq
����� ��0�� _��	"Z���n�`i���߃����J���!n�J"܂��*����],�Y�PKE:s�w��x��Z�s����HW���B�鑜9��Q{ɰ�M�ς>
�	��؍UkƖ����{�B�|nkn�_>�z���<t��D��P���z:�D�@.�W�,pit#!i|Ik@�C���"Vq���-P�Z��є*�>�}}��{���ؒ��j\�<W{�&�Ү((�+~<��ө��IS_T���kVU�p?�f���4^�;��v�<V�]��26^��QPX���F�\f�Dd�t"C����>����5�vL��~��\s.�	�a&$ă�j��-��3���v�D�҄5`��"jZvÞ(��iv��|�L����}�m���A�d�$d6iJ��@*��!MV|��Qh�,�+��NDE�0d޼����^Li<Fa�!ȇ9��C�H��iJl���*��E��z�r�eفۙ4�&�0�A�&`��d�4<� �Z�{}&�V�"�-F�:ph�6��y��&WDB:�KJ�-��cxN��r�ci��)�?`��|�)}��Tҧ�7��F/ z�R���Au���:n%�tT�>5mPR�D	xV�rj�!��۩��5<�B4i�c��|�L��<�W���o�R'
ƙ��0m�em�{��Q���lݦ&��H�q�J�zl����4��:\w�xi}Z3%w^��$s��c��g ����i������a��������/�ުN�x_��"`�w�O� ZF��3�ca��O�Ǌ�s4�M��H`Ǐ�3�Ľ�X	�1�`)U�g �O�]�i�8:�[�=�k��V�ՠ�+��%�����䥓��uߐ�P��6l�Ŏ�n�y��m��R$���b�,���1:[^,�z~���%��.�';�a��P*��������v~N1���K/�HV+"^+I�8[%�Y���`��ߊ\s(�[c�6k�$A�: p�,ҏ��)��r"�tS�b=�q�я�!�IW��OhXd"���p|��<Y��y��#6T�wZ���밧/�5~*�ŕB+SP3�#0�Z���������/5zڿ��y.�<x�z�ǟyh�S'�w	��x�OR��+?O<ĄG���\��<�.|�@��L*b���wj��QҋZdu��!��M>}�#��!צ	�@*���:Q�`e3$A�OH�y�X�(C���c/ho� �5۬��'70�n;?j� 6��!�G�ى��0�to���գԿ�=�=�;4+He�bջA�jEު0�)�����g^�����c�	_���Tf�d��W&z�gb5g���"sG��߳�F�b�Q#��iz��)��@S1�ި�����voˊU�:�J�G��^������~Á�ڈ,0,e9�3�=ȧ����$)E:?�I,*��i�W��+??�#�����\�Z3�%����==,��(�#E�M`�(2u?�I�Ģ�)ۜ#�����&�5��d��t�Q�z�I$�j�v��sRd�c���N�]z�	,��I����M�B����� �A=�ϰd&�Wm��L�;��>����4�>��~���"������
�7�Ʒ(�α��:�\�`R�" 5����������B�o��\SC�,l�c+a�8�A�P��1�]V�4pС�?~�� ��Tu�W�c�V��R�61u&p��3`>�;[d��;N���Z"��إL��G�9�,q�+]��(����ki�͓���t�����U�;�vc��D�Z���I����,E�5R<�z�����p�9ߢ���V��5i��wu�
���n�cf���б�r�d��u�k�o0U�;�Eaߜ�����H�O���ɡB�c�=���/�R��7 �3��w֞��~��i�}>���4`Սz��ƿل|+���nR�$8�S��B���n��_N�B2c�g�e�Ta��C�7}���F�+A�h~��2Q_�|�NRȮY�K�o�Y��ҘM��_�:N�����?�F��*S[��̭��WR���c@|6%POb�����[\���A����Â��z|�|�b��ЛX*9vo ��Ҟg�9x��Z�z.�I��N`X���N?��<��Q��D�C��^��Kjы�����Q��A.�j`V�Wo��~�al�L�{���XGf�[%b��r�tnJ��d�_6�z��oRI�a��gQe��7��t�z46� ��ح��pl6]!�\�Ԅ��a��%f�8�Hj��G�k7�_8�1����I��M�׵�����\7��'�=�e��j��Cp�:��D��G�9�u�,
�Ah	ꉒ^@������̸���*��6��0Na'eHj�FPk�Z�J���)j�x�2�Kq����.��7����IX�JtOց� ��h;Vr9e�Ϸ��g��	E�f�o���RK����ޟU�x�꽬��}�=���}N�7�ʱ��6��X�e&�QZd���^¢��;Q2<iO%�c��f:��k����j��:"���߽X c9
������UUw,�b"͝�QC �ج;���+�Z��;e��y6�"š=�a�,���]���_Q��}3�u��E.|�u�?%�@g6��%�%{@F ��? �į	���9��X�^�5JS�J���X^wdt(�vpϛ��w��t�
��7���v�o�����T38��~�4���1�83H�r&�'������Ǯ���aS�<Y����t@=�W G=H���<K�T������Ѧ�V!�8��"�
Ǖ������pk��lC�]*�}Z!ڢ�[�\��������,�Ïp�3VO�H��=O����x#&��V=��Zd�*�Z�x|9��y�f���v�&�Hs�^�e��خ�CU��4f��l��U�h=�EUS:�����ߞ��� w����=Xn����*XP��VlS�q��~p|���O��}㤾���uH|n�tlך���{*)�J:9�����\1�ß�yo� i0//~������d-�0�����O��� z
Q�N��w>"m���/9?�ȼaRz�zU���pͯ���8�(g����rα_���ĖZ�3�Iu+��%��V��vȕJ�Ɩ@��-I�}���'�F��Xh$a����:���ްQґ<.�}�t&��\��m���㈋P�v�1By}�|I.�x�́�h%�ԟ�+�(�1��%��=�Ⴆ�3R?����Qr��m9t���Y�b�?�M)�q-,ni?}��<"��)`����DE�h�0+k�-�q�|Y�&�9����69LA��ږ�2dl1]�>!�~:,^�:��;��d�j��&��)��$3yB*��2�z�/Ӷ�܊�?�Ѹ�������:SJ��W�*��K�v���}�#�
g�[?j��@Ȼ'�O�O�'�^T"�jq-�;��T_$,�ǟ���y�19O�;ځ	�O���A(|QB>�?Dh��-.�(nU@Oa&>�Z[�f��4m�L����7��O9�@:+���ũ>۰Õ���G��o;�ՓA�I��dt��2<tw:yVRl��O)���o.��'#a���>k�U6+�.���M�(���	�:�6� *�%U���{F�̌�)�4��7�T>�=��FK9lp �o\�T����{hw�#�O��U�R&�.�\�"�8*%�K9s���;p-ly��K�L�2X7��1 �SF�6jɶ��,�W<lP���<p�.�����=����`��X���J�V���^��<���.��w�����Z/=$�5I�p|4d�GD��W2ݶoX�}j�) 
�8�����!�����2�D炧 ��ԝ���_'�I�TI���@i?�Q�@��R�Ҏധ�ŷ�¹Qd\_�B9%�L7�@�u�b�hg�G3�>u�wF��yJ�Z�SB\*�:oS7H2��v���?��]{��w`9��yl�����xl)�fe\�ڵ�Ĥ#ؕ�� ;��b�� ������D��6Q�ﴬ1�E���P��=fzڮjw�Þ'F����X�����X�ae�aVV�H9�	�ȶ��)���KSd��/}���r�)X�h�}3t10�g�
��&z�`&� �X'��lhk`[d3�xB �U�t9a!,��x�i��{�l��y47iY�B�1ז��*�Ξ�"�_�s����a�ݪ��֢lGZr9n��b*	��Jϐ#j��)�yɷcb?�a�h��g_'-A�^dV�H���Gt'�2t@'����d�@Y�$O�fͶ�������Tc;�^�ٺ��|�Wbk��'�A�oK�S�5�9��5�ژ�a�!dV�ᤔ�ʏifY�o��� U/�іrm�)�̿�^ �<�}++H�/�!2����F��O�W��)J`�N��s8�R�ͭ�!�;��z�?��8�y̕G����#�1�6�$������6�9V�z��h���~���r�aa�'��'l��¹1��sꃉ�y�U�Z��n�ߚ.X���_�c$+j2\[�ٞBjCD��Q���Md��c���h^�h�W%�qK���6^B������������%d%�S��8�:�P*T[[	Mp�W�r_�Tҗ�{4+�� %
�;���-�������~)5�~$�G]�.��_y�`�8��t�����T�eԭ;�|�N�3�iD2)$��ɶ�~y�dϝ*77��Ֆ�#GTۣ	�X�g֧C����[���+�0yA����uT�0A�ڿ{'�;�ܬOa�~��}D(���X�Q@���ﱃ.#��WTQ��FSRE��;m��S��H���g$�a]1��!��퍻�Yϡ�_��H��kh1K�U��G
I����Qi�רєd�;K��e3Q0_���V��E�p�LeΠ�����1Tߕl0,r�O�-�0D^��v
Z�]GX�G �����y�],�>?Yĥ�|�(Z�:���&�At.�U�{��Hx���54���]���SP��$YHd&3�^���'�m��졔G���9��R�#�0o���ឰ�ð��oq��G�,�(�c�x�^]�pH��I��W�T�	c���_/ax��� ��+l);#�����3b�NƑ�ڛXf;O&;̬ �X3��D�M;wW���34m$%��Qb�*� S�]�s�s�JZ�D7�!6J����=��\V��0�}c)%MQ�X���_/c'���o(�&C�:�B�f�j���uI�+V��2��`q�X��P*���x�Ҁ����RVV+O������`�a��RM��XP�XL��Չ�o�F��낯[�f.�x@u`��`
�s���U�!t̎����W�����bFI�MBgu��f?�Mm(�p���E�!��[�x�2H�-)�
Cf�£�n�X�j�O_e�t����|C��+�����w�W�z��j��I@-��a"��
�|��m�d���tm.�	J2�ؙ�r�Z^�4��t�T� Ci�"��iU�ho�7nj��*�F�^�@�U)��W&f�g�v��0�ɚM-��l|~�qi���6#]Y�H�xM��wK�=�_9.j���ү�&;�ٕ�<���ίO53/K�N��"d�fs3�V�T8�"�4Krf������\��(@�z2��Q?�RU��-�.�i,/9�U[՝e{x!Nm=ҋ�c���:�ϒPPE�d�+ޛ���i4��������5���F���Y��U�#� �4G5|��Op/tC��g�z#]�;��ٽ���m�[9>�T���ƅ<����F�f�^u�\����%8�#hK��J8W��7���r���ld��o)r��{J0���V���5QI�>�^��e���¥�+.j��*����9����"ơUD�0?O��>�g�/.�s�v�m8��.�U�M� ���������F�8L=~9y�V��W��5D�Iο���t03Vy��l7�Z�����I/�۰�����D���ad`w4n6I���5�"�}5�����+�LS|�B+��K3� �r�v�ŏ��:mzA"`x5:���w���:��dg1�]���nֻH��ř�"��������K��`q�(f����~��026H�?~ز�jݥ/�����ൈ)����m��ɻV=f&�⦱�5����g&�n�7]���װ�KI�&�2"6V`�|֙��֢�	�߲��#n���f%8�;[R6���ז�<�&|�c=i���|g�CH�1�u���qf�{�TǢ��ǘ�4)'G��������b���bI��]���b�h��v��2n�b�b-���/9/alΌ���zm@(��8����:�L<��I��r�"Z�;���o0^�����jq���M�9a�����|l�X��x�^�5�l��]z6d�u��m���UqIG�759�1�̀��j4�~����Q���*,����H&Xcf��5�����o��o���,�<���9�����ˎ1A����K[�f?���4迌k��I�?�J����?E��47�Ϊ���b�'1�xЈ�M�_�Ʌ��{Y�M���]�R����BP��+C;�����~�Χ̀T��>Ov�+��Kf7��/�1�V�b6�ُ�?��(k�w���}]��U�K���.#��C��B�~d�A�ź�&om~�u
x��Z@�oM� ���" ��؏�L23˘e7����0�t�}Gp4��-c�icry�%��m?��W�^����(庸A��-4�z��N������dv+Bɂ.��ԛC��y�O���a����ƷiD��V���w��2B�����$��ّS���1���ޮ:���BQ���a(КXi��t����^��Ӛ�v�qŰ�=)��p9bJ��bڗA�� ��
`!
�������L-�4���0"Muj�����O�L�O������W�M�?O����8�n��R�Dů���/;c�$�-V;e�z�*̒S�g9�w[��P|&FŇa�����	*�R��U�"���Q��������>�?��|�VE��4��v[�YL����"��P4U�x�1=�n����߆?7���Gшq-Ƀ��쉺���:p�K�P���</��`��a]�����'*Ւ�8�<�
�\i�J>.���M��[��T�N#�W�n�C�W��w�	&���#��*b	��Q&T�I&PB&��7-F�.�6�ס�A��+�;Q�~n�ٌ�a�~5'?��/�����z�oF	�	˝l����]�����u4���?]?�^�y������*�{�k��I�Pm0�EN_�oPt��i�QS�7f$"x�$x�>��UvzEz���Ǹ`޳Hdn�XN\wQ!��M� X�3���`��9T����
��+�W��۴j$�S�����R��+=k#��� 1i����ɢ <J>LȉíA'FS﬒�O����� ��x����I�>����{6�?x��[���L	������\��Ɖ�נUЦ��.m+���TF.�]���pv7:K��M�WDJ�!F�)ϟ2��c
�}�Ɯ��iU��X���f�T.��t�g	��9d��\l�S���FW{!�N~
d��.f&�p��,㺓W����d�/�ډ���@�s���(���v��^쥲<��%ڗ�Ľ���<�5�B�ofa�6õ���_>�Oq2��>��vfmt�}tf���tW�c���ZX�������!Y��>}<f�$���
��=�X6�g���_��E�>����|s�ẜ��.)�p~�aM��/�I&hL|�o^�խ7Oo`:�R���ګ�tѯ["¦^�:��:�AbJ��V�M��b�$�����&����cd��i��6/3�$�d�9���$�.-��f�y(�S:?�[t�7\�������6]p���3��9ݭ��B���P����r7����H��$�[���=fתM��V�4��l:�`���0V��FD[�xU����Nx��q��uM��&��&��}�Tj� ^qh<�Y6)�~�H~[��`@=�D����CuZ�V�B���I
��չ,��� Y��������a֧<rf���d�(�<¾��}xy��`��T3��)a��Es3X�$�t�`m�7=y߲2�UK����)����������S�UX�	j45�3l@8�̖�+R�@�ݵe\�t.BZs9J�6��(�w �:�N�i�ÀѼ8uy�"����2��ܬ��(�d���$0�]*�� �p�i����h�����uA6��H�Ъ��#���� �kk�=�?���F�}��y�"F�֜�4����ZR5���.hE��.�|���(~�N���}�QeMd�G��q�"���4H�y �s�j� ]%�G��?�hK���oP#R��y �����D&�P�,�ŧE��d�n���Ob�_�8�tW����[� [����%9Hx��\p_dȍ�g*�q%|�%iQ8c�9= ߂�������L�������'�	�`��w�S=��x"F�2/N� BY�8j[\%%���Q�:��Cx	�#�AS�]��|ϥ�c>���}τ�����͖=�{�ȇ�޹.�����EoN�2�& ���ޤ~���J�sk|������Q����nAB�BqϿ�c,�dB�?�He�ʂ2��5(��8�%rw��O�ZҬS�����@��6�FX��?�VQDh��PfMT�cu(_D��~�-Ε���B�<�?���Y�@��̑N�ދ@�������.�}0A�k���"v��*<lܽ�������hȷ��d��[�l`�"���7��JfLU�/Ÿ��J���&A����U�e96�D���3�Vu���~f� -#��!]�=����/ى�=�-�FT,�0ݬ�K&�W�ڛ�1�i� =*Ĉf���+j�[�z��À�3���02mu��!~g���Q�]�g׺Ew��;��YD
�R��ۙ7H�\��N�0��{�[*��B��;��V�:k@g0��&k�tZ͜c�Ǳ
��M�����t�Ģ1p�=@p�-��$S`��-S<i�
�IOh@�{��]�qqx��T����Tuʮ�U���{`�F�MEk^O6M�����Q�~}��D��g?K�V���dn�GA��P�	ڛ9 x�n<��T��@��>����ت,|�����&ƾ70�g���]�+���=�2�K�$��1���l%�M[�{\�0���� r�)��ťPǰK5d�?�7�A{�}���o��u0�G����D�*���I�@��YOy Hd8�(�� �Z�;6�yB���L,A -1sz�� ߓ�-�J5��uzڲ}ڙiU��<�_v�%�ѦX[�KD�����n&������Z@�}��O�_켾g*��r��!��I"`�]��$�b=�0��eO�������ߝN��l�&g=|0��bR�E�?K��V�}���PX�ci����5�,�y�������ê�:.�%DF����9z��լ¦�ef!���&\D�a2k��<��<����3[�����
���<h@�q�7t������q�F���%֊p�[F�E�=!�k�<|Dyn,
�\�38�/��h��^sP��1�qqjx.����y�8?ƍ��UT����I%v_�N3�)P�����EN���G	o�'�׈�s�Ǳl]��\�A��������\6Q�`w�g!�=AoE2��
��:�7�l��p�n���k z��*�J�����IYe��V���E���+ڷPK���� �`Լg�[�;��DM��������.�J�첦�os�?h}�`�a�6R������-GH"JaT�T���z��=��"��E�6�b.��Y�#����lߑ�s|�5�Q������%�W�y	��EU#��0�� e ��\��F��sDqB[�y��7��ZZ�d�s��v�!,:��kK"�����:곑=!'��2�&�;�%m@S����� N�i�Ӗ�A/2�X.��q9nL����q�k�1T� �!�+���\����N�˭п�$޾[ �-�-Ǫ����:E)K�k�}�cr��E�{y�s۶?Ɓ�����iE��fC=_>e�x)��s��oLY=PR7��#�c�'�Y�+�)cq�sK�%[g)r��j�4ؾg�}���\s���u7����_BRe>__w�PDE�8.H�\�Z�"-	x�|f�S A��u�0�5��
hخx%�Љo?Յ>�p��Qj��o�S�	���D��5Y;�|,ݑWE�[l!|оn,_.��&�?9������pC8o$�BK���:�E�FF71����U� @��$�(��:��1�US�r�t�f��kx��!쾨�|����+|�4���Ef� �+�H����#��k?�G|����!�,b|��ˎ����)s"��Y���#���C��G����*o�ws�f����ջƎ��8�'pL�(�`	MBOCbf�S���!J�yj�Ow��&�����b+��sOV�d�=���^R~����P�Q��+;�"uL�_yC�
��kW�0WYXD�x��z'���@����u�v����)6�J�u�)�<]�u#��%صhYy`#������0�<�2�΂����h.[�'����QoY���^��e�ӹ��dG��y���j�vh��o�U)2��
ՉT7>.�Y�r4n�Ks�L/j��m�t��mz�X�[�$߰��X��y���;�S蒫u�je)�kz����Ru�cj�	�-`1�h���*����`z�[9�£��4Fv�޸�9������R����ɰTo=��U�o�g��hyOnw�=z�9��;���xF5���db���V�e4�7��j�N�@��%��o�ä� Z�^�^ܭ�ᣏ�[k���.$��ގ�j����2�U3�-�%���»\�	t �C�J���{[Z@���;�BCXB}sl�*�릴?:��u���
5!��iCU��FӍ䗺��'���+��8��OԹm�I���c�{����ob'�.��]&����3ha��ه�=�QCa�05����-
`-��i_�S�h3	c��;ց�����Ntq�/^�}��\lR�����־*�\��DeLz.b��7���9�'CH������V�f�+�Jf�M >��6Jͳ��7�o�g���R��[*�>��r��t������?���u���+�����?�:mѭf��P�L�Y���&C��`ĚMׄ��C}|~����*�9/*�{�W�筈�^�����r֜{"ky�$=��Ö(X[R������y�v�n���\Ii��{���$!�`&Q��E`���#o&�п�lm��C[{]�o��6�t�7��&���=�]�`)-x�(�#�o[^��\�����*��C�kf���'֮�"��a�{��4�<��9^�����L���H��Xa����@��������LK��ʦ�F���W$I�3��yd���� ɷ�#�Z����)#RC�řv���5e")��kҵ��8���y]W�.��!�`p~k��ևLn0����� ��)
Ã'���~�D�_	n��S8D�V��}	&��y�'��!�TZ��?��Ө^�J��Ĺ�v���r©��I�2�[։ĺ�P�e����V��jIy��J��Q�"�+�yd�	{�O~����A=�
����z���ك^T0Bt��pUQB�mN��-i��͊�,8�5��N�-�)@<�73f�3��VЏ1?+D9��l=�H����'��+�Ѡ'T���O�C�fؽjA4�B��r@���x�������t����`"sMv�W�nŞgzrq����#&s���'�}�F�쾸qX�mC�M�� ��M�����W%L�*nN�Lu@�����l��e�n�@o��pk�=��#�����~������
����G��*�v�����(��}�DV-]�����2l��P���j&���Ӧ��"�=�
�R��$����[%jN�������O�Ua�9�Cx�zY6� j<�v�4�$�[B �ɲ�x��o/���XG�ʽl�|�>i��V*��{�bG�܀?I�cxSv�칃F��:�G�
����m
�n֠6|��&!QYY�Ѥ0�P�:���k�q	�LE�:U0�@�����W�7�C+^+b'5�m�M�;P��U�P�/\A2��ۭ�3g7�(��P^���u�RF�X�+k�V��L��N����:�΄���_�:�	���T������vS�|���W�L%�N�����Q�/����g6�bw;y2��z�'(�3"Ɠ�:^�%���0������X<J��H�JS��9��l��d�f���N�I���	�KO�y�r$�����&��1�T�h�|���i@L�n�D><����)�H"Z���D!�.5�=�b�Xv$ b�N�G��?M�Al����fa��"8��[����A�2��s"��K��)�$�¼D�/�f|%x�*���&J���!:�,3���0H*aoiʱ%+�͘X �%\[��V	2�_cI�{��%~�wwH��Ob��
D���c�)�Zf�==�Y0��}����2�&�5x�=7X�z�����U�S�ho�����+ ߂J�� ��-�@���r9ꜜ~-ǳ���S���I}��<��x�(��닼5�Eʇ�d��}݋�[�P�J�s+�����ӷ,(�+�;�<o�$���I��<�QP��O�!� �/EvT��2E��?���,�+�菅=�?���%�H��w�LV���v�C�՘��JI���v����Wmz~^�*K�ej@id�U�łjX��9y1�5���W�����=��h	y)[n���Q K���h(���9|�o��כA5}�b�1��7����"-�k��˥�IY9RO��xM[�� �ڭ�A������g_&�MtT�y-��>���.��V��'��J;IB�h@��A��)���B3a9��%��e]^�1N�U��ف��i�z��stj��~D�%�{vޭ� �f?vݣ����e~ ��:�X@;��ڈ���D�ݶ���ɫl�z��D-�\��$���|��H��$�x���3A� �5ᾍԧ	���+%�HX�m�C	�riy�o{p��K�pV�!���>��i4��q��>�w�Do*�2�s"S6ݟ���-�/��˴��!��Ef�����+�� ���*�໠jqԠʉZ��s�7��7d;4�Z��$���Y���ۼ*#w��A<řތ�GP=��8	")�C��b��B��K?�)9�������\Ӓ|�3Aa�\	�c_j��3���� �]?�	�����NIm'��JQ���
�����Ȑ�
䶵�5/���7��U~������a��O_YNTI�{Q "��[	����f^q�f�D��`-Vx�]ǡ�߭��)��M�g��t�'�	��f���	��p�a�����lڥ�`�Q�-)���)�כAp�Gg��h#�W�g� �K>��Y~Ƌ�o
w�ꬹו�[�а%�U�fA���@N�9O��tH%䉵��Ȯ�*�V]֌�y��t>���5�w�]CY��>P?��cD�a\p�sS��z�D�T�b&\�R��	B�]��vBp1���})U�&`��I0^��B�g�
��B��X��f�����I�*����ʞtQ�9ܶ�b�$�qU�΋�n�?���o�����χ����x�M ����)QKK���2ݘq����*3RVZ����[�m����r�63���� Ou�Ƭ1��k���Sa�x<��w��1���s��Y�����������b�_xSf�O��v	I���^�uv�E(�c]EN��u��y���^�謄Ń���2�蒩!�ѽ�������O�~v����T�w��/�O����bvA�C���<H�8��d�/U���u}��9�{��bB�7q�ֽ�L�h$��)���Q(%��ʍm���/����5�l�}-(�f��Dޣ�_���c('on|r+/qy�.=s�Ɇ�w
�4ڨ��,�u9��ޫu���>��#�!!~kG-��==�Ő%����b	�� ���xU��)�l 3NJ�7��-|�2�9�V
m�i��ۊ�9�O�xH�_uZ�����H#�R����{���m��+j�͌D�{�bA��`i��� Uּ�E����r�>+CP�}�w��T�X�KDG�Vd�l� $��[����L�S�Ւ�L�P0�����
���\�	�S���Q7�bp]R��,��cn�k]�R�	x	%��
��x�f�i}�� ��fhr'���b��{��>VQ���D�Q�qOV���ٖ�A��Oao�̶�:"�;�Dt�?�16�|+�v��؂��e��LL&j�t"�K���ڞn�E.�� p����<0�6ɚ�3a�!|=�mY�TP�,�͋����R
#����Llg?v���c�;�j�S�G.:����:yne~C����ő��G�O�d�6�� .���NOzz��a��E�_��vm����ҍ5#y~&�
�w U�8�:4>0��1���}Ły����5d�D�����UYH�J�����Av��-Ɔ+�	}eV��3}*�e^��|Uǖ49'�zP�*������9=&ï$�GC�[k]"j�3��@�HS�=�-����06"0�p�}�o'F�[��<j�eg9E��=���8��C�Ԇ�I��
������xӶ"zFY�Nes���,3��&�KE�ПZ�3�g왞־����$%���^�J)l����[����Oq�¥~\~�C&���v7-E�}��NA"(���'�T}X�k�?]W�$�{��C���Tp��X�&�Vx7ar�?��WR�(�-�j�I�k��rii�����_,��ť�̡���
k~2W�h��,k�E@Y�N��nx����G��=�\f�WK�o#]0�>Ĩ�h5�Ow2�j����v�pnW#�-�6o"5^��R�
����9+a{���C�`&,��,�Dd�N-Y��{�B��+ީ@��V��hTl,�U��eW�M4v4.��~I��T�>{�ΰCNPC c5�#�sf���.����6�d�N|�RWCOͿ���ς�I���a��l�I�O��J�:�y�݋�4��b	�=��R���}򩾹��֢켨/�tJk������mH�K:T��F۵¿�
2��x"�l�k�o�5{��]�j�îE�^'T��e>f�P��_c�u':&��ܧ�Ew���8��]�֝�
3�PO���frJ��D�W�(Ϫ�8o���Ije5�H�QN[0o0&ײ �Z���n�O��i�[�c��_y�/�Sr��]5��v�����_��nʘy�X�e��͂���	�<ɗ�].qa���{��?�^*��CE%�^<4{(��5~���J�z�9����nPi�
��PGs�P����O�"�$��;)���A��.,�{�����9(�^��\X�]Q����'Q��
�􂬄@#��kM�{���bd.8j�"��r���/=iI�SfPMpI�%�:׽��Jb��-NSf��Z ��¤w׸�	�����wl�Vt}3kN����ڴ2�V_�X�P�er����9ٯ���"}��%[Q�Y.2*���bf>L��4W+��v�Qں͖_�l�*�?�&���x�%^5�����Sf���+�@���� �/Q1�J]�%����l�r�/3�A|�c�R���uK.
�V2ߨ|�lHa}�6eԱ�.ܶ_���t��'��jl1��H;S|�	��������I�RHY��$�m�2Ii;Kv?��K�Pb�e��1fe�P�{�p�!�Q1γ����X��^ ���vJm��s<F♤��N�=g͓�eɜ������E�~����W?��5gk���ԅ��/lY�?���t���M�ck��V
�L,�/~WƱ�=}�&�cs�Zd5&�8v����7%A/� +D8�<�� ��
V��@��E�i:���R*�����-�v=��+9Z��������
�nZh�΂�X��$_�U�Cn�M�,B�' ���{	�oϓeʅ� l��־�I1TS������2Ѥ2�׮�8Y��W�,�Y��a�AѾ�nJ���sIc!ab[k��Z�`�a
�zg��+��%���u,��8q�o�b�K��Y׿�ܼ@�Y�4���40�*-��(.����7j@B���� �.*��ջ��� �L����{��VKf�������`bb�bo��O��C-z2XB�o_y6ߞg�m���02L��0Z1-;FO���������]'
IFw1E��U6��"�#�V�9���|_p�0U{%ʼ#�����T��s\���Nc�� 8��:;�5�M1ϼ9z'�L�S���K��1��o�/��c\�;�M�b�7Ǟ�2���<�c'�"�J�DX��`N��$�t�5?),߬Zp#4U��d5.=~A��˖��^1�0y;����v�|`�y�FJ�s���e���Հ�6,�:�����,&21)�!�Xʑ�ፀ�r���N�+͸{ࢎ�/�\ #_U���*b�o���K����8�ݥV�g=���4�X�9�F<�8ڟ�xFu�f�3b���ʕ&zC�iB��h=�`� �:oz����;�r/I���E�>�pir�U3�l,��^f���|$a��yOn��l�!�7[��'�n��3�K~�$B*�*�A�y%�6ۭ������Ә1�`O��j'K�0^�V˚z:4rDԊ��p�Ŀ��:4��mH�#��W"SϩU�ϟ/ӕ�3׻S��TQ���rFa�(LM�����ϩ�itS���jm���˱��?Uq��@'&�r�������]�y|�����^���t���K(�d�8��j#�#XL�[�]��GRU�
 Y�l�E�uc� Oq?hdϨi�9��?.�q�/����&���a��n�ة�5X�V��V)��& $�k����͠�nWMu�(ɂUx�L_���>�͍��D��ע��f'�$cmX&���Y�ĳh޷�~i�c} ����x:@W�s^���܈J����
�ϕ�ZX�mls̐hUE����k��>�>����~�i|�u���k��%��VM���4�2�>^؇��ɰmm �fMR�*��"��۲:�U�%զw�FV�O��,�����ꮢX�2	O�_k�����Oæ���E���0�))Rt���Y�ɖVN�|3�h���&{�B�1dp)�f%S��&���9���G��,�e�m����W͢�����D�$�Y��l��z��hRȴ�����!��ŅBHu�4t�k�ޚ�z�\��t��#��fUy���o7WH�T����,���F�.H��A���'(�*+ڃː��}tȶ����6���3���]��۝��~^=��a�q�o!�en}�s�A��m���p���T��yFI#�і6/��7(茣���z�:������Bo�+,5�E8�{��J�Yr�1�5�fI�8��4��\́�[4�㹲S�8�����~���}LB$���i��*���H|QP����D�Q߆�_/��d膕��Z�a�����ƭ]#�mK�)�Ej�<����t�C0q���
�Y��]JS|���O�ۧ��nA��M����ڟ��������l��og���Y�d��:��&ȵ"���D7�}��*��fߧ[5���Ή������ڸ��G�A������I��ƽ �A�s����f��ޗ�p���y��o�%����u/yˇ�ZXeºׯ�3�A]��WP�����겐�3��/x�Wd�C}� �9�2R������]�#j/
��>\����	��u	�)�����Hā��1�t�_�N����u�?�RT`	3#%��XH%O��$G���ms���ޮ�]dQ{�G�s��;E����%���ㇰz�P:�G:��mr��[��2���h�b��N���>x�i�?��|�zx?lS���7=<�cP5ofiʸ������$ },��)�}B�r�0�GD��Q=s�� ��}&�c��`Z)�[S��؊� 2u�܉��%'��`�Q^>>��I��9D��U�@�zRɨ�M,#��cZ}~���5�BN%��e/�X��6�7����<���N�6���\c����jQ鐈�I�.�^�:߹�"�ǧ�>�D�yXM�t���uK�h��<*���{��kz)�M���X~<�����eX�����/v[����HJ�oSV��^y��Ò4.Eł����0蓥'����/In^�!����[Uz���!��F~�$kZP���ձ��P[4�V��F��w�q6aڤ�#�9�����&dv��ڦZ��$:�?��+k%�ƅ�ԾʟBbI����D|��KZ�KH�֬A7>������+Q'5R��p�G��P�;�	�K���K/�?�x�#�7�*�� yC�=Y�H
��+Tݺ#�xX�k�8y�#���B�#'Q�Y#��Qn��01��x����	J�}���5 ��bG�l�Ru�>��N����7��4�5S@cM�T�� ��$���n5v�c����_������N�fh ��Q�.b-��'����� ]�ǌ|q��if`RQ���A��1�b�W�'���j��nj:�6>�OL�: %'O����Տ@���t�g�j��FLq��(����v��ꄪV�=!�$`� �/�&��]eL����&�(��$b�{EW��ac_��)z��Cu�9e'ɲ��8Q�#b���"�/�h�������f��Vj�ɦ,��VD?�yr�U��z1v�/�4ʘ��_�;B编8�fe�sH2��m2k/>�����lz��5�:�d8ʺj�Ev��H�/��h���dzS�mD�h��g�%��QN�6r�� 	OXH�2'�{�arl.�&$S>��n�^_@p� �(Y�}>�}[T#/�[�T7�,� )�t*ѡϫ|I�r�Ȋf��鼞W�<���~��F�f�s�M	�y�ύI�m�p��!~�YD�ߝӢ����1(�((�'����-�\ǻ��B��A�5]4��b�9���T�N���IR�3�0i�g��wr�i�\��=�s	��I�-�"� s8X�2����w��Ѕh�O�T�m^�4��ۊ�"��	���#j^e�+�K�C�^���Ĺʳ��[�6�P��l�x�P��!�I-��p�1��Ӑ2g�$[���ǌ?4���'}���޸��)���aˀϨ���WW�ST�J��j���2X� ��8^MA$�s������`�^J�B�[9���-=�Y�8h���2��_8����������,���^��.Mׄ��0��^Xá̔�
�o�C��5J�{s4�����j���'yƐ�R$�S�$���[r�	�%J�3ؒ�Ts$T��{�`�J�-ЍM�L�>��n|[�(5zZYD�^��]m�F���rU����˯SI�Yf�j���	~�����ܷ'"����\]�������5*//��F,��q�yU��6���j}M�@��.�'�}�ʺj9WԨc��sw����u9�c�����%��8��K�e�;�����Sk�	�F�KJ�#r���X���1���b��dD��_����M���SDp�8�o"�-��~�m�uh|C��������Zr�9��8|���r�B��'��S{a��Nv�J�H8��#�yRL�-Ɇ�~(&|Mu?0�w}�iB��=�#��`m���~�~j�G��fc%O���m�O��4h@x,��d�`�8������E�q	a�>*H�~>[<},0@������v.��G�e�K����a>�8ҽ�r�Ƹ����jC_���s�D�E���H=1J�sga~����(&�ߜq0d�����������|�?qk�0�Y�#�H�<���C�o𺶟����s�&���PO���J@�I89#���!W� P���r���A/kA{�u��"[���)��f�8��{� 2����cP������|��Q�1���-l[�Rv��\�C�/��&���r	H!�@
��4�<6����H!X�O��X��^�zY�㷤��&�����!?���"�W_�Z��>Ei��z�D����q�N�h�[�~��m1$�����8�m�p����=�m���TA���:�oV�Ћ�O����\����lg���I#%��Q{�ڬE@ � �V_�6PSP��`H��d�]���{8�Z5V0O�oa��&�U��\�\�Z����c�Iata��ҧ�H%ta[�&�x\��aScN� ?�m�u���+�!�-U(Ë��	�wШ�g�}^�&���u:�KG�>'�zʆݬ�:dj��@ �V�Q��n��=Ӣ�?Oc֜#a�����s�1��^Yx���k���m�l����%Z8��k��q[v�T2H/R/
q�8��x���}R(�k ����Yp8�^��V*��#�����K��'L�����j�L��.�l!TK�8r�%$�v�F�Ch`V�C㊻;YN�iZ�F��`F�zB�TKi��bK	h�i��R�9G�i�E��7� �SY�qz���W��-�	�X�ۣ�����-�&:bר�5͈�<t� ������|J����:�aK�k�r�z�#zK�%:&X#v����տ4���/zڅɟ\m�7S��ytj;�4��I�$+�[������HT�}�fB��B������%�~Gi�w��@P?0�v�v����_L��~e����G-�,M��y��6���:53�<�X���<uя$AW,�z��(G/h	Ynli�=j@�M��	W�i=Iކ8���P6����6�j=�܆\�52h�F�؋1ߕ��T�`"����+�W��\�J�FX*��+��� ���K��e����?��h��S���eX��>&��:�����a��[�4sEqT�S�1����f�����ɭ��$ئ�G����X"��:�=�Z1��8�װU�fg���J�Y�Շ¯�0�v�/k�ªZB:��r�U�b���"<IS�=ZҍJ�I"B��ՙ:҆�FCK��![�L��AT���xq$������n�A7{���s\,^����|�i2R~�{����Ǖ7���$`�5�0�j�A80ݔ)��	k� ~YSP�	�(|߭���}�5����D��f-��*��r�R�R8b51s:���FO���91	��٘�?fh�i��rd���DZɁ$ۀ '?yl�eƥ8�ȹӧ�E�2����|d/+���a*����6_�8���:&�f�;jN��b��PN�Ota�i�.�׻" z�[�odiTx�U���b�,s�l6�~ZH"�g���9�*�	(�b������z�1Si�$�?l�_w�*�)2K��l��8�/8��h}���`�z��/�'t���fFi
p���A.�"7���>4Z���ޙ��?߰����:�݄W�~�`_5Z����R�TrH�?�aZ��@"U16�i�&��O���@�jn(�l���[J���پ�q��ٴRD�	�1ęG��M��;�M��)�Q�G��WI������N������[>z.��1!��3�MNH<je�H`C[����{\�iiQr�H��b'3j#~�99%��)�p�
��Vu�[\���[W4��� ����T(���4��7ΕO�d�٢��!r�	�ԉ����^��R,��F��0��^1�(��|*C݌nʘ��W"~�������k�v�w�ǵ���E����}uP�L5v8��R=H�!k��h75���,h7�8Hk���5���t�s�~	 �𱬙��t�,���?@#rUr ���0/i&��ı"�kX}�����7�]�@�������p~nZ^.t�|D�$��.�'4=�����)60�&(j+~f7,�1�p��*����Ëo��Z�NdR��?���������l��?��<HT�ַ2������H� ��:������p�$�p��(�΁q��T�2YVH'�Ǘe�^?(�0�κjxzu��Pln�����y=xC�����r\��"ܵ����U2���O�9��������d`� �Y�<��g�i�>�5�O)�J���a��p��x��SNxh^h��r[�	H�2Y��Oo��Du�!>!(]��%�M!# ���5ST��tX%CH���h���>bs\��M��Wf�����|drx���G&�h-�>z�@W n��g��o�>���l�*�I�탍���R�3��]�l�D/�q�}�FC@4i�M�(CȰ���1,ɜö�jNI�ZF&NW��^��ņ���0��M-�e�ٯk�����ߎ��%(�S�1k��6K�9�b��'�FOR�bn��0X�a�	t�p��-܄������_u���u�$аY�
f�tR�-{|��!��TL�+[��1풤��v)�d.Zص�����'Û.���Z�X	�j�y�%r�Y�;
yدGpuS]�SA/_�����0Q�N¸$̯v8�=���`�u�B)K�qbm�ot�mL=,���R��+@�-[�@��R~� ��n��5d��S�(���I�ʧ�)�B��e �#��g�v��Fu�宆yx���������3�G�#S�3������/���@���*�!��[ ������1t�ԅM���\�d;��1�wM�`�ujCBnr�����}�q���.�D[�S��l�����U�۶��C��ޯ���܌��T�2Ffđ������RJ[(� U4���SoFS�4u�k��HU���C��C��k�q�4Uco����W�确�];z��eL�8祫4�p]��o��ݭع�͸����S��ƪ&C>�Nn�όu��ޝ7SJ[�rJ�._s#~�K�%E��y�!�y(��G,�:����zhs{屺00$��>~
����k*�޷@��a��mv/�#g��_}������;g�&����x�Ī�t%z�59�q6]������Yå�"���gSt����*�)wY2��"���c�)�v�ӷZ��tz3n��8�3�,�|ʵ\�IsOd�C�/	l󈸶8>�G⹍LWՍ�>D�ٕ��&~�T)�	�Q<0�;�)q;��(H��I��F��d��U�$��j6,�רc>��K�S�?��4۔��*��J�|>��2n��)ƥ�U����)�	���,���✇@���$M����?<l[ǎaas6��祎W������
0ZE�[�`)�>���:��S+�ٵ��j��,S��Ν�-�[�dW������B��PߚL4�SIɼ��P�tNE���*��RA��>S�s��$��PDϹ<��\W�ޅ���t8��`���(��_	q�
�I�S������%"�fe�A�`���b?֤�QT�Gy0o���eۭ[еVb�cI�x��H7,��2�Ʉ����X z�/?��Vܙ%t���P�Ѕ� -��/�I�,��;>nI��LŶ�P"��j����Ԑ�5���d���h��=Y��>��� ҕyF�/�b7���]o�� ]�"�Hl0�P���%�h�7�z��s�K���x��U��u�u����J=;��ё+�yS�$��ed��Ky�����6����fx����c�3� u��n��F��M,�9em 
�KkH89L�?*�L��l�
@i̲P�!�j���eJq�^�O;����&���NYR���l��8���%�%v��� �}��i�,��e[,����Z�I��p�YR�!��"�"���1����5��w |����g!�!wN�\���~X�	'�g �nr컙�1Ja$�]��k�De�b�κmCq��T	3�Ro���V����n��\��>"��`�������J/_.y�L��sDl-K��/퇯�S��5�����/�������[z����I�Y��2�r����s��6��I�$�,����]cb�fdc��	�^1T��)yDT�lk�x2mq67��B�����Gן]�0���M((�%�C �\���}�a����5�U�ת�:8�[y�c� Y��CK�]@0J-WkC��s��_o��#�>)pzc����{�A r8� w޺ ����W!�	�i�@���>��VwQ��k��Q����	�Q'�c�)Ms� ˄-s��s�n���u����\���A,����yh��H��l���[gXfOz�fN��q����B0�<��k� �-��ۅ���()�2�Ť-\?_Ǡ[��N�XB��R�0�|�DG���|�>�h�\؟��ku����)a��Q=�
�֮>̘S�T�7e��AF�d�O��R�� �̷�f���A�hK���6)4z��yV�0ߠ%�C�{F5k}���b<?R5]�2���6�n�m��ԎD*ߊB��|�O*�+�]�և'��R�����IU�R3՟��w��|�^�
���s�VWiqAX
�ݔPJKNi�	�O:(�x-6JD�_s�r� ��	�M�����=���"	�ɍ�G���Dl��L���݊��C��N^c�14����2����>�����Ĩ���B��a�M���~��;E��ְ;恆�k�;4����IvrHqDۋ_MZ���|@�Ї�klf�V���D4��u���".'R�zT+���#�n�/��'�D�]o�[]��x�*ɐ�昚,�$%���f��MO�u<����x��[Ώ�0.$�!er�j?i�I^�^��Qy�b� $�A�U!������dV!fe;5:���rή�m-�f{͠)��gU�a]R�w�������]���4߹��GRB����!� �*e%��*�F]\��/w�=M��϶���9k�T��P,*\}w�(�ٙ��S�m)���*�	�s��;&ȐU��W:�`���K.�B�*�Sf���%�*�,�G����mvm���F[���]�
6���d���\��fj��z�%�D7�I*�֍�}���������x�X��S� ���v,6T}��9-7 �5w���V8�7��h��ʅ����e��%vv��7�jem1Mkw}}LG,��>�}	��j+�MQ�ز^����$0��mՓJUE�]��N|�}v�.4y؏�Y/��9�/�+)�@B$�FШF��u/r������#L������g�V`>��]��1I�0i5%�����}�w�GHJ�F4�^�ǳί��;q�Pw39E�e1O��L��eB����ɵ0�3�q�
�U��KxShV��@!�oU�d�swy9_|9�CK�^�j�3�n���j���29�S{���M��zz��U�>�_iԍ�\�&���,ޠ����C��FiMN����SЖ�AL�tㄌ=��%a�>�oNR2��FQ~��:43kIg�1vc�Y�]Z�(��I+O��\���|���+�{I���3�p>d��Yɶ�Ŝ*���2�G7e��Ə��$K������x����ک��7�/�谣�|�:H��V[�/Qڢ�G�B�D�Sj�$.1�|�O�����%)�������s7�L�Ubo)���QJ��[�gD^]-�p�>%F��<�.I��@�����S�Y�	�:�e/�6'^4�W�.i��`��Mam	֌O��Y"Լ���:�:9�_)F��(��,� ��ӱ�1�X�G�҇p7=O�ąd�{f�,����I)6)�qT�"P��b{]���3�*���?��[�n�NN�J�2h������F
p�J]���;������f�O�1��H�+���./���5�G5�C�z5	�z�3Lq�I4/!����CS��B�ת��@\THZ�
��RM���<�!���ܒ��y����)7�>��H�^����ٚ ],%X�P�e"��HZM�j;�k�\Ep��Ұ�,3�9�܀w�T܀s�1{��HC�l���i `�d�tn�{�7� +�c��Ğ�ܐQ�o��ғZ'��HrM��셔����P�;cf���\}���Fݗrc�Xwj�f+�b���a����v��!X��KA�;Ϧ�{�(�F�Y��Q�Eդ��:��y�Ql
����������܏��ӕG�GA��	��k��ƕ�U�0�=�E7���%�ඊ~A�NdlT�7��wa�n�ݢ?��]": M�Y���V~|`��ɒ\^���!J��tٕg�4���|ͱ�~�VB���jƝs�O���	:>��k���O׹��!���6�yR�5F�,����yT� ���0 �k�	EU�z��
��'#7��u/t��l�o����Ϳ7���˶7AE��ͮ�E�`�����2��1��b>������٤1�78��i����/0g�Ƶ�K�3��rma(a�y�ewUC�)Vyb�:��AҡnK��o'���2��u+9��U����Ҵ<���t��Q+��Rqm�]�uOg:�x$�V�6-�Vy�G��:I�vW��!���6�}�|�`C���r���6_\�/�@x�C?G[���W�E��Kf��z0^Y�э�@lȪT[CGcT�1ر0���}R�e@zs�_3?<?[�B_� ېGn46h��,-V��[�|�M����ayw)3Vҁ/&�;�^mi6���Q%����� T��}Z-S�ۉ�E�æĠ	5�	-b%�,r]6u��#�5S(���h^޷��H���8��%D?~���k�Z�Kh/��7B����r�Q������C��o"�J�౓�)<~��L1I `�_�ְ4�6,LB9��d�*��CjR[k�Z`f�7�C}�7M����@�\$k).��ߞ� �����&lL���:\E�zS?.o�I�0t�*�n��>5!f������:1�-������ @	�!2|��j:��}�nW��$G� !�x��!�*�C�|��
h�f��~�<�T�-�i��uE���
8�9�d~�mu�v�(���	�c��;_�٢���U]�����6 A�����K'���cܣ��j4\���&E�fB���|X���Pj.�}�h�'���ic��TmYa'�MO_	�l�(ֆ�ZB����L)�"����oݫ�P�H�tk��GV�ZG�8�+�LJ�99wᲤzF��(/��u�������%S%���Ҽ��C�� x�ql[�dCD=����$m�꘵Ym��њH�Jn�����SCj����1�@��,��9��z냄���k4F��+."J6)��n㪆���$����wNp���+��p�[���ά��4���?Q�wdU�^ra0��S�^e�QeQ�;��hF�2��B8��A�!EU@ݱ������](H���	�$�_���m����O�2%#�G���P��
�|�%�`pq ̗nq#�:QP�̔m�\�r�&�xj��-�=ؑ�^_�)3�f|�� ��)��
�X�,"a�����H��,F�J�'��LW���'a�͸zI��LDuT��9z�Y�g=X�`p9��	�1Q�u_����a>o�Y�6d9�f{��D��t�E!����0�3��������&2^!��  N���j�W$1X�#��B�#HU݆���$�W�&K-��B�<u��k���mF���Ù""/���z��/	�u޼�Fc>ՉzW�cM�U�In�� ���]+��q�Ф���j��^��Ȟ�@}��N&�Z�X`ǝ�c>��i������:0�¬��B�0�n0�@������.�.�N���j�������|�$�K=/��?�Ċ���_UݓX����Ԩ_]%�ᷭ$'�@�|���M�4sE��K��pغ{Ҕ� �P�{�6�� ��
�b$2~�?��0*?T)e?��V"�+��R��T,>b�gs?,G���;a1u�&.�V/6���T�M4��3�v�ȫ��5<B�m o�%�L�{�o_/�͆���^�1�qM^�7tU��5��`�}��w5�C�@V��xjW������Kz|+��8�A��Ɠn�t�`�_�����MڮA�~z5?	�f���ݢ3*�JXě��\7�gm;t�湷Zh��[%UB��|�������~��������v��k8����5�3�I1�o���w�25ѱ&�i>�+-"��v��)Kw������K��(n�[�Ԃ�W�B��+���z���'�?ڣ��A��mG8�EP����-�����p-��[U��YT#���	E�U�ع���w�7��d�m*�\f���A�.�xo�&�	����p����A���ڬ�XҨo�.�~:�a��>�Nr��x���@K�x�}�ej��(g׾�oZ�:���m+[*��&��;��
��������z{�N��Ú%?|��i���T�LX��hK�W�GJ�Q��qQ<&�*�X5��V`S��X�8�",�|�k� 9F9�r~ý�Bj<'�;��>�"�v��������|`ͮR�qrhn8߫���~R�Yz_Ɩ7ǹ�q*Ȟ�8�L~��[Í�-_���`<�U�>���k+�j>nn������l��P )�a�����F�8xN!�P"�gvǨP6�[7�2[��MT6߲�J�?$�{�Ue>���J�<1���E��`֭���Ϸ��䅪���:� �Ҷ���C'�(�f��P_�"�!�c��a]lՖ�DJy�a5�~��.�m�Q=**���hD�hZ@@����)�2'X&C*10������7�V6�%D� [K�{Ғ8�r��v�����?���?A�qp���X��6�O�(?i���O�ql���9��^@`I�YJ�O�,�UfаP���MPb��s�E�M�uLyz���-��s鍪�B��߫b'g7��0�_f �'x�V�8�����Bx��깳����]��_�J�#�̓�;�#�%,_	�P��_�7��o�h�����`q�� ֒6>�E��|Ae��?�RPqZ��C�z��-gc%]d����X-��A������,�a�g�r҉�p��F}4��Ŏ0����,���u ��$����K�BɬM��³(Ya��g��9���|��[a���O�Jr��i�j51cq��LaT�\%��r�m}�r�b�|���`cԻMP�o�`��M�v��x��o�mY/�J$����֏;�L��U�#�2�qp3�����|�k���$>�uav����I�*��1��3:h��?��f��
��u�`G����&\Q��-�*��{�<sa��R����l%�:�de�j�4�����l�+D��8�*�?�\7+b�
� }
��0"��V+�$�4�������5��^~���f�x	�N�,��V�jVIͯ�	���=As@{�d�A=�]���Vֳ��
����.���k�#@����=���d�7�K2���-{�θFB"h}�<o���z�rM��֪:v۫�s'�oYQ�?��Ua�vEL<�s1B���-�9��=�C�6� �&��Cb��J!��G�+��0i\L5­�2HZ-��a�k`�Rn�����DvG�w-.����1��e��G_����A4�3l�nY�FJ�U8>Wb6%DG�p��rq#x�MgӒ�/%N]	�V�p��@~@_�&��/0�>'n�ǻ����ɚM
Έ)0`�v�s_���P��#�V I��R���DCz�^,��>E9-����Xv��'N�*�dq%S��Cп�s�gf���ddaQ@�x6�I�F�
K����qi��	�
./�,�uqO%�Wp|c�����)�OM�$0�]���)D�s���^˫L+-&�%���R�#��V�+���:�j�����F"�+2D�B�方�������UXL��?3�{zC�F�2Q��l�ԫ��V��6t1�]T­������ f<n6��?
fS��c�	E&�Z<����Evr]
�>Y�O��E�TE6�Gq�jB�QC���A"CC:
Y@�d�L<�5�߃��A_�c�	
�>g��-�Wsn1֜b��/.O��c��q��إ���8}P��
y�����[��F��c[̲6)2P�3�N)F���ޖ���YG�f��峜�nD��S�u!��)g���X}�c�t�N�����h�)$5���[y �~i6t��f�3SgB��3��ZN��E�ϥ��
��4p{�
@���ݛ.?�֝��_qR�U��e�D�� #Xt0�tZ%oV�b���Pnm��.����Ht.K�c���c����h:oV�_5�e]6�����4��z2iN��tHL{K~��٣Ԁ�	 vg�?Q���n�I*r
Lw�f��Ts]���S�4¾�L��7��#	���4�\���+�ug%t�4�gK�یN|�O��t�G=.h�g�+ LDVc���A"�V��z���- ��gs��l��$� ���~��!ө���������X7�^�v��Q��=� ��/t����s�>��[����0��d����6=2�S�`T�h��H/,`݋��-S-H�;C"B�OW����r[	V���^���$g��ζ�lי^M���u���?诗oMi��kF�n�c���Ԏ���)��H�?ݧR��J�s%#ԓ���	��E���'J޲�5��AM��>@�+�O����1��L惸�`�H�v,%� ���>A7}p֚���ATÌ	Ơ0i�4�c�7 �(�6E�M������=�H�k��+��I�	���m!�{{a��Z��A�,��i����c-�6���z�U�C�����V��F�c��7��IG��<�"hKV=�1=t�}��=i��8������Ob"��9*�̄�Nwr�b�6F������%c��j�ia��*y����X��&0������yU�-G�����K~�����{�0h����zi��	���vy��t�?�_&���9�X_�֥Ǖ�y.ɾc(RQ��/���$N4G�ܞ�&�����GT�4ȳ4]Ej7^�Z����g�0 �`(?��������e��F��D��m79��c�d��*�]m"b܆�A�1�B@���`4'��0a��U��k� �e�@�����D������@���꠼��\\�O�W�HQY:����B#
�� �ko\���>���A��(��%���C�HE��4{��%�v�:�+ `P�?\�S����>eT��p�/2�<8�2��t	��a|d���I+���P��+��9��_�mT&���d߉y��w-o�M��A��%�J��S��Y���$R,����^���$S�� $,��@��!�T ���d� ��`����舜�j�O{«h��ΠPv�ի�v���g������ ��|�,h@_g��H�*�O-��حŰ�[zDL7���7��K�i������j��JV�t�gcrҤ��7�����d W܉
��Ak��1��b9���>M���Kq'�������ͨ4b�'��fk�J=���d�i;��'�u��~��|s���	+�+��X���o�g�a�P�ݻE���@�`	L�3a�&J
txQ���?�R�i)�_=9z����{�A��K���Ļ�0���Vvɂ��엮Ո�*�8��9�WɓXV�!��fy�RH�˪�YN�� �1�`��Ce���d�6oBb 7�E%1{���S �չ��vg��DT�v��`/�'�;�	n�,��֋�'J�@�\l�
��Zw�[�U7"19��lSbSn��Q����(\����Rj~���	ǣz���* ����	�`>xde�rBY�SYK��yk�s�`=�����k�Q-{�	�bJ�����3��kW3���#��AJ#���8��y5}t��8Uys���> ��/6�W������_����aq����ʹx�����~�o{g�|| E����(U�$�R�&�l�M�?]?�g�����ԫ������W��2�K��B�R�,�Y��NގYY��sK%�$
)�E�_\%8�6� w����Pn6�8����ZD�~*��@{�~��9�,���R��֑Y6�����O�}�t4R�v��t+@���rf���`��/��[�-ã���y�[�P�;�Q�&��m����r6����|���NA��|�fф���D�)�có��P�"z�.�-���"<�]i7���r�Fn�H�Y���<o�5<}���X�!DD�\i���׸���r�A���`/�`�H:i�T�(+1��kvE��ܽ��?��y>�,��vg��E+�g����-k�P�4�Q��t��;�m��^�0{)A@�z,���6�8����y�s�U}����qĶ� E�S�S�;K�f������l��b���������@ ��3r�#��Ή����V�<?�9��`J������T�p����׈H.�䤐�V�܃Rv ����B�֛Ыa^@��U�4��l/;�l�9��!vrO����}��]i8z������y���0���[k(�s��ϭ@��%�{�?2�Z�rJq/.�Lk��K5yB;��@F��@�Z����>G
g�yINΙ �aY����S�ګ�B؞�8d�W���O��F~.�7�	`oH#_V�A�o�U�`�EHd�^���.���2��x$���^F�)�=�u����RڦjV�uo �O�
`�c6A����o�}8Q^��!��A����*�D�T%�B|>AX6ls0�x؄�y���]H���+m��◔�{�R��@���.��3���x:�����5�s���a���x��p#sF�`}�[<[�[� �̳3�t������w�Ց� V�fs3w��pl���^�(��+}2��f;:~�)[rbn���\��V'�C`sHz���#OnFwl�O�N�����:�Xx���7#�_bo[g��@�dYL���=�v��8u¿�g>���C?�7}BUNXB�# �B�2
$���T�Zy3��k����:g#�����f�=�����D,��Z��/��aM�jT�_()Ԑ��dnm�KOݲLԅ��\H.��ZiaS�Z�1O��z�!�s��"1�ň�x��C��)fek���t��}Q��uZv�c~
u��c��u���0<B�g<��I�"��O�D������ؘ՜�r�p {G����Λt Jǭ��2�Y�q�� �H<�<��؉����w�0��_�;�v_��� 	q����$J�"/��������'l���mu�S!�u�l��C䯊>S��2O���%��j5��sg��vTUM��L��-�4�EI8�
�m�-�	b0bxA�D>��B��E�9�G�W��u|C��Ϗ`���["����uMoQwR2�h�024���i�>�?������Sã�d���4���؃��z�<����3P��nD��R��T�Ԁ�2`����.�A�>��,c6�sajy��\�؊�|��D=[��WbZIC�;����>d����<�M`3T�/T�e^�i�y�a��
�c���SB�>�j\���L���6e�C&���b�@zy�hzG#�ѝ�-�٦�b�a8�X�D���-�ȉ��T��TK	O��Wj��/{:0)ǈ�?��zI(>�&s�­.�Ӻ���Q`���VO���r$��L�&c����\ͳ���'�ϲ���'���r�f�7�L������H�g�m���A���r�&Q�ĳ���/�g����1�Ny'y���Cƻ�pa�\���M�UR��\8��<�W�	��br'��Q:�@]ZԦK�'���J�l���FZ��t�R�o�(�b���6���wF��ƵNV�]�N�{V�d�!к8#.̩���(L�D����*�������Y\��ө E��I7��Ѹpx2�Q�L�f#U-4��:"�Eo�ϒ�q�2���u�
[ۼ��I��nU��y9J���^�i<U9�����TE>��6��b=� ��?P��Y^���>����qB0�7U�!����e�4�k>C��������ʋ/�4�X�;���} �P���ȯuip�2U��/��ǘ�h�����ۍ!���=A��N�q�(�~��}���2�B!�ƣ�F,��'itT�F��!|Ko��#�%�TJ��ؓ�+2�Sv�,N��\�7��ᘗ���ayS�s3k������:h�O�]#�D��SP�rOAl{r)�Ё/�X�5\���JjN�'�&[��yx(#[�Ђ�>D���`��k��o�c�ֽ�p�ߝ����=ǅ��Is�M�z�0s�嫛|��Ȇ:c"�
��tc%��?�qy<�OU��]�N�a��O�<;����A0�����I,����B�5�k����TR���X�����K.�}l��u����
H4p��9,_%�T/�q�{��L�l���?�>9�y���'�l�V��ҹ�4mQ�]%�"Cs�h��8%�\��L��bX�-"o ��Aݒ�Mu�`B�eE�;O��k\/��c�H�r�Td|	8�ni��6�M�i��������G���������;x~�k�d�f4�҂�+�|o.M�zZ�x����C��O$�{��g`�Pt�'s=s�ltW[xi��lF��B������p�|��Y�}�x!x�d���ƿ4�����]�Rܭ�i�$W���q$+>�<���F��y��MA�G�o
�H���w�-<99�y���K��F��u�������EV��P�q1����՗%6Z�c�����t_������
��O��<�k�4�1�k{M5?�Ih�Y
�Ϻk����)`a�i�xzX�@1v�{2:�y�l�t_~����z?|`�4�hk�Q9I���rS屬�Q���/6���a�3WtǢ�>��^����)tFbo�/Zi��{>ͼ0�=s�^���� ��\ϼ�
��qʰ����Ay�8��l5Có(������"ď�<���U�kBK�\�u��
b��ϯ�#Y�PQ�m*ݴAȵQ����5̴��=�+���Q�f�=�g]��[L3�^������\Un�l�<"��Z1l�c=�4���X>_%Ifk�)�.�؂W�?G^+.��fEِ���@�{���k��L��V%a�G,7 ���Xfx(%d�A�g��,���s�'��ض�1,�=ֳ�Z`��n�<ܸS�K~N��IV��trs�kQ ί�4���LQ,Wt�6RV��4~�~���j���@��`Y_��`��[~ӿV�h���ݳ��u=X���\ш�K���m�3hl�H�#�)<�0�����(ix�u%��C��N�F�ݼ���E$��ǿMC� t����I�"�����pΐ��*��$���@)_�4��=Zz�e�[�P%�4.����ga􎩜g!��^<Tμ�u�;�s�cЎ���gS{����Y��W�9o� V�W��o�0IؖM��{n���X��G���9L�c֌k�	�F���ѣru$?4Zf�sM�
�Y�I�)}KI��p��!h?�B�"�{q���c�t`�c~� 1j�����"��<KLfa���ْ_ݐy�Xpٺ������f�պ~WQ@="����Q��R�h&cָ�ϱ���e�4s	�C�F�Yq�w္GT�����ps�0���5��L>$0%�4�0 !��ݨ�BAf(���w������Z1=�:�)�{�u��vGxܨVl�آ}�1�l���%g�P6�iwӷ��3O���h��=��+߲���؃J�+���{Jn��B*�����ԨÃ)H�w��GH-]����P`+�r���1�S�$�*�>Ĭ�[�OmǙm1�t��W��1���C<Uk[�h��r)J�A������]�oO��ƒ�������3���N��XB{�%;�CD"�u��$_�_P��/��i �-�G��ԚV�[r���#W(�/�al*�%s���Ժ���9�QJ��S�g�@K5,B��c�VN��T )w�q�ֿ��v�!���^�U��q�H�qi���.�y�
�hs��>i<Y��֘'=X�ftR��o�66F�Q�\�`�`j#A"�v�SIR_RN�<��P�DB�΅�W��p���[;�-u��HO��̋"��(`��[��I��ִLq�Je��V��0�W]+�����iv�qg¡Y�ю�!m��6y"v��fVu��k�"�323n�7a��پ��.e؂�t8q�@�D.�s�I3�X�,#+��1�K�L���4�w�2_<
�A���ne>�+����0z�4������wI���?*�p�
Al�9i�q�W�'YGcA��m�	4;�.)Ϭ  ���9'u�lܳ��`WB���}�f~�_6{ﮑ�#���跨$\9��&˯NǷX^��i��Mr����#�j�_�r�{ͨp�=oj���$����u����==��ti��\u��%&a����֞��&��Bv7�i�I�	B�����2��V���U���/L ��?Ĳ����s��/+���	��	ڋn��oa����)�|N��J�kV���P�[��H�ߌ�"�	�4rl��&�l�}� lJ��G��<���y<��r��O��8��cbn��;�,
?~��8�m\ܕ��V�K��� 9�}�'t��KsAmX/S�6��^�F�{'?���vX��3�(�G7����/@1ߟ�*K
{VZ���쾻X��E��N����	�H��{*�P.(�ݪ��[LG.~j�����;vZ?>�/>�O@n+fV�t*KUC�FC-�|���&|h��kqG�41�$Cl�7i����y["�\֩����3j�6�F��,e�E�zY+_�ٙ97�&5t����A��DU��=f��$,yd��޷�H���!#��d]ʓ�_��tt|*d�QEJ�=��?�5�Ո�v����4����cz���Y���,�\H;�j:�VZ:� |����D�qn4c{�N!�4�^��j�	<U�Ь�
G�^L�(���}<��p�d���0�Z%G��p�R��{Q����ʭ0�<���8��@,o�U��R9ԇ��I�D2�W��a������י7�"� 0�v����
��}qL�^��qP8� c|"Q�S8�4!�	J����b�FZ�re�_oP��n�3V@������s�!$u@a�������oإ��M�|L���8�K�]{�Ҿ�K��<�Ė��|�8�A�ș�׼]\V�[�}�[8�b�I�ʋ��Balry�hQ�� �~�-yt��F&���{��Ȼ�.D�s�"��U��NC
��!1�-h5}�!y��h'�K�܌�Ypɟ��z��'���}�6e/^��+�N���*�֣~�
�=q���LI�8- �J�8�;�����z\L��#�8��z&[�d����,��fp�|�j�҉����P7��*����Gx$V(-�ƭh�%$2����ʦ���5����qİ-_4wV���fFQd1 h
������y�J���E������l>5����>N|F�^��|=�,���-�kV��7M�_�r'�;����l���v�e-FZsCJ���TuےW7@�i���d7l)���ϒ�z1��R�3{�ؒ�Q�)�ߵg�(6�K@�{c������3����0-�������H�r�uz)K"��GR�B�="�Z	���L�%�`�A��>n߱V��[�>����<�\��ܳ����w��nΤJ?�1�v�Q(c���IV�C�y��|=W��g&�ŋ���#��	� ע�hr�˩GT�M1��\��k(Ƚ�j�_�E���I}q�&���b���EW +.�'x�j���7��}�z%ES_�V�Uj]�N�
>!�K�c���0�#`�>q����.�9�so��,�O+�?���ŵ��d�*�϶Q,���[��(��.ƒ�T���>�M7?����E|	5�z�A��]��V�6�����Ba�1���w�u��4:VOF>Kř�q�a�	�kj�~��҇Ͻ
';;�(������Z�+# .���W)��ל<�-�T/
�ip�d��czFu To��T-!Bo�X0�}�b����Qӳ��@�#�+g4�9�T)2M�͂��#�^|i�ȅQo�\݃�ڀ�aQB�׉��uQI���E��=���L�S�N�����gڎ���C;{u�[���خ�,~,����z�K���V �n����y~1U����HMA���r�#���O�r퍢˴�|�����z�n�j��:�A���mt�n�$��kڬ���%�d%Nla|�ڵr*c;� :K��l{m#�e��_0��&EÐH̞�������D6�3=�$������8#��ff���66D��g� �"��F�W��O��k�93=7�'D5 pӁm�>�m,N�yoe��$8�s�楍u}oI�
�w֠��Z�(�K����ty"����RM�`ki;1���KO�>nrʥӛD������K@��>����.��,�����Lp�Ο$�:ZV(���w-B��"��7VIF5l�[b��?�K���;5�#w~29p��	 y�������,5ӪC���C�p�(�~����j�2Q�i�R��[�2�$,��އz۲N���k���C~D��Y����m�2$ݛ3�'�Q�
f�I�N�icGP�x(���NɎ�W���4����ⓉI���11G�[8),��Q�}]P�7���o��g'�������_�5as]ɜ���I���RU*ܓ"Z��*3��DHk���-e6@�B��.�Ӻf��&�81M��N`�p�ͨ�ٶ�óg}��8�_���k���?KT�	����o�zdG|��.[��E*7��J�����B�^�������$���}%�8cf�il�;�%�Y�����2�,��s�k�e���DW5�;o�|ܰ,[m6a����`��"�/�樦��x3�Ȳ�_����/�3��Q�����[�R�V�7�}ln�d�������k��qy��-��T��EA��(f���Y�?-�{�]�Z�b�}�U���!����QPcJ�ѯ�^���YWzn�(Gٮ6r~���' ʞZ<pn�ղ��O���T��m��A~�!K�5��#�	Ŗ���Y�'��ji����)����1�eN�6�D�^l�A�+� :
�xB�����}�~|�QuR�Fo��n&���i�ӛ�����rfl���O����O_E\�F����3��8��x�-Nsf�[
D��~j��ǉ�&�'S� �b+IZ�Z�N�$
E[�0e��4�Ԋyc���k�<$P���6�gow �1��Y:⢵�Xc���W3 ����dw*'������3���_���ۚ?X4��DR�  ���\ͨ'	�J��?���pq�
F��/,�.^��|�ܴHY���l�k�:��5!��ܙle���i�#�?��{�`��)���౦q6%a�����f-R���@�fE%�|~H)Fh�97?c�N�y8�R����Or���@�ؒv��C��4�.~q1Sb�7��hs��cvn �يL|0�848�a�4���p\)��CG��{6_!�r��^?ͥa5� �?�G%��g2�/����"���!hs>�+�� ��I�J!�=�B}>����·���U����Q�H�4l}^>7���%�0�o1��-sFHR@��Cmʪ��X���Էg�p�����0�Nk{@�{Z�c&�<�ER����z�Q5kBȺ>����h2gV8�5v(Re}x�7�l���+��^��s�8��y��X��c-�QkaB�Y�����`V�� WD|
-(�z�~�^5(���F�X�B���s �M�*V��f#���G�1������K���Am�1	�sB}�0��(���/M9n@�=��q.��� |*��n Ag�lo�##`X��U)��~<?�F���a�[	�s��|�AjŇXg�u.��yV��
����,y���-�b����0h4�Z�|D[�6_R���	C�$:�"�)����h�K���®�x���R�G�Nn�z,��3��������qa^�`j�;Q��B�W�U�خx�
4��L�y�_�����������,M�{�����M��}lX+�ң�ٌ�Qy�y�	��V�~�yxyW�O{ȿ�,�PL��erF��p�K��^%R��G���ANM��<�@S�=g�.?Z��>��`1�d�����p>h<3᠋�ɜ������|V2K1�������V�>߂1��^�b,߼�VҀX��y��;S��ݓP�ʦg�w_�����g�IlXO�lw�{�i?�_�
�Bw��RO�2e2a$�� iAր.����s��i6����5�&��u�(D�o����R��g���V�������{�z�71˟����i��+e�xc�D[��<T������������R��Qe�	�,-g����t�P��E=�5/N�{�u�sc�0G���O�ց�1�½�[p�r�¶G�k�#VJ,/���ZnW�>��9���/E�X�h"��wP}��
W��8~|=�����&���?�f�3;� �o)�����d���y"�X�E���Bem���~��Lt�	���_�o_ǰ��s[���W�[���%����\$�+ʺ~:� �o����!) �2�'���"}
��CZ��q]^�n�̹-�2����6�ʪ�m�ϫVÆ��&��Q2vk��ƾ��b�9��[���hf�Zƺ@�Y'�.B�t���h�^��o�N�PO��&G�ӔR>͂��)yn#~^�$�mi�1<fsYx+-.�dh��G�c~F�[H�F�z|�:^π}�Z)��F�&xw��J�|q�Z�8�m h
D�E�T?�¤q�����Gb���;/���6^�NYE�T���9�>�؜�p���3�Z��9���=�<z�էգv���2"�c�#|`i�׳���)�0��c��DM�]�Wv���ӯ�����ka�=#H�~���د���с�x�f����&	�2���r-H)��E�ق�4�K��F%oZ5�����$�{pG!&�j�l}2ZԣSS��[L<�.E4b+���>@�(���105���7�&H}�Ռu�&65�M�D=f�+�4}�6�&c϶����8w�Wrs��&̛E26(�A]�<�ڥ&�q�1�u9G=����®	��q�*5��!�<�c��"^�	�+��^���X�Z�]Y(�Qy�l]�
�.U34��]���h����'��~�@��Id��y{_����~y ��.sq9�O���v�:��2b����]_3�3�����s�MD��ۗ�c��� �+Vc�L#��w��ݘ;����B�jSY��*�䤸6� cL<��dʮX\�n�=�ϹYK>��u`�,\]�k����sKC�U�`^��V�bNMpX�X߱E6}�%\������e��Da�Uvː�ڞ�����̘���wf�(G�] ���9�͟���Xv��^3�'Q2�]��ڽ��V�5�$	����f�l��p��m��)��3��:p^��K��*��`���@]�в�7V*ݼ�3/}�D�%nn�K�J������;���&{Ɖ��i�|�v)^ʀW)̣���+ |�dQ�[�O>��8�㪰����_��`��Y��Y�m���JU_�ckӽL1�/������!]p^�Nj���4iA�|���f2
{U�S�S/be���0��
Q}�4_�.���N��v�QS�!��`����֓� 7�fC�az����O8��۸���� �N6y]�^�Z6��S�*Tal��b�z��d�{�9��GZ����[;A�1���j����k>m3/��lGx1��u�7(B{�z6; ��L0-�?u�[�|$^R�(~;�a��nECj�1>X����(<���V�{v6�E��+��F�>L�oi�"�M�>�� h�)��Vq�\WiĢ������G��X�6�T/18��Q���'<ִ��W�d|�9�*6о7�ez���s���E˻p�?��e��Q�5�Oč?���_��r�}�N���5��N����{Z��[��#Mc���Z�l�;�ɕ=x�K��})T�4�%?�EⰂ��$��O�Piσo�� 0�!�4j�\�.rf��su���:p�c�/?b{w:�/�-��:@���U"�<F^'�h�Y��I~�2�:7�œ��qqvY�����"�k��e���h��tZ����]:uVq�݅�ն��L�ĎĄ�|�K�~=����k�$~�a�?s�#�-ZΘ��@�D�K�@����Ll���X�h�`4�:<�����C�N�V ��P����ᖯxad� !	Pd�/��0�v��\_>����0ٙ-,�آD=P���ƮnIX�[Q��d�@٠����]X.{�DMDw�:�L��/w�m�K �7�j/�o�2v6���)ZW�{�Aq�m���3V����P��� %'��p�f�t���
��?��u��%����|��+t(4�Δ���K���7�R�A��6lZHg4[�.�c��iB�Ц,�p�^�z�+~����%���J�c�!|/i6b�iq��߂��ʁ�=���H�Q-]6(P�g0����G�0�#I��N�8�Ͷ�8
���u������ �5)"X����]�p���;g���J2��� ���s_Ċ��k'���4��)��'6uR�C{Y��Z��������mu�M	[
�Ś
U�u{�����"�J���Yٔ��OV�9Ջ��~H�Q~a���2�5Uo��n���@�p������{/�CUA/��7���8Yc���5�W����_$Ģ]k xI���D�\퇉�w4h�,�yz�	�O��XQ��(��<Dg����k��7G��i/*�X�6zW�QH�T��%��V��n�N�U�)�l���w>��ހ����3b$���3&l{���2���q-�2zT��D�D��}5��~��aq��:M���l���78n�i�k�^��bL����/���/cj��t���	�3�iWln�Y��~!8W�kZ�,?B� ����+'�M��H$$ �S�1!b?�Ⲥº�X��M�`k�M�g�S�<k�c�)"�Ǩ�-�̽>wʶ����g��r�u��R�B�!*����KcR�%�B�d%��U�ෙ�f�	��g��.�"!$;6 ����ժԏ����0���������x�A�*���I�iI|J�U�	1C�FJ;G������������"�a.ç�e���1����6�~O������TY������:�:N&{�R���=���?��sJ�J	j����!ҡ^f��<��4% �����h?���+g�5?�����ʼU��k�ʿɮ!�.�^��*ʷ�;�`g�A�E��)Eb���I�����d&)�#�K��8�YM�X��Չ��G���+LhK7j�!�9:_�;�j ìQ:q�{v:w���y�x�L��Տ�,֏pc���F�� ?�ƨ�/<-^�K]y�.��E�6y5]�`&���J3/�����O��>p�P��CJ�:C�8t��tr��r���4tWp�%��T���y����qm�A<ۇ��%�`Vg�����`b&�ˁ��ـ*�����R�M���2����Sv�a����k4솄�O��#c��B_�_Yu�q���Ly�SRXs�y��}����H��u�֔���X���F�v��ۄ����[_�֬���qp��4W�K'/����S|^O������KU W����1L#i��P�(i%H������E�� �*J.3K�?TW�劰�� ��޲*1o� ᇁ��U��pwD��	b{ ���e^s)FW��sLo���� Q�A��
�$���?9r�JK�t}�e�22E���]�c�V������9X\D��f�x>�%P�����$���������K�К�}�����2�����)��ދݠY�����'4�I�W,	���@�Rc�EW�Ei�P�'���64W��i\����ɮ�����I�E��aPk���%m�o�x����i����MB���n�t�Z��P6�)�Ř��xtMzG� �G	)Gs3><BC"".UO�)N���[v��Da��	�MGj����8��xR�ն��6	TH��0%�7'��S��$,~ׁ�Rߧy���l��܍@����5�olƔv�yG"~��H����%ђb�'�������sSsj�xp��:
�"��3���FrJ�#�^����ӕ�tʜO�������ŧ*�R���`�@k��]�AB¦���Px�$}Tf�i}��7
�w�����l�mF=�MOf<��;��+��V��*��̻A�e�/ǚ�D ��J(�(���U�J̈́��@fF��6�	ڪc�u����2{�F@�]�
~I����=�YSȏ�Js�j7>�!�|ۂ�Uʒ�Y�=��:�4)@:aB 	�����5���B����o����I����`���r��rם���\�{"�W�ߣRs-r��w�)�;�J��{�'{Qi ���Q@cV�4�^x[� "�p�N5J30݀�n������Z��\}�������o����U@d�ۼ��!�?S������kPκYUӻs?�y3��Q\0\A�[�N^����9%P�s���A����ܬ���+�ί�@����nEcv�#a�HJ�Q�Z�����q��F��K�b
�l�-N9@�������A�m]�����Ԁ���\8��ɛ��0`���0�8�h��?FC�8ߟ/����9h��A;�p����|���J,~���0v2�uT��y��b�åW�1�Q�S���}2�4h�o�[
�O�cP&�J1���x��i3p!Y4��6�wj�7�H���m+;��_`��,��{%����ð��7�;(�D��'�i�o��0��g�H�����@D��O��g�^;FY��dEhq�R��d�r��&{�	�����3z�oCU�W~Ӥ�+kY�K���.$����B�4��3�)	�T���L�5�����1qz+�Cr�:��>�|�ض���/
�%��k��:�8+�J ���č��������(��d��|��8i3	a5�P�����{���H�X�X�	����yl�ĕ�g���mJ�q	�cׅ�6[�p1������h׆��L�6j٨`2���T�ܝ�9�	.lQ,�j�D*��q�y=x�������+�\e��?�ᦎyH��RE&gN�7*g�bi+��]�8��jw����_+a����Gp��H���~=D��4!���9WlU%KA�:�fx�T�Lё4g�t�9Z�P��H�CO�ғ����);��.(�l�,y	��	$�%��LW
���EC3�A�S�@x��V�Q]_}�g׮�?Mw��B�K��%|���kbK���WD�����c���<��t���Y)�pZ���Up^�M��J�O�v�a"K�$��4-mE�j1��q�	���PF�/��>@j����_����!�X�c�v�ڧ�#�{B��"�o�dё䒀��21W��<`b�7�r::����_�	���Q�򇒯��yFe�C��9���\�2��K�gׇ@d�Bk.ui<����B9Y�Db!rA��B�;��o!gyb�Фj�N?�P��~ɇ�W�̕�I�&g�����ڬ1�ד�(�F'T+Eqc��N�:��FsLy<��*3y�<��Wn�e��"����gn���Bٓh��͏�[�K��:�>5�y��R-_9W׳�;�c2��GI��Х��z/��T[A69/��k�=���X;R�p (�5s�MQ���k��3����4�a��&q��u���:�zQ$��ܱ�I����
.b��2d�1<:��zkʔU"�����ٍ����$�9e%�:��LP"��M�(���4�����.�G|(���X?�����i�%�1�� �L`H/�c��ҟH��=�(�9��s>k�,��m,?�=A5bB��WM3���cw�f��w�T$G�H��o?yx����9�{>c�?���Čy��䘮��D���>R�D[v��:s;��Z^�5r~����S��L��iQ�.���$Uۘf`3l�tn��-�'���p¥
��$�/�`��!�}kiR{��)�C���sF��/t�%w�H�������u�],���0�������䧵�0`����_�&�<��4֐�g��4�A)?�xLTv����zqWs�D��wb�	N�)K�s�J����@����D�@q/��7	�V~C:���-Yt�>�b�~\d�?��Xi����p��G�ȴi^Q@X���f�*�	LHc0!ݺ���W]P�|���D��U��n���E�$�K�O�q��T�eY��T"݈��*��g6�%��-��M.G���d���H�I)��NmN��J��I{�uNpDm�[�8RFIG'Ny�����b��O�/$dȸ�p�~Q����K�tCˬ���L�����=j$����cl�ТzUp(�>�~�rP�ꐨG��i�f9���Fh������!�Rm&#ܨ��Iǹ	�~[r�'�hZ)!�y���>�b� �ay�m�0��Ӂ�������G��3x-�� t�$Y>���b����zU��TE�4��Ȟf~w�l?c_Vy���rvK�)M���؆ك-|�AB7)O� ח��Ʋ�16T����5��ncs�� v�&�/�*�N��� ���ּ�B�iŢ���+�����X5�k�̩����_��93�b��L���»= H[U���}�w�1*Z�ϊWoY�L���!����B������z�[GDE���Cѭ?�{��#�&�hp����xB�W�^�)!w���+T:3��Ĕ�;�tb���S��{��O*�_O�z�B@���<��_*:�!�jdV�։.N���z���h�L��{�ɏ�b,�Z��$���<S �-�v �4�-m�kޯ��J"�Z���:�w".6 F�\�1ǣJ����3m�#e�4��~e��;Y��`Cc34��k"�B͝��̳��'C��гw�eI�;�
8rH���h����[��Ό��Sb�w3�j|8��9�QA�
�y�Tx3\O���p4Dmv��������6Mj��&؜� �!�<|�U��̤���j�W�����發3Jd3�3K[HXNcc�����M�qP&��w�qȻց������Z[��4N��|�ʚo��.dB�������K����p^�:�RY�?�������P��P;��pi������+�Ӕ��C��_έ�������`Gs�3���/�x	��AS�c���T�Ѻ���O؄�������f�/1U7[�ϥ���q8T����/5���������w}���۴����|����G�b�,�����@�^� �D>⑛��v@�{s�V��U�ƒ&�* �Ө^pG��v^aABDy��'��8�`?����am�����BZ�e ���C�U�*[ ҈0Y�*��l�ea�D����"��gN+G�zL@�#���%66�$u�Px[;��09:�0�E  ~a�&H��#�Kxgh|�,������撧��$�Z_[��!U��_?p��8r~�G�G���� l4�d�l���q�؏mH�҈k��P�g��A6�(T0���?��˶�&6��)̟�5�14ֹ�ݷ��h�U߽q��P����Ǹ�B�"�c\�Y�zp��#�ݐI���%n�(����V6��/7��d+Z���z�f'�k쪶s����E+�	Sڮ�,��ZQ[�1�K�1�S	�	�Y���ݴmOtdw��2L;���&%������Q���?��H��DS���UH�T7��j�F �H�^I��B�X7Q��tP��.<�����,�]��]�-i�"dv�_���LZ��4��=x�q@��^��*>�1�j}�0�<��@�L���D���Im�@�=/��-M��4g��襥,�+���`V�f����E��̟�/ B2Dl9�3S�l:�c�&���*J���Q�V:C��ɶ�J�7;>�,J[V�W	�ej���z��l�T�ІO�	�L�����NֈX0g�f_���+�%U��gy�f�/\)�a2?Ξ �4�ՅZUm��o�I<���@�t�]��}��� (7�N���ы3���s�{;�&SR˩ ���]��w*�Y��l��(0=N�<t�j:v}�_\�%bT�i)h [��{\ǹw�����T��4�U��$V'O�jk�Ж��
oo=a���ӊd��i���[�vm�b��N�M���,�QV�6sG��y(��=f�_���\����{F��x�Ѧ
C`�mY)V��R$��J�`x�h��|�F=����f�
��W�{�-0\�����_���[�[{@��<_��6��(�Σ\�i��8��3Rlww�9��[�%c�W��Uު�e��m�w�2'��;�E��C	-w3f�k�WEBm��i���*��ڐ�b���ԊȖOu�oXW�����)+��n��֨j��	��q�|�Q4��S�^KD��G���V��ϜJQ�ڂ�0�r��>��8-7���>���.� `3�W���v��ᖣ�5=�H�<��{\�R5�hM[�TN��w�"���]�}��:w/���*{1s�}0K��RsS�{<�@���W�vLF�|�9�xkcW\����};��o�m�������> M��CJ�Z,�X��@�	V���lf���0߁zs�����裳`jt������s��0W�*����bH���O�uZ�m?���M��A�<��[_"aC��(�ă�G�K]&8Lܖ��Wr)��1��'���TB#�7�;A�5񚟰���������(���7GJ_������ٟ��צ,�'��i�`�R��Č����J��W�<�g� ��K�(q���=��(گ��R�LB�yj��K�T:�(j����j��˱:js�|{�ܓ�3��Ca��bϼ��у^��6�f��)����;;��q�ϭa(D�����t���^�.'�	QB[9�����%�M�fV��'G~�8[�AcH'	e��46)��<�7���*z�y�������D���@8��}gޜ��fN��'��~�j�
��k�E�h�!�}g������y�L������Į�БE�~��ɩ1��=�j�,�:�����JT�>�
��NC���'�KMS=�;C8	^N��*?��5hRϭⅲm׼�/�3�ʠ�v����{v/
�A�ߢ�[f+FI�Ä���y���ˑx��C�`+���i%��t�V���Y��9�!p%�Q�����$k��
�>CͰ��%�Ҙ7��=�
w��1?�h|�X+��ǩU�[ۼ�_�h0�1�31�:A\���_���I���;�H��X���q�`��px���.秊�(�`@��L�l4=�c:6�ͅ���\\g橥%$���*���QJ��B����M���|d���8�O�Lh��o5�������X_��8-؀��F|�Fg�?���mA��_���}.0�UF�[�fUB�y���01-Wઇ|ҌW��S�(Uu���o��@X��)hӯ`$�=k )U�L�N�w2 P�ao����Q) ��v��;P��q�W����u[?OV�}_�ȵO[Xu�jAR؈�q�J5��r�h���ͅ���d��{��trf��?fDfK�J3S<}2�tGI�^�������������V;�b�2�0Tk�X�/� 8F��KЛI���$����v:��[�Z�С�5�VC�%������~.�q�̪�`��r���`�AG�63
����e&H^���v��L�C\<�r���F���G���5ӫ�v7�G7�@v�Dμ͠�$�,]Q���v4nހ!,��e��Ry\����.�/Ņ$�z�+�[cVz�����	��:
g��Y-���u&X<cs2NM%���p�Gvh�4�?e�2d~�����s�E���3mɪ�,(�w��Jߞ���P/�/�zi�Hm���R1Uw��Ll��V��%��?x�LB2�Gt��X�������j�k���YgwzL.��zh�E-����U}��v��F�����8B����[��Ɵ�2��k�{q��:61��$ǣ?x�`ϝ��j3j�i�m~��A�*[c�Nt��Ud�k�}��|���z���S��.Xu��"�h5����xya8��9��,�?Ɉ#�����0�Z���J�R,n:��zA<�����?(�x6<�h����~�ь�6v��vx�o] ����-�l��ͩ��Y��Y%:,,���JZ<��;w�j�ĝ��`$������3�*}��r���! �0�u�c����[}b�Z0�Ff|l����{�cU�����^��L��Q웄��W��_Yg87�]�����6�^��B��0�v��3w�d�TZ�
�t�3�]
��Y:�� q�Wm�/*��OjN�b� u<��ܷ�^�g,��\��xm��>͖,�0��6��񱦴�<�R
�^���`X��� y����bnS�MτH�wx��KE�|-�	��*��F�a�¤SX���y-�7S��i~��K��X�6�S�hV�6�������$m���-2~X�ǡ���R��Vm>h+8��_����>O�y��y?�p9z+��2�d����[�	o)9���M��:�ַ���2Y��D�%��Ξ:rHl"�@�\ ��J�uOG������!+Q�ǀP�JJ��?D5�����e�`�M-���(��pG��A,z�H�AdPBzs=P�0@iN3q�~������9뀹�Yp4�)���ヿ��3��o���|f�7J�q�G�zTLލ8���!��d��,��м��(挹Ȯ�������xj{էq|�ȅ����Oge�^�|�Ǖږ���h�:��V~&z�h��3����aӓWq��s��rk�F��n����P�MZj�_'���UA��V˰�e'��\Pi��[��>�
)�)�"����m�{�y�ڄG�\p����,P ��&#��5G��>�gӮ��B���L��N�sv�YX1)���)�Z)�n�83[C�;?�ehP<�?yAl����QԅTf�Vn�������$�&1z����+ٴ~����Nw�d�Z��*��,�56��z�=��]Hx枆ծ��t>A����솿��̳�yx����e5�1���-ҙ�(E�˕�L0s���N�Vz���HP.�(�8��Y���^{W4/҅�ҕm������_�,��~-D)�z��X�!I�O���>!z�j��|����ş�pw�
Gx-#������(A�e�"�yDT�&��
o�Q�ۨ�ƪꗟKŧ����3�aK������,݆g����`���[/(�;Us#�J�ci����N�m�1���x��
�3���|��IƷ���r�kf1F��w���Н������ ����D��-]�j��a�d)=�7؟Ӓw�Ǔ�U����:���P�>l�Ӭ���6�8�G�ϻ���B�

� ��EuW,JRS'�,KHY�e�K�5�a��W��_C�d��&���5"�W�slA*j*S�inۉg�&���Fo�|8r�_�(_{f;���l�kR�#5�,���n�'�M�&u(��=���l@��n ���6!�M�J�F�@i��eٽ;"�k���S��Ʈ�
�W�NUK��Y�t��6m�l�����}��:��{�Hs���KE����m&?�?f.�?
�/#X�B�b�բ¹���h�[��|�}�h���-�T���8��.����\���NA���u����s����.!�����D��D5� ��mx�B߂d���?������X�:��-���ε$J�@2'?�f��ŏk��W7F՟��1���m����^�BO�O0\�����l>!�^��d�k�D�*�n�������6��rme���UfF��{kI��.���kK7��2��X��̏�;ޟgÑ��K�E_�r]�an�o�]�j���N���}��Ќ)7S�{^ {��Ko!�r��/�LԵ�9(4�@�Jי3�㪲�3������Q7�
�&�Ih��j�E ��S����pcy�F|�=��`
^��_J90�\T�<�����>�[48���&�Z�{���$7���ٽ�Y��ۇ��6�Mbs�3L�8�uF3^�kI1���轹5By�˝���uqO���s-O��z�r�5�Kd�<r��q<)�.:$o�]��$���P���Ǚ4�䍺u�'*�[g ���'��Î�ㆄ�)�F�b�1݆o����:g�����k(�tnN���5��F�6�$7�JJ�E�S8x�0�2�~>�dQf{����Owb��U"�5�Kw�6̘MA@,�
7U���X��*���C�}��mk]�y���,��k
�w�����"��\�f��.Y!'-�
�V����2��T�u��y��Z]��a%�6r�x�a�0��q���t���:j�$�'#��Ϳ��v)�*5��(݃��w���W��ÏU��	��a�/t����Z���/LP>'��<����6��K�\�`�y�e	u�gxN��=����kUhnwL�����g�ö�Hyh�Ӯ"J>p-|eO�<t��l�Yy8���_'d�˟�-a�(������o�h�#�jf�����O� ��3�%j�#�8���Di.��b�zHI!�POB�C&�������<�*�(�E���r�=�ғ�E�d��A�l�Li4Ff�p�nj�|ǲ�c�!�T��.�/jcYu&'�0`�ݜM��i�W������c��7�R����$�Z�S�[���JڌO�·���6��н�%9��洲���5�;��DCs�*M\�K�1H�?�U����늴�̀{��^70B|�Â������zPh"�w���V>��.s��mb'�a��+Ō�>��\TX�d��U�=�į>k-��'���:$%�d̺�1x{�n�QȍE�P��P"M�3�����aXs�	�w�����B�*�q����{�?m�{��o�����~����FՈWT_��J�)�@�!�_y��)u�ni�]��Kf�s�@Jtٝ�k�!�N�-�f�^�cK��ؒ���0���vUz�[@����D����O�.�GI,�9y��[5�R�l�����jN���u��'-��-��]dA�>n��̱l�p��¡<Á�w�cU�3�A��?���̼G�$7ftjxÌ�3͸ vN�$���L��l��U$�إ�P�~���	W�~�v)���QH���ʕۋ�
�F]
iju��z�\G�T��^���kd-x׋T+��Y�J�ȱ"s�J�pt|f7�C�1 r�5��W��m������`8���7ы��?R�Ie���v}�,�& 㣊D|Nَ�_@��(z�`�$E��K� O��;!�{�";�������5��f�o|���,$VK1����kM�P]p|��8�|��&��AA���3bv�nGgT�WfRA�9�i��u��Xs�A$��[7D쏥Nꕛӫt����V^lk'[�뒩�~%4�*�W�y��������?%;�"Cd�2ul�3�G�	�����^_�����h7���4���\j�N�a�#��qd�W"*�BVyFG��с��+��Bq�AG� �Z��O�bRn@�ݛ5%gʟ���8�:)��zn�P�i���R�X�Z�\�?�:��T�6T���u&��P��}O7�������m���q�˰<E�G��\�='��f��� ؘh�M��)�����OIe�=�~{5�V	z��͏�K��6���bƷ[�_��f��=���㋬t�J>3A���f~Z�,�aPWw~G��t�`���V���m�����n��V�6��fȟ����v�g�����ꮑ����bY�]�{�^Q��g�Id����dP� �Ve� H�G]�c2bUN%:��覧-�I��T��J2i�l�^q�C�j�%=�"�Q�do���QM퐢X�=w�o�=*^��9�C��:QRv�8�B��a�nhv��S~D�n$5¯�i[/��2��d�V�T��
S�N	t	�-���[��V""]�e�Oa�1?c/u
�:���4�}#3�DS�LA�R��[�y����X���wO"U�%�v�`������E%��K�{RCcn��>��Z�_9�|ù��Q��HOk��&��Ȱl�m���� ��%�8�ʌ�V�es���Bؕ@v��)�v1s�O���FUiD�����������k�e�9�]�V�av4���O�����c����1u�����4$X��<w�h*jD;}���RjQ���<�ٷްa��������j~��rp�s�_�^�kQ�Q�Z�]�\!��T�b�%��1����q�qj�u�/G���o^&	�0���h��^�#P�������J�\����$O��M����=��5y3U�'EV���.3+1�N��i-�0�<Th�-ɤ��F"{a�m�u[��X�"$�Io<1a8� fB�qh������U�.i���1^&�ݺb����1�!)� ������<�����<_�����m%=;%98�h���l�e��1|N]Kч
�g���9��| ��V���TJR�~_Z����\upCM��j�0����<!ϕ��	�;���{۴�Xz�(�HL2)��P<>��}����Q#U�	x�����,��rW-� �:����Y��oڍI��^n{�*�f����>�4&��P�5�ܥ$��pd;w/��8��E��$+�������Z(�������Z�-u ��Í�ź�b�-"�u~M��|�6�����; ��:d�����	ɲ��u��M��Z&�H�� ���n�Έa�b��eL�za��y
�����MȢ-2"��@��33��m�2�n����by+�P-~�ן�T�!�jdl�xg{��9���v��hG5w�T�Ɉk/l\�	�a"�hВ
���7.���".�֩~�z.�>�D`}&�� D��Q{u�ƨ���$!P��J/�GQ�m�ˎ����MA��C�=8�$�h�)�A|��3�k+mJ�jݟ�;�5�!��P�T�N����ͯt��Rb�xE�����I��w��~���̆h�kJ�sSՒ��Y�,�x��!#�tH��R�"ml
6�|6'����5�Ǵ�7\oa��ƏzU��{�X]��Ԕ1�Tbm޴���S�ع�l�,��.�O�s�Z��ڀ�㲁"���)�ȹiO����褔)�$��GJ�c�e6�>�*�Z�,Tb�u�>YM�8�ekz��3��]$�|��"rs�G ;�xrѠ����̀}(/�;�7���n���&������IR���._�j��1��,3��_�yyW�gI]I��Y���B�x�Cg�˸���L�� �4<�)`P��J������S(��Ao����^HpY�Ӱ��lX->w�,DW��7y���\Շ�/^:`�ta�Ud	qwQ��l�'ߗݓ�M(�0B&�BEMG>��-�$�Yp��qpY8:���tI��T(�tU$[�D�h���2V�Ԗ�d��W�/�v�ǇuT�������7"ٱ[Rx���=Gr�>	O�|�l�4}�������V�AeH6G����������\ ���׌:�Rl���p�5<���?%A(p�F�qjѨE��邸�z���f3	?�E��
�շd�T�"C~b���Jw%�M��g\�z��/;+�u���5ޤT�q��al�9�s2d��f;���u��f1@�>HlZiHBA�O����?�*�����qv�-��-u+�^d�ON���=w"��P���t��d�`��6�RX��"S^7��=���YAC��Q�\�_!l��?!��q��=$���N��sz���>M|sV��38l�t���/�r����C;B����ņH9������'/�^p�o��]�N�*ծ�>�;q�؏�r��<�]Unc}���m�H	��fYSj�R�F��sw����54���~���?��~���,P�i�x��(��:с?�����E��?拸��:F�5�Z��1�enȲ�ӈ����I��EN& ����ɋ֓���Uԩ�h�^�5h9'��}~ay�d	@�����Ե�?@�m��+uA��cÄq���E��3/����L�y�4�59�2��ԉ~����7Β��]�pqp?�h�A�X�K�t<R�w%Q8j�T.�ZF���КM��/6��s ����056���`o���Yk�98L�)������Uˍ��o�c!�l�6��V'������e�v)��4�څ�:�~q\�9p�{�6�)�yGy�k�f!�(�2	ئ.������<;�s��=���?���m�S�w������0Sg�%m� u��j ђ�/.Ӡ�;j��G\���擮�2m����]]��M����OJ̜�b��=!�z�d
(�m�e��0�(&����-�����r[&��6���:6m�=RS�^��Jt������A���|��>Й$���ˎmcN�9E�Q�.��<�����L'm^R3#�(B�(��D��X���VQBJ���f&�E;�r���B�f�<�~:%'_�ʨU�10������W=&:Ӿ:Ml��rO3��	�.Y��V�Z�%�Թv�q��K����B��!��y��q�=P�0��N ����~Pc���q8����8�W�e�^��yI�{�4�h���z�$�u;�����d�О�=�0[,-̫
�*��9e��"�
#k�`\�D��93W��3ْ9.2�A�v�S�ћ�CpZ�B�V��Ѻ\6k5+���O�@�}���P[����F�"�_1��k�����ji���L-$�B� ��kDs�Ҟ���f�r@�>�=��OI:B҅#�*r,a sF�`���`U�Ϊ��p@�
x�D3��ehF�4�A��Ί��K���Ӈ�>�������lC�S��۹G�d�i���]�4Y#3�� D;p��6	u���#Tp*:�B4��Ar*?�����b��/�ބ���r��5ޕ�uF��EL|A�zd���\t�w�����,�÷A�J��Z%�����I;��t����=�i�LJ��VJ��Of�F"�5P��׆��a=�&,�(L��4�� B��Ue�*����՗���o��h�������ˑ���x�*�dGl䞆�VV�p�x��p��؈R�JE~t�4��Zn:A�dB��T��M�*M��a�ɑTU,i�Q-}U@+߭�d^����v�$����OH�ma�a�)'w&M\i��6�?��=F��b�]-+s�ڡz��$ �Yߍ�8�3�B��@򛻐_�{K'�W��j���"���k:�)*�?N'Y�
��ZJ+Ռ���Ŏ��u�<���p�1th�D^�V.� Oŭ�v?��y!�����V��6M��	�o`��&�8�響/����G���ۻfF졝,L���$z��K8��i�A��;��ퟔ��aߨ�IH�}+$ڻ��{^�5f�tT��]��H�7�l�z��Z|"a��R�Q�"T�PcƄ�R`iI�x�JR���Օ<1�1,�~�"���P:�V�����@�r���J&��R&L�L'�?%��~���?��+.�Ѭ#ڌ=��n<�$�@�ů��R,���&��nZʪ��=�O{)��4�q�06CQ{�/�k|�y��<M�=�ϵ���|��e��,�+�-m�K���S^)���g�_�h|t�/~ٓ�n%��(�����C������'�����#1	�k��. ��i	T����C̻���pw���b�Q|�����\�OS��Q�7�&):�έZ�0C ��g�*�Q� M�qDrY?Ky�4��I��f��qr���,O��(��){�5�׌D���"}��:�
� �}�3����˿*�[���	��W��Sj=~�<��P��D��g��N�X�����n,�T1RU:�3!�S���{���g�k����j������G݂�l�Ԣb��O��r��y\]�Q���>W�&y��~�&�����~ak��Kf���$��coe�d�o�%�~�Q���2��N�i���^��%Y�+�@�&��^��~L��ׂ�ZVv�t_)�At��Z����C3I�2j�q�ɏ�}J���rO\e�X˪m�A��� r��)M�SW�x�?�8q��-���h��<�:���!E	3��r��kQS6�%�D���\3텵�[�Ul� 6��6/�m�Q���͜w6lu�NC���>���҅<�Bn��Nao*�ߛ���n�
�.����*���+�c�w�� >d����?m�� 33c����OѤ��A�)�y����q��[��&NΣ��j/���Q��mbܓn*1�/�w�b��O���=ם�K0N�P���u��%(�#T�> �ַwEً�8�a���8��V��E�&#�+H1�v��A"������#�����>Hz�6H����w-�_T��cJ[��Bm�ݶߵ�.����������\fM���FD-s�v�Am�Z��-�+��]�C|�xG��
o���J��#�bj��Q���d��Q���ku@f�
�v�o��%�X���`�4b��y￧��!�������T�)���K� S�Ν�+H�'����g��J-yүy����Rr`î!�m�`U�5�e�
fָj������f�\��]�W�쑑�=����Q�ʺ����,����= ̧T,��J�;@�)�2H��}��9>�}Q��I��D�
90�.[o����,�O�ڂ�o(���c;��F|�k[��,��_\�h�vOT�4��v��ҿ&x�l�R�Z���]>4(���y[��3��t�Ɓ�⒅#�|* � fgf���p`4O�Fӛ=����<�ˀt7M.��&�����O�c"zg س�wS��!!�A"xq�ȍk�1�:?�Q��0��
Cp��'K�ً"����A��x��
�rμVj�f�C�_�RH��h���GT�~��<d���ޑ� 'J{c)""�E�u�L��W]4{%�4� {����2��q+�ʏ����6�\@c�i���{ G�K��4D��Oǟ������S2͊��B���1e)�Q7����~�����%�T b��oG�A�e5ϋs���?㯊�P}֠�l�[��6��,;a��'m1ca]R���'�2zOr�A�����	3��U	�p�{}�3a.P��P���:3���˯���o��`]%�)b=16�Lw�>'�0���H��W��2=@O�dX� �F5��32���8�Gm���G�����\���:U􊿟�Ha��'Ϻ�x[���_Q�'���ĆC>6K��\�G������A@^��{Q$�S��Z�N���R�M��3=�ԡ&�CoN�7M{x�]�Ͳ��j���|���G��'���� s/)~�o���^y���nn#��{�.#63�9�&9b����/����
�jH�5��$뢁���|M�T]��s6[&���Ə�8��p(:n%�ߗmI���HyV�w��������?O�]�L��((i�.��Z,i"�])½��<���7@��7���} 03���U0� ��{��˙�[<�r4~ %��ٜ w�1X=���'z��ݔ�p%0�oB��]�p�d�X�8`���{��i|��yOj���d���"ie�+o� �U%`E�v~��/��nf�0�39�f����gd�����'�V6")O7�J���u��d�9����������؞�"4 :�@O��c�DJ-���t~5�/=����}��cP�S�U�� ����,�VS�������[6�6�������&�e����/�V�^-�s���mt������Ŕm8-6b�o�h<���Y�cw���'o|C$Ȥ�WN�I�sd�_�uZ7��u����L�"�����x٢�D&�΅+x
vmf'ȓ�I�4�B�n�n����m�$f1S\���׍k�D��pD�����i&wjb'����x���g!p�5=%7xɭ}�bh���vwh'�g���{û_���}V-	�.j��mK��*����M/#���W(g�sw���N+��:{���	�y4��ml�4�tZ坍ڮj�ag��[%��&�1զ��ǹ�-q}��W�(�HR���𛞅��z[�c���?��wΩ�J ר
3d�Ŧ��u�%��#;�����T��r:��b!�܊������8��x�
�;��I{�~��C�� �N�{��g���b��ٻ��w<{�F��22p�&A��s�L��(���)Z�,�Ų�V�}*)<�aH;+��{�Q֦�Soʉ��U1��>e�VX��N!��c*��eا��N�">�����j�C�x�[���ҝ1KM���YO�) ���?5�,�+c�á����fa��v�s�IC��
�(���<�f�m�/'�ܥ��I�ې�A��-!�^��eW�����.:�h��:�����*Ns���}@�;�d`H����X�O{��YCʐ�vg3l	�;;���Z�ׄ��n	CAd���4��
AN��/.����� JG"�ܸ�N�On/��!�E�b���}���� ���Ơx�ݧ�oTJӌbhЏ�8���@�d����t�,Xy�����F�.ܧ [�R"��w6��«��ۡG���1�PǊR���NXw��0~J��,�(P6<׮��FŨ�I�+䚗1G��g��ߩ�b��]{\������5x�#_�3R�lö
�$ZV2T���Cxtt/_���S���l29�R��)qM��)���f���K�y�a.�־�-�S۱��
;Ǳˢ�]���-`W�1��R˶�IzQw�!�yG�kd
s��*�X�Q�;~��F��R�V�·ud���p�I��:������hDlD�q�b�w��z�)E�&��)FP x�ʰ��@�o$����R��d�L�*���e�!���!F~e0�Ŷe�&��4�A�C\�GX���E�\��6�"s�H�	ך��䇂rG/^a8��Q_d����JZA1�AJC�bm�g�4,�)A��[�m���?��0�ߥ>$��#E7�G\�&��gm<C3U����h8g�#�oG���@`�]E�����_�S:�S�]�Ҭ�_yS��ϊ[�B�X�B����I1u�R��<%�4����Ҁ���]!�.��d��\��b�^L�I���5�-��{I�C �v%\�5�R�E��s捿L��k�on����I�l��2��I��
�rVe�����b+��Z��+3���JG�\��Ô��]�q�Y3��N���E6�,���0���m��J���J�ڪ�Q���t���J"�@k��Q&"�>5r���nCAo\c��¬�
�)�3��5J��T�$� ,yq$�w�Q&��\����g��ô��2�	������,�R���ѧdLG)�h� ���K��$�58�<Fk������3ɡ���@���~��?(e���u� v�CO�'l7���d1Z#{���*���m���Ĕ<&f[=�:�/I�	^�����b�d��M�eQ������3 �,MS���#p'#���A_�O���QS_ H�%��̓*�7��.R�sk�����j(h/Q�>f�Ȅ/��O��9ʑ�}'x@�r��Jۏ7Z��=}ׂ(�ȿ�Q��c�ϔ"Fio�a���ܯ�"ġ��6ZfN��P�-�F��,Wv��k�F%4���Y�l٥��u��� Y��Q����j�]��{ s_{ɸ��x��0#dw���4�$�|?������jo�:>yOq�@���'�vn�B���PDd�rE�Q�5���gΩ)���]|#�
���s��,�:%�06��	A1�x�R�uZ6�@]���]Ā�D2����<��������������^`/l���ǫm5��Fx�| b]�x�n?����u�;��Pw�gZu8�HT���*���î��P�����)7�rL[����y઻��x��i���;�
0 �6�/���C(6Q�xD��O	�'0�P�54d&J�џ�'��e���;8���1OV�����{D�<���nAv:J���y�1�ңn�D'�N)>����W��S	�x'Π��QEڵ����?�1R�E���Țg��1��;��h�-��A�������:�@����S�H�����sP4e�z[2��y��svi{����A�A+$`�w�1˝v@9��C�lE��\}O������L����ͪ�� !V�!�_X����i^$\��Ŭ��z�Yq�4��<V�N4������_9O��^x�e�T�����8|>�z��Rs�B�_Ԝ�b��ť��k,��;%��H��Z?U��0�9���H�ۃ�����s�*J�j̖�eڮ~�ƴ#ͷ�D���G�Io�D�o����&�D.���M	�T��4�u��J�� N2i��PFA�r�[������Bh��+y2vN��<�Gwֆ��/��6I"��p��!�$���ǅ%�wY��uYQs7��0�!L҃JW������K6����|�Z�Fx��"�3<����}\�Kkn?P�lL�͔B��J@���vލG0p�S̆cxR��HxVjL�+��i
�0w�fe1���4 $J�ie�{;�D�.����h�HL_z�_pbxB���_U�
D����mQ���oKܩ^O+�Q���� 9_�>h0��z��Y�=z�tf�$ą�t�܍u
X4������#Qj�*�@`벸;�'��|�����p���X�k�U�ς�l,�y�����;e0.�Wvu����dT��vh���e�@�7�u�x��F����QWy�;�1��QF编kZ����!� �	H7(9�1���ǈ�@r���X��s�	Yo�"�-H��"�`���qC\�u�OE�E`��	�_mH��z�=غR�ų��]�� ^� }�\Z�-�W��ꦼs�������U��B�7D}\���^f�v."4�%�+5�k�<ϣ����? Sw�}\�QWץ��s]E)�"�\�ǒ\i`vv�|��J^��9b�Č�����{`ܫ�*���
B�A�Hf�̈8��0��Ȫ��~"S�U��O���9�p�?�F%����7��-6ϐ�^4`|�w��� �U��K��o$+zsbCNCi��nS.8a��H�e:���S��r��`R�
���^�b�Dh��٣]��FAc{�����*�lB��6�Yܮ�y<d�+,0^� ��4�fx΍BDFl%�z�k��"zN��ž>�,���]�㋻D"����g�|��
�·G��]����0���|p�TN���3���0�A=�o}�?_�5�570�)��u���4 �k�`�R�f����Z���֍\(��F��3�d��C�����Fo���,&uH�"��uf5@N����e'ơ�HO3l?��"�(�X�:$G�3ݵ��(��^�q2.�ns�{%�,
�\F��b�8��{`y�Q����n,���ϱ3��6v�X�
	�&���1ܠ7)%��ۨ�L$��EVi<ZH�{��q�B%�w��ޮ�%�±��e[ <Z�_ƤIT�ۧ�3�J"U(��8g��Å�v>��0�bn�5ʆ���J����11�ذ0��ݣ�rji���c5����t�;k\��[j�(ͪ<���(�B�� E�N���Y'۵4j�Q��5���@u= %�p.�Mt2a���Ӵ9b'�O�LJ&��F�~���YT��Ș�:��6a �����:q=�����*@r/�tG�䢕:�0�u �`��k��������R~��VL�P��i(���PHsdI���h��N̪�U݀���K���0��;�Ď��#��a��wF+����.�5���ɉ�B�A �̸��^���h�($����s���	G�� �P��ո��9��W�N��Î*C��F�������I������?\MHh���ÑCa�dqhb��sl����vV��ѱ��R����jb�������$��s��Nr@4�둗4���}]�r8��}�k �)���ؑ�G1{)L�l�z��,����'��@�b]h�H����<��&2�_R����hImz�oM����ՙ&�aK��~��;LI+hn� .4��!�8X[�o 8�6G�1��F�ҏ�aО{�y���|'�O�������v���=��!��������:%d�,_�C��,�Qʉ�3.���G@���خ0�Q�,��N?����3X��*�s��������e�ݐFF5��1�IO~iq�:�@�fX�	�ǀ�:7�Sӟ*�}(�?�k��}pr(�fŢ�\\��\��	$���Ɯpb��6d#3~Rs��� �?bk��!�\b}�&�3W��ݧ4�A��1@�'�a�M�,��t	�"��w�`�}�w�?t���^���ی��ñ^H ��5�v7��)�A�5!�Y�Կ0��)uV���W�Q_������D�M��ܮ��sާ`�Z�����&�^I�{�-;�J�eڦ]�و�,��a����}ϙ�R7�6�%�X�]��b��Q57�� qX�LY��Q�\I2r&��v�=-}>�8)���,���2�s�UEֈ��E0��V�aс�:۔ye����<�M�5/��",<���- 5k�]?��D�(�K���P�@[�9q3 �zM�����lk� �Ņ��ժ�b�zw[jC�X����[�{6����"��iR�+�ͷy�E�ȠafD8(XC�
h�f
����,m�kv��:Z��U�zY���8�K���Ř �����"Nv7������+5�я�)
�����T��?��M�7[�/
�X�%�62V�t��	�B�Q��~�����hBO}���4_�t�^�+�$ѥ������&e!��VȦƩ�������G'��D�����w
�7��7l�)V
�[����vY��r��K��;s�U	��ζ�r۩�͇m��k�����5�Ѧ�/D��(B#�z3�?\Tf��`�% T�
߾�l�����	%^��'�f���nM��#�a	¡ aNL]^+*=<����n��H��K�(>�"��ҏ��7<�H�g�ʨn��i�jȚ��ء���F��p�<�H� ��Dy�<�\=�V�7Cɕ8B��M�]������ԟ�X7A�HW�z�}�[�@^�)��*Ǝϊy�04y�$ї���橻�x�?��T���<�������l�Q7jP Y^�bw˧x�h�)��W�\��1^+�Q�|7�s��t/];$"~ڍ�AQ*<�z���9w�������҃�?�l��v}����U���t���u�`m�b��7��ӾAR�@\���.�Ih&���V�_�FLz�ᡝ=IC���o�$(�ftjUbo���K8��t�:{sx��"��i��>���oMx�D���g�JV�����d���c��c���t�?r�&�I�;;�)�
�W�-��ׯ~g鏕��9h	qo�f�8���f�4�Q��.��*��A�\���)�d����s�%s�h���u�8���q�=\t�XnGB�<+�� q�C��5��4�\7^p�O�*Y�����u���]�j�z̄ 7|��I��X�����/��'�FSa�l��Y��~��k��C�dQ�Z�+��Ʉ�w����I�D�����{���QB�����A/�����|F�Z��*.N�D@_��� 6�5�����K���*w��堣���"4Oa��F��p�M)�^����N�u�I��b�+�X���Q9�0.Cl~��H*�03�IM4��κD����CD&21���{"�f~�ġs�N+�/��pޒ�R�/4$��a��R�<^=����g��`����t��Z���}n�#����G��I�!u��JV}�H�����#T,�v΀�6���A�.�c�|�g��@��IJ
�U՜q����y��xԧ��R>����K��1<��]p�%��1i��t�|�����d5��{H}��x*j~ �����lY�<��Mj���2��+JɾZ�Nna���똩�Ƴ�v'��o�Vˑ����)��H��k;�{��2x��=��%����������]돯NI\����OD�i���E*�V�4ᷝ�aL)S����~�p�c=�hZG���ݜ�\������S'�/���2��@S���B�K��
z�^�����J(C�S�˟6vE43n����O 4 �ժ�%A��"��]_|��+��V�_����/�d��N����g÷3W�Tw=�����Y^���DG�gw���kP)�C|�~��ݹ�r�A?� �O����@��3&�=GG�e4��4�'���^ko0�xxy��&-��xr��{�+~�N������B�V����Ⱦ &9��!��	2���N�Z��h
b\L��҅!F����kF�~Ƣ��"�e�� �H�%e�������4P:�,l\�ab�#��)�_`i�ʑ���@1+��҄ޮ�o	��<E��Z��u�tA=�S�0MnB�Օ5�Uo��Ai}��,����ICo���K�k+�Z֥6���W����MZ�u�`(�k(���0�yε��Zu���Њ��\��s6� N^J �,�d	ɞ�a��&����S�ǧww�f}*KQ�oCݵGNB_s��9p,�K�j���Le,w�v��"��y�٫a��7,�����}��,��Z ~�]ȍ���|	����t��)l`�)o6M�x~
Ҧd��wg�b8FT���m(m�a>�g��_�$�R��8�z�2�V�&u�O;5R������c��@��C;tA<�7*�X�3ǀ��D��	�}��Z�.��c,U��{�Ѩ<�����ˏ4i����1"Kt�����ES�wHF���h�ae<� �0�w�4���X�,_�$r�
�5�.�Q���Qs�@U�6��*yrۚ&��dO�R	�J.W\�"F�%�� ��GP�Ro��R&�����%��?���r��(cueE߀��D��ǉz�Y���- sG�H���e�Ȓ���#ܔ"$`Mf5Z���'�Zgs��v:����a��	ӧi�]��MB�T�W�Tq��� �(�
\9�A!M*7���k�@��K�����%j�I�D�i�U��U��͘��9I��#y�ְj��Y��~e�&�o�����g��Vu�Ш��O�6Jj8�!,�(r�ůBj����0��*�$��aO�D( �h�&���s��j�
�����E�.4�EFW�	�d�B�_�A��/>S�L���F��Z-���P�5	l�y��$w��B�yY_�	����bsxՈЕ�ͧ%�/�@�:Iir�D���$��#�H�Q���<�ş׵��ή/�"\7��J��|x�d�Πq�z��i G����\����'/��%@=�����y�T(�M�b��E=�E�Iv��..��eֆI=M�M2ݗT�S�h�ڤU�1ș �5a�qM�}��"n"r9��e�?U��h���*onVh�E�ĽE=���E՚ɠwT"�v'�CI����ύ�V��iMf�Ϫ	$	�p�����ns�q擓�汰\��Wl�i������B�`e����N��ݏ��tjB�q>#��ÛAD��H���6Z��wd��7E���Ca��*�G�=΃.���a�i;�v��x4�N�
Ŝe�Ӣ�iV�3'�N@�Dr�"eS����S���w X�%��뵔ٳ[=�zi�R*�	?���Ud)�G;��wŰ��I�VK�<&VI����ʲy�{;
<��U�ԫ�єM��W�m�K�$���&Hz��M(���[-tǤ��+�;��S�v�g�4E+n��o�ہa���{$9����91i����M�Ny-�f3$&Z�b"��؀i&�N~C�Hf�R��<�'��+�:cJ�@�`5�5Q���uc�F�^�HC[��+��VX�&��/��P�M�V`�9^�2����c5#�w)��jb��T�w��o�v�P�������o�>����p%tHYPI�,{��uQ�_+�W�i��vP�`:�������u�ξ�I�LkO�;8*�K���1Rѯ��J��&t?P� �8'��(��ٙ�qUu/��nHJ�B/3r�?�j�h��)��+��*�� q�]���ۘT)4.�F>��1�9$�d�p�2h�T������=�̓�[�(�R�JUa�6ӒD1�\*��qh���a�T`6	�8����Xh��<�?�Zֳ�"`�<�*�i���a�P�'�ދ�	����Ыo�<�M�Kuxvz�Ґ��=����+�1;�}p	~Tg�{��^��w�V'U�#g���e���X���|�$��T���[r[�g���eBx3|ŬN�b���%��LJRh��x��+��MY�X?-T��&�˔ԍ<�:�?���c�yP����n�'iBE�1�>
.���OZ����J��g ��Iͧ�o|K\�1[�M�
QjnV'�����t2�>�l�;Nn`�!9?_�\��L\~��l�ۣj����;�|� Y3a!=����\d4,�.��7K�2$WT��q�~�xwFpW�����[�ygF��Iu��
	@̜F��pD�U��pQ\�ζ�S�^wά�Jd�A �����J���o��βms�5��9�*ӵj��m��l�X��b瓦'%̈́j�I���!��V{��!�cF��y�wr؁���nF��ɖG1d�#<�,�8mk�6?��?�d�zM��`�v�]���3T�h}z�}ݾ���P�3�@�R�D������S��_Β��Om`�;0B>*��/������|��� ��}��c�ӰȺ��F�5�Iꋯ�e�:�2[5&.*�����sF?����x�)��D~�t�}�T���ۀ���h%v��P�q�ȴq>�*JN���r!_�9��X��7�Wf��o�q�g���J`1v��pe�x����o*j�:�tަ��Ã^+s�I�#��9Z^n_��b��6H'wJR�YA�6�����AJ��"d��6W7�����K��=�8�?��f��U�w����OW}�h�S[ޅ���:�`�~^Ҧ�*�P8�߿�3ScTK�26���>J�ql�+S8,�q�E�4m�/�Z�Q��~�����́�Mpپ(����M7N���M�mY:���<�7\�[�F=ߥX�s<؇���劑�{�Ľ�q�Ff|@`���������^��B��Wx� |�X����j'PlY��ϼ�%�E�W
^ԑ�#���3�p��l�?PK� /��^�2��h[k����ce."�8���p(��JO�̿�l�4�MMav5�%�F�8'�|cs��������rTs�?�-����|��:�mI�؃�_�E�т�ѱ�bf�4Փ]�	�f��B��U4tn��{{7E���<	���Ҁl:3��E&�DG�$����#j���r�{:�Ք�8d����Ɓ2=�����J��,+��[(��!}aT˩����{[��ǂ3�ㆬdJ��7���?̌�l�����S�5؛��H��{�L�[�zY#5�w�V�����Q�r�������Hg�QZ���vJ%�X�Bߛ�8A ���,��\u�����"����hs�����:z����~xR[��$4��-u߅��u۟E���CQ�}���������D��۬��,O�����elA��·5G��M���\�ͦ}�h������4A2�rw ���$�38"F8�QO�n��0����ƺ� 2�L^����H��6��d�Wcj,�o�[�(�Vp�l�2c�����Q�s�XB��3~S���������kh���P�}�^���ϼh�L�//j8�j7��3�.�sZO-�_�=�'sx=����uc8��\�x��zy&J�������ȹ�@�B&�������wʐ%���Q�K/YY4���>�Ϋ��ׯ����w�{/F�uL���nꙘ~��OC���O�Ǐ�&����o��#����K��� ���Q�e��Yp	�y��T�V�g'�q�]Wӫ��oo��-�������o���<R�N�|����QZ꼾c�׸?�����٫�!�2j���N�P|�]�In�l���..o�bT�ke����X�"N�Z	��!�ܿqҘ��@�_&G�c�+�HytlQ
�����v��!�����WsZ�Ƞyɱ*	U���n�5O��ک5=����o��4��P����Pq�1@x6�۹��m��5Z���Z�զg��r��F�kH]���1�Jl�/vY��釥:��a\����F�P�e���! �`�ƻ��S2�~��RC�V�P�tU�����w�byj4O�۾�}r�+Ȣq��y���_;�X�����@��E���kQ-R�k^u~slB��$���.�:܃��7/0_��;!Z�e���d�ϖ�5�צ�a��D��.��v�����ڹ�$=���YAx��D��e�0C$�߭�`��7C�t�7�Csc{�#�[�ϻX��J�;�����g �{ |u8n�/ؠ��N
c�7nq�a�� �߆Z9�$���>�k�Sq�c4{B���̊�Tpr����W�a� .�wL5ke4��|�J�\1��QP����n�R��]msEyJ���3r��gٌ�Y�B�Q;q:|�h�K�ŔN��C��wr�����r ��&��_w��`���<�����P�ϱ��i-	\2�8�d��KS���{���+
�m`�+�#̉�\G�<��>�j?�]w(� Ae��頒��툇��b`���͌�D���g�R�t q�4��3�8�g���ߺ���?V�0�����r��u<�Y ���������#�򆆐.�W'��{����:�`�ު�Ҥ�V�r���0�Nl�Rw��v?��%�29A�Gk�ލ�:\u,�6�j���!32��W��X���E�ꞌ�ݎǪ;-R�������Z��N���zr[h�w� Q���vf��C����e�lK�!�5�W���^�;�Πp����ZS�y-��U��A�q֡8/��1�,IП���x�%��9�XO��~�}å /�i�ԥ�<>l��9_��x��N5�3�X���HϚ�y��I��i8B�h���#~�T�Ǝ�:����K���$IOO�&�:Hr�,��;�|��&���*q�f���xZѿ��2#�G�p�M�0%�Ȃُ��3��@�l�+ҵ���D��Ar.y
l�!�^���1Q�8]��\/��c�n^uԲ24/���t�w^�Ya	�)�iq��p��(]v|��T�.�6(���T���� �y��� \��1����4\�%+ȥNk©M���0;�ti�^����h�a0�G(���XR�w�L�p��O�d(�/܍З�{���5���x�j�鏈i��h��dZv�G��	��M��c��,{���T��iT{���}�j�}����NޝHz�i�ɴ�� �w�(
�ɕz/-�O�z�Llߟ<_b��bboa��� F�h��#�@�O����y���4�0osĠ�Q?g�ꕔ�b
H�u�.���"�G�s�\��
� �Yȫ�����!�s�=bݧdeɦ�E8�D� ��zI�14�ǧ���EWbd��ґ���b�/!g�`��d���̵���;��`.\2Y�<��#�m.�C%��y�OóVWϯǗ�r~E^��e��`1��A�]�6�ا�t�x炛�x1�=��|x� t#5ĿF�3���B6E.</�N3����^(A��s���^l�w\U�z��R�2cD�a'~(w����;>:mk'���D$)\�Ɔ�CZj���V����/������G�&�&���7�)�W�n�����b��x;�s����7�Fo�_��<s�%(��^�:��P8c�B)4���[`��σ,�u�q�=����QB��9�H�ώd\:��T&\��9o�(��a�GG%U��䙂G�iaED����0S���;��j�Y�h~]���ͣ�⬧�֧C�E�H}��Ă����&6$u��_���Nu��^���n�?1>qt�N!���X����j0�I��je8�;��ҍ
|պ�o��ͮt	��ϚJ����Nt(����2WE��<��׭�e5T������G!a�ma�8Q��V�B:����@�J��_ȼ������&�8�=�f%{H�µ��>�k`����L��&���$-���"��c�C��&����x��,|}�oB�7z�|7�փ���U����BIU=̠|~#�[E/�wy�oo�~\"����`=����9���������;�'�%./�O�/XE�ȫ��W5�Ӂz�i��'g;i����-��Gֵ�V��>n��j��>�H�
!ǽ6QG\?��`�q ���Y]�><�h������^0�JV����<�޺�><�ffcd���ݨ�$�e�NSH/�2��$`'�x�5�3���A�7ſ��ڏryMmV��,R�� �!V��t����>X0%Ԃ*�^��ћ2�U����/����Z�q�յ���	�,��#���@R�A���H�R%�?�B��m�ԋ.�OM]������6)�&��P��T����rY���ϋXu��<�k����.���t��G���݌"��[�i^��{j?�ѭG��t���QR*1�v����N���y�#I��>X���9���v$�C�L�����Rt0����㣭s��X@nVXOzR�Ǐ�$�����hZ����� �zk�X/n�]P��+L
CZ{ާN�f��w�g_�ġ��EM�$`#�Gj�M�+�B�ׯ�T&�џ������K���'��r�S�Ԟ~{Q���,��h�k��ޟ�!ܿ|���e"P3��4�``D�z�M�0h��AA|{[|��=6l;��az�,��.�4�ipc�n�F�
As���b]�Ex"��?���T ��e����/���T�����oȚ�FF�tl[�g�+:L��8s4��d}������`�S�_|��i����	Kt�?�t�<Yr�![�U����o�ג��i��y��jD�8S�,���)>*�0PA;��,d�d4|N��L�h��`wx�����E�KZ��qSf�1���Dk_LPo8�f_55�#�D0:5�'zJ��P�J�(*"U;���s������ۿ&4�ߑ�{ɭC�Fzd4���5b�ā��m+�� ��I����>�b�{�ɽw�ܟ�+b�e�A��q;�+����-���|= �z9kb5�P_F(���p��;CK�%yM�� <x���y�ō��M�Kv7���9� ��s����V��,���de
�y�a����t���Z#w�\���X��Rǀ��Eb.�"�H��.�Q��;�� ���Y��٨�"pc��X������S�θp�<v�A5�*���0y��O����I(Mp��O#b#gM���}�,V�"���ػ�������@GV���G�4�WE����	�D��Jfw#]{��(�i}�U�6�e�N5s,B�`�j՚`j�\���<Y�&t��5��nε���ȵJ�C� =�L:��#^vkk��޴�ya9�:j���~��c^��]� �3G�KT���������z�$h%��T�D��D�9��g-�I8E��n���/�@�RMu��%��W�4uٹ�0^Y����&���C�
b��$��r&���#�\.��Q��c���_1�P��������/�||J
����$X������Eއ|w�O��]�SS��3�&������1�[�R��N���H,��݌M<�� ����X�N�/�<R� 9�'fKPS;,���%�I��B"Ռx�s# �8���y���ݧ�e��?�G�ܖ�¾�D�v^C#���#�A���&������+�dd]h�^��Z���X���,�EVe��{N6 ��E}���v� >,5��G2��N`QT"x�kh�;�.����ei�
���k��|�F���|@J\y�g��ۙ+��J�jH"Sw�𬠏Hߚ�TE�VT�nѱ�}��q~A�_�6�q>���OT���$ʬ�4�B��L�@S�S7{KӇ��FtZQ���5Zj���$��g�#q}?��(��o.+^)6Az�����a�� @ɡ��qz�A	l�|.wO;���%���wq�^��(����>j5����H��mdb�c�?Vul��p��br��q�}׌�O�Lh��EWM�`)�p灉��`���m�͝�rR}�C���]x��.�;ۋz����y�&:����OO ).eU�5�f��hl�IYq.Ѱ�����3����E�9�s��9l�t!�=�u������h]5\�9^��7�Z8k���Z	SM�j��8�B����x�����1��=��fz���I揠YQ�g��4���u��;���5��OK�ǘ�|é��+��ѯ3���������2��r�B�<w�������v���`C;a+8E�qs{�Rtv��6�)A�o�H���%62z5&�T��4�nj/�OJn�O>֒����G�Z,? a�oR�n��"U:od����q��D����j;��C6���Dp/��9��KXw0#i���]�3^!o��&��E[;�:H��y�E�9 �L  3��ނ�&�"�M{ы��Sr��:�t �g$q�D�z;x%=�;Sr��ZY=�Q�&��0�u|qSRY���M�g���(V����B	�Z�Z�@K��	�^�pc��ab�߆D�ṝN�����R���Xy�`�����᭄�A~kb�B�@n'�#��'d�`���e��.\ ۷>��=?Is�B�z���\]���	e�Ѧ�ӟx��+�g�N���8�{I�z�q,�
�Ս6��j�؟�To�!T���-�0S1�~���ۓ�QMBnBoNɀ߄�t70���T���w����=�&7W�T��Dn��$�)��9�$�,ף�F��P��ǵ5����x�$�uz�L��i��þ�Qe.Pz_����'E^��`�<<�U�C�8ZuLs��X,=��s@�j�*���>"`P0�@#���>�N�����+a��q�T�>��O��Ei�wRG)���e�x�i�6%J9�d��ܚ�}M-\���.�c�R8���X��� L��=�$A��o�
#��v3>|�+Ok ��]"��\{�Ҽ2 -�a�	�aS�O�]Dy�KD��+k���VNv�L��vw�W�ROo��Ws�K����av�}G��2	���ooI���kN�L����[Eܟ�n/�J?<0+,7V�lu��3
;�:�"t>�?Yݪz�KT��I�������IJ��=1�	�k<_׽S1�۱���uV9��u��y^�b{��'���BZ�K���VE�a�����C�>4��F��k��ظ��u�Ջ��Q=@2�' ����$������2w�Þ鋕���<cc|���0���� ��y�Z���p��o��&wyz�J����Hh��m��e)��w���Yx�ޟ��S��'�����̈��.�,v�#��/�������32r�e��2�4�FG�߾Fvt�f�~<�� O���qӺv�Hb4�*�C����=Bi��:��������6]�a��F_@�<�ۂ3G�[��	�p,4���Oz�8��|���\��U�wX�$���Qm�Z��k@B�ec�^�3�]s�x�һ}SFd@� �3_L`��N�Z��&C��@��}�Z�x�Rk������(�6��j�=eTN{s�Dƛ�!����5�P2�����+$#_f���2�+�{��##5�/�*JB�*�
6�N�1��2
6�ߴ��p+��r�7�a���}�Qد�އ*�gF�m�sc�ʗ��,1d +EK,�f�������}8�R�h	OH_/Ev����UI#}p-����c��:c�vA���$��6h7r b}��bw�Pj�O�IW��ё�`�� Z�[��g������r��WyJ�R�x���;\�o���'5���G���i/�,-�v��c�y˪�����L��p��˰MZV#љ�M
6�o��&�e�������z�������i[��l��k��H��W|�uy%`tj��.����N�z����������4,�u�a��O�j%Y�%/e�<���R|���[XN�ɠ�#��lwgF�@`���l�n.�ߍ@ (�Kn��zD쌗��������}�O��?��;�xN��fW�/����R�j����9�ܠ`R惻"��|ѕC/S����˛�]L:�h��� �,�zᑜ~=���F�я�?2P�c�}	-��:@�N@�"��p�%3�˥�4�����ɍ�4��=��&��t奜nN��+!��I���-���i(�R��g?mi�"�va>���<��KΈqd��|��"��= �W�r���Vq��@um:�q^li��}�B�'�kzC�����Yx����a�&�1U7��ehc`������z�wg��Ր�_>
�n��`����DZ���r�xDd'�����Qgj��H8J�
7R �x��m;�'*�
�W���k�˗�.I�h�%�,�ê�y���̇X�~R��ٗ���2�[�wX���UmO��������z�S�:��֍NVp�Y��?��Uy�3ߞZA��D����PF�N�G��K�%��x�<�����\����캰�L�$��F��%/��^��+i1�*a����x�d�L��m=�w�l1˞�M9�f<W�@��]*��
�k���ϢM��Nc�ض>�:�g�2�X�Z���� _�N�,�g;o��ʁ�G]c<m�!����^��[:����'����rc`�R��N�~�i{�\����h��_E�D^<��w���;�7ѵӀ/C�u̶��wif�=�(?��L1bUk�5�ŭ+I��P�^��?��,���|�Cn�)�#e��_X�)�BO�GձX�r6�������8��ù���>��hG�f�x�&���.�$6��w\-m��L\�v&~V��I���I+B�������J�m�B�=Y�m��y֟kw�Nhp���@v4���ͱ/c�1�;�I�!�o[Ǉ
-7]���A�����_S7�h�v��-�yN�V���w8��a�,�L<)C�l��a8�}�ә��[��iB6��Ӝe��Nl	�����m��.���0Q	F
�6����)��� N�l9Q���������GT%�Q�����n��\x�?ߝ�+d�҇��z�}'�BFOpH	
�A���q�A�0�nq�{'x�D��r�����ևol� r����X	�b�X���]/�OR+��8����(`��t��ۤ%�V�+����_z�yϚ��Q6<���;���<U�wQ������T�?ρ8�4�$����P����yX��(_B���x�J���]Ye�T�����o�7�.E�� ������[)�G�2�h=o@t���Ľ�Uko�O��>�߇Q�=Q;�����|1s}������1���Ѩ������ O[�@E6��_��W�F�8HV#!�no0��Ĩ�;#��AEDlІQt�����,�	�"5�3�D���L��pig����'@�_t�&��~hNE-N$��Im�CڮW����}4��իC�,s��G��>��\�A]%)]����̘��s{��Mت���#Lb�7�W&�Y��cqltk�(1�������񨣗]���"�z@@c_` \��+�@H�:�rqG''$HwQ$Ȣ°�G�DI��ɇrGu��ӹ��*�R!���"x$�F�T��b��b��Y���K7&�ܩD�x�sFR��l.�$�%x ���+ǩ��O`���e'���-��S�/�ǋ�!��|�)�/e	�T����"'����
�;a�gZ ��Ja����RHZ"�OxUb��{*M�n�����?��8�V.^����

�@�ֹ��߻�V�i.�*M�:2�c�<���i��t���zf�	�������X�wqe��k[�dA]�C���3�CgoG��rNX(�U��`���5�y�������e�%��Al,�'�(-tl5!���NTu,��0�[��!���;؀�}7M=M�o�_W���zT�����2^u�ņ�ڡ���.��5pso�F��{��6�X1��n�W���$���Te7��P\{0���+�Ʒ��ue�."���m�X�
��ek���b�B�l#_����b��:�G<cق�]%�ױ	�Љ�^y��֚��8��'�[�Hp"<��kyf���n�PgUG)l�KuF�X�?&R�� �zEzL J�+�{����0<Ί�U��!r7�����p]1A�b�Ƙo�_Z�V/��V
"n�����
�S���M`}�z�B�t�0����]�۸�õ<�d�T�XBL���3��ûipڗp�P��Dl]�a��?
tZE2kHR�Ov��3�܇G�dx��
���v�Z	�{��]|,~�HO���@�[���)�wb�)�w�?�PG)�kN��S�(i�]��&(��>���0�?�Fvk��3&�o4
'm�jN�{Q��9�fKW%�y3|m!t9��Xh�G��o69X�}ͭ��6*
��hL�ҷ�&��}����E�
C2ƭ�8���Am�)+O*�~����w��h1�d����>aN^�`�Y�����L|}�� +^u���˾^���O��j�+� tÖ��>�1>$?U���6f˱F�	]&�h
��ΒO���|�ߕ��8x�`�s;�u^�#�"�n!�wڤTuPz}^���e�]9�t	e|P ����D�W���e̷J������V�Vny���<����-���d���Q�TL��/��Nd���D��~XF(u�F��4��xĘ���[t������ �-�C���@��}>ˁ�����$�6����}��"݁�0���q��n<�1:��S8C��@s
���Ξ�HQ����#P?%�������IP2kJf��@��bS�~��D�.����Z�a6�)x/۪�C��Q��
2D��&Rs��L��F��g�1�''�C�?���O��/�M�jX�G��Sm��2��JcDj��q�"Yݬ�m��Fg=��?���Z�����Y,�ۗ�B�8HJ�eƪ�Wd[����}a��qS����l$+J���-W�D>h>? m��P�k�^��<��].���%��4�Y�1��m�ix[oqo;I�Mq�۾���Z-�ʯ�I�5�C����2ޠ�o���x��
V���a�
��[&��=�zϊ;*��*>��D�o��&��C�Y�']��[��?�p�r�MU������b�,DR9|���CD��Ъ֫����H�\���X��E�^�@�%8�r��B�6l}K]S
���妼�$���F�s'����Ӟ.�Y`=��}�Fgf$9��>��t�9�� �E�+���9�Z8��jS�����z��<�VlZ�w&eI9Hgi�t硼4��k��_ƦS�Y�V�.L�w��+cq�����H��V3�ܩ�5a��/xA��E]�fAA�k�[' `�P��W@��r�IDyKe��[ʴ��̎�%=�'m&�E{l�p���_�����7cJ���u쒰�[%��I�
c�S�I�����!�6�ܒ?Ar���b$�h�#��;�lO�Ʒj��n���4�#Jg����;��v��%[�@Y�~��JK���7$�]z`�<"l�ԛq;��g���ް[r�T�|�?;IK�"��H&��󗕚N�,A�M���u?	Q�,��� x��C\x
s�h{A�}�\
�""�ѐ"�7l�iO�'�bP;crP����`��Tf:������pY}?����6�%tr���"���0��� ���g��Ⱦ��Ҁ� ���r�{!�:�5�هj<���l�6��1��+]�`��G��i�0�Z��K��b�g����O�7Z.�N���z@wQڌxSB}vf^Ah?�����q��T&;x&C�E*��V~'0��ԙL �^�9A���\��xD���e0/��[�x{W��]��"�Y�"n���}���`n�&uYT�Y���$�Ȇ�A��Z�ا����H���,թ�p���Q!�Ý�B�33��]�e���O��u:�OZ��e0	)g�uL3h[A%n�3\ tvD?��(��E~͑D�ʒ2��Ё�I��V�R]��Uեq1�(�۾��aۧk�<GC�ma�lU����*�v*��/؞=�5����F��~���6����=�����b�;��Hou�n�3��V����v�b4��ƿJ���+9�1l�m!2�s��)b��*���o7��`��7k������m���U�lu�bx�� � ��<��&%�'�&��4qKK����0�A�����݋�B�9k��.��{X5���h��oU��#+=w����L�6'��mlw�Z�û}9�`��Y�Wm�u��T�q|S�%��l�΍ �B{����`��Z�/�o�GN����j��m�SX�I[�h�>�s��8jc8<��+�6����n��i�Z�i��}�2H���¿����T�h�d'B��a��y���]K����z����򺽾�CF�hR�@��f�ы��OE�@��R0��Q>�0e#nA�c���Y�I�$X�M����~H�=���</*$�����㰪�nS4�p\�Г��'4��:��G�q�ʑ���mRk}b���﹂��<�v�$�i�լNa�T��s�j0�V��E�~,s`�w��kY�e�Uod���!��?��o!+�+��Q�q�撷�ى�nu\��-����Lq�˶c(��xw�b��zA?ꌹ}T�񝯛�9i�B�2X}�K<�c���+�k�o��y��O�xV�v��Ê�)�jx�.�U�����0��Og.)��m���>����l��-}c�o�B ���$|�,�w�+^xjֱ�����K]:Y ����Puő�Qm��
x�md�j	���T����@Sz�]M���h��<�Ezq23gZ�:���]Թ�}������G�1Bd��p��N-{�!;�:/48-�^�ݖ���E�6ͻ�m)E� ���"��KKh��A�;�-
᪨Y�q�:�k\z��Y��TY�/��IOūH2Mڻ���b�1rk�w��(0ߏ�=t��F��S�)&C���BP���9��b�%~f�P����b�:|�{��tE.�̙5"Nk�a}��&��Mh��_>s��,��4��IN���ع�q�F�Y�*��*�bܑ���C
B7�}��xk-�ǉ��a�i��>�8slԯ�'�C��g��V��ƕo��~����]�ƍK���#m,}9[5��ANM�]��b�]�o)���)<�C+&ϴ���z\5Ε�4����>��K��ڤ�B��.�ct�Ӕ�9Rmʎw������ԝ+2���ٔ�D"�\�/�]��Z;�8�B��7_�f�����*�$C���CC����f���EZ�˗tw���r��Q�Q���k?�%�&�"j�s�����h-�7'��h�P�&���I,���d.��&^*�j��7���(�)�q����~9sT�dc%Ca��m��=gL\}��A����3�⿍����C§�,���ͺ�M����י]6<�y�xJ6��j��bU;R�}��\*�v,~7��0Cx�
.�"d�@����嗚#2*��qB�)R�;Ʊ)��"�������3�$TL���"q+��ht�L�#� |%!��F3��?w��aB=D���Z�3`�+�?��Z�L"�gҺ����l�g�E��<�&(��}�i����L�<���Su��,����t<�z����x�+N�J���h(��I��HV�����+�&���F���)]��d��F�*�j6�nZ�L{U�{?����&�#9�U��E0��q��n�C�n��f��F
�疂iE
:.�jԪ�ǦaOl��Xm}@�Z�*|����H�}Z}uf|pl*ɐ<�H�leRN���߁bҌ������e:�?�)�)gj��1"&/��8R�&a&aJg�"��*��0
���-_���VB���H���ɕ�-I�/~�7�N���,=:/�*٦3�)�$�Jz��8
.��=�9\�ϙJc���<J/)C� e����ϱ趭���Ul�)ZJ���_�]G̠5)��(pn�f�.��[�M��=�͐k�ߍP%eX�$i{g�k��)���'H-)���o��r|��^O��C+U��_[ �bҶV
�\	��_� �晏ǳ��K�����/d�����9��:h��ع�mն��\�����x.��u1k>�uO Ns�Y_o�q7N�i�BS�n"�ǥ?� R.�Y� ��אÐ��C�W<���K�B���-����X��9a6l/f�Y�-#��^��j�>,�9��dJ���Z=b&3=����bFչ����w�>-�ҽ.�ȧu��y�fͪ!�su�c��	�԰���1܍�-x6����Y�E[+��읝��s�`�7�}��"u��u��R#�]K�X �w�9s^r����hꗿ�A������	Ď;���N[{(�9�A�� 줸ɏ��l�a���	�j�� �r���4���-Hz[{�JXJX��E��	���lA+"��"�o�K���Gv��D]�Dz��P#1c�k��-�߻�HW�F�B\��>-�N�Aѣ7�����t� �� k 2�.9�>�y
;o [��~!��^z���~=b��z�w�F�R�m�H�*m_#@L�'�"u�&.&]��pwM�p7����WO��q��ټ;!(�F�'�Q��r_U��6��dccF�V�(��Nը<��
��[X�I����;)�~�@���,ĸ�F=+����c�d������ ���l����:㔜�k?$V��M���Z�Vr�Tp~�=���o��ڬ�=�Ja�
�7�TΣ�����_��(��L.�$�5 U�f�a��|/,D?8��8��Q�\��������5n���_�,!`d��j1��nX�>Aܤ|Tn�=e:���TBBt�P=�i�!�bk�X�4��q�g�vk7l>Oݳ9��D�gh�~XK�e�]���	���Чd��~�k� 
4���#�����Qv:<Z��[h�zU��Q��9�/�\��R����n�������ٺF�=Ɓ�x�#�95�F����][��ve=� Ԇ*���W�W(	?�cXNYc�������Y7s ���o�a2Dz"�%Q�G�N��@:�xS���7�f`�WB���)P?����j�*�9I"��j"� am%����8���P-��8q,�kC�S�Ɗ�}{�MٕR�������`�_~�q��	���1
j�QYV��	��T/?م*��ܤ��a���q9?M���:�9eۚ�)o�u>@�Ih�eܱI"����/A#���m ��OW:\.H-	���%3ǘܹo��~'y
���-"�-[�Ύ�B���3}`�P�4��� ��)֍���Xa�'/��3M��58�i��O��L��d��`ٛ*����w0:BE���n�(��.�e\�T
W���y�_�,� ���!�ʓ��e��W�m���rF7�V:�\�YoE769�+�q����B��?x_�S蝌�z�Am�Ӯc����`&��a�^z�2X����k����J�&�D�5��ɴ"N�N�3c����\\�9�6z�����p������gY�m���u8f�?���_g���oC��i|���9"�V�΅�Ι�U��ͅ�P���4L~���Z>����ڛv ���y%��R�������K���I��<�*��Ek��;<�]�۱�Q����>�����Q��CM?���������?������eZS}���kŊJ�?з�́�H�ƪ�m4[�j�E�ߴ=���J�h��ؤO-]���� 5�j���:+�D�u���K�b�s�B�#��*W�Yr�&��,~��o"��>0�ᵭ�������5,
lM�WJhA-{�x�� jw��
P�~j:�m#9Y��db��vd/�p3@u�8������x Ґ�`�������m��js]`j�Õ�;�mj�GM�mYv�S��ۅ?��blo��Y�7d�X�ן��h��:�@����ذ}�V�	Q9�l���RYu��VBᶲ����n_�@um�S��l����ļ �p\@���pi��J�xZ�J�I���RH#�W� ���N��08�":>�ň*�lzM��"���E�:u��_��$�l����̸�;�3�m���C�ص��]��y)@�ٳ�^|U[��O��#ǫ�gF)�=��ނp�}6c?���cZR5�P�4A�+�?~5����目~0�lE�Jp<܈�G�\2<|	�������:eU�|���o�!�N=G�:���"�pv�(V�sD1V�����̓�lp��f�	8!���5��#��ES+j
��h����t�����D�f���l`�I����Kc��iL�+5-�5����v��=̟�0��������M���D��<	8�W����MYH��/�HxŪ����d�ݖ���r�F��ᆶ�����a��� :��Ȫ%��aղ�1�8j)戉��N��Y�Wro�����O��xŒOF魠{�cR�
�T���)�Wq`��S\p�Ԃ~5BI��iŤ
�~ {ΟF�����<�B���jE��g�皹�'v{duW�%RB:ba�Xț�Y\x�ԅo�����B�m)�<�	�/��/��2 "�� �8�Vy�^��a3;4�1��+��hH�C=, �:�� =)N�@�R�迶.�`��(�,H!sRn�{߸��9���X�dP�^����x6��4�v~�ֲ�8�󞭕vK�-a��hTENz.wډ�Pg����GV��	<$~��8q�ҍP	�vD���GWʼY�F�y
�l��	1�*�����/�Y��/��Z9�҂��1�6�^SƚP��ٟQ�|W�hL�d]Vup������>�M��cC�w�΍�G�I12�?
�M��Gm����#&�4;�s9����~�ί��4�B�<�盰���[��-�ˋ��5�"�y�f�Q������ |t�"lX�u�kfj�b�,�9"5�?��>��*DVL�ǚ�K��1���w�m�0V���As9��tikX��m=cދ�J��{�0�n�1#4���Lh�;SΥ�h)׬{@� *[=��9f�k��2�8{����+��E���F*қ����g,����I���ŧ�(��Z����?X0�;��85�+�w�:�H �Ϛ%V�
�i`a�햫Q��;:-�3�N��ܔW87�݀ � ��LZ���ex�&WfLi/�5&i��ẑ (+w�����`�{�Ҧ�V��8�G6h��f��-���@��"J�z�pΩ��9�U�"�
L*����B�Zj�_*�nl�:���)��@L@�z��1�i�q��?���R�l������k�c%�pQث��Z����0S���D�+�i2`��*����sk�}�c�g?��u�V��/گX���)�q2��W[/�D�cq;	���i�됸`�Ry?)
m��	h�t]��vMvŊ��s�x�O�W��+��Q�}#�Wџ��u��<����[�w�gH	��`ՖM�c���bĽ�/�Z�� ����дq.3G�BH����-ּ�xY�mٿxW�r+l��!���/��X�S���/m&�=�r���V�b���Q�ߗpm8(q��Oם?�"�ꐳ�^���5��N9���=���B���&T�	J9�堶|\�f�s<��.+l�/�"�;`��}'��b P,���?�׈����z���3E̱�ZVF�Wz<U��sg�\M�����{S	�j��o�����UhV�u_�JAZ%.��#��t?ń�>RsYPh�dt�J�c����mL�М�0��'�t��u���@����uX��F�9s�yV���	���J�o]7�n��ŵ�K=��"��W�+5 ������0ZeV��XM^'(bKC�l�Le��C���Q�XlO�σ�![������#�k_�~0bNz��������M�?c�jcrn@P�e�S���
�}��[����{�j ^�L
L�7�8qۙ�M ��V�}�J�R�R��OS���`��z�W܀m�:\���ã�'Sΰ���-��2���ABF��թ��i"�,�;��w}t�q��[fͲ/^k���AW����O��D����LY� �^n"A�typ����E]+�*�T�__�ع�_<a�[�3Hd�bpB�c1��!���zX�E���&�z`3D(c��fxIa7�h�U�P����fw���
��,�������3jY���^�^�W�<���k(Hh#=�g%q�����蓓���q4�x���GʭT����)*�L�Ne�7���ɬ�ăJK����V�E4�գ�9�|&����s&���=�w��Q��J�`)�_����ƀ�m�1�4dv���J���6��2S�҉��0���3�1Ŧ*���0�˜�=�� HFֻ�FJH���T�j?U"��=�Y�m�h�z%̑����W�X�NZ�~����}�8�,�����>ZA�r�"�y�љ�C���L=%gE荫��=Xc�Ky0���rdM���ɒŊ����@����nwc|���z1M�������pj�*�g)������r&~Y���K9��G�}��ɂ�3��'�����Ȳ
�T\�0w�Oj�ɝ��o'��W���[ʷ&n!��0�"��l���)ԉ�8�Ԡ�P�F��꿫G{�:o�e�&���ǟ�Vc%��Ju���ߍ�-x�^w	�֔�H���W�LXB��j4�"����m�XQ!���&\��=��DG<�%S���oY�S�3W;ũ�aN^)��z�w˽�ⷧ랂�ЈSxl��U���A��!E��n��C�Q�٬�k�$|�l��p74G1�4�Ԍ���S,:㔴��E�O|�>�=�X�J���)�����,���s��;��R�뫂GH�'�r�xb2� V�K�	���5&@�M�4��(�&k��}�w^]�2n�:)�ti�4�_9�b���&���6'#v�I����@�,`dQ�������cr1Z�x�,�@٢Kw��R��J�g���ֺ���Хվ�}��>?!��a��A,;)$�����*�������?Ai��-u���n�*���W��KH��� �o�u`��φ�� D� u���Y��������{ g�L�ڡ�W�2M�W�_%�|>R:^H��O�J
�P�HK�YJ�%N�j���+;Jg�o�eu�w�g?�������I�G��^�������Y1~��{�z�`�����Qd��*��l�I���T}x��q�<���u��Sr�Y�C�_L���;q���]��cP��^��c���sO�ň�� �fړ��]�ͤ5"�(,�4���4�Q���O���3�KH�Olt�\|g��+����+D�!�iv�[���]{�p�ӆ����2�mmѴb��E�wF���^W�zx�es��U�G�#zʕ3b��Zn,41�D\/{7�ǚ �.�U�p ?7�4� ����P�7���9��]7_j��C��`�ʻ dW��vrx�Dnb�)�|�I�[wX��Ⱦ���ڥ���rr5F}2��b��,���v��,��h��0<A�N˪1z5b�޷e=Ӎ�"�1je�H`����3u��m˿>���y�#��Uo:�iCE��&���2��wC�3��D��?<�UIԅ�u�_#����n_q�y]�"��?<������?�(fo�u�������5z�>3�i��]�߼e�����nU�Q��}ʆ�Gٜ�oCe���s Ps��o��=W�mS���ޅWk�&E�^D Wv�$0J
���U_���hB]*_�����L���ş�ѻ���[2?e��D������n�������C���l,�>�<�p9z�ڭd����},{��1&�1����}~k"ą�Vj��
)��wEDb=�O{��w3�H.7 coL�Ûf�!�������19��P��o�z1s��O��3n[W��;�ڻ��|���(�F�|a^e�"1� E��Rݭ�I��]���e����i?le<�kyX#�IFc��
g�ք��7Q%#ŭWB�<��d/-<�5�:�F��'�6�g��}e�.L{'i��I�]h>z��X�@-�l��z]��󄛝u)�۳��/&H2�/k��by��O���gБ���=�����6U����"�d�GZ'	7��V�,;�y���#wqŵ��!J�v�c��$��pc@hT�J$�������J:���H��^�2o�GMS5O�i:q}%���.60�=�~�`���%�&8;�EV1����1��be�5 ��%*+�b �$�'��L;��W9���֞M����wT����*z�n�-���{	%��9,���s�y�I�Z?�a�a��}0���mn:�Wo�ᓷ��C;()EGl��i��<=�8�K�~{�&��]�K5N��j��d�%�F��	Η�u^���p���Q����'`��n
,�@4�;�x���΁�(yGܿ&�覕�Ү1�G��|�$�Z�ѡ����y��{	��n6��O������)�<\�D�>��W�����d��Q �3����;8P@d9P��t���(�#�����a�`zXZ%Wň������'�Dl����>��=uמ� ��T�m%e���c�"��R��%.��[{Ͳ�2od�GחD������=7%s��C��c�4JF\��OП�w���E��h���0<�6��N����*�%�/��zK~�Yk�2��'�}Q�讄/T��Ԏb��p��<��7n�\��45eTNd����j�����4y-9`V�G�,���5I�?���4Y��	�ǒsz�ش�o*L���ߡ���z�-���Υ�t9R�OH�M=�54�n�ɠ�s`g�Z��(m~פ�5�O��?���J�ϲ��Au"nI^�L�}N�����z�1U��zˢ?�&�D���PO~���u83�q��!$�5b��[�5�횤nlI!�@�n�g�B��C��?)� �?�eϵ�b�%�	{M��rYx�'���DpG�T̀�W�聐��b!J��'�ۖ�uG�f��z�%d� Z�\<��vq�ڥ����m[�Ir�-CC�AmS�2�a���c���wi͙E�SM�
ƀ ���41��Hܥ�j�2-����Vx�FbMK1|h��|k�9�/�k�Yݛچ����%rҬO�1=��68�E �0���~�ś
���rk�u<蘾�d�
�yry�Wz���$�(��g~#�D6Г鶞~6`�uX;���D6튋R�Hy�C�C�Yͨ�r���������	ǟ��#�\��\Xsrq�l�U�ұ%w��#��$�ֱ[w
��{Hw���[� ɠ:+�"t!��lV��/1��@�F�_�����Ћ+d������Ӌܟ��הK�ȆpG&�M,�Mw�Ǜ*0�O!u)!��gW�6/2=M>7��������3Xtea�һ2�Xy;?����p�ȡo�*s(��������Z!�֔5p��eG�zjۤ	vc���K@*@R)��B�p��#��I�=۲}�@ͩs6�����FS;J����������h�t�����!qA9�%����	;�I6�qS�i���>�yђ�+�O׹�+[��}�ԃ|m�o��B *v����@Z�d���7�v�	>�ߤ:;�:b���ī��.�ݙã�B�P�\��P�w��w�!���&�~�.����)��,��W��<asl�w�M,
�6���\lM���b)����O&���-��m�љ���kn'��3���4�j��`��i3����P����>�m��[ĉ�b��:��a&}U���e�z�-q�@��{�h�Up̓S����O��$F�Hmx���­�`�8Tgq�[i?K+�F�`����Mj��~�3�W]q|�\�v�9@=G��.h/O�=�/��������O��}As;�,$*�
��9��$����Lt:��FU��zT_k�,�nt'؛�kS��ӓ�9����J�X�hO���4 �,�V;l��}J|�\������=�ǯ$G>�2:�!b~�������nV��Kn��dׅ��?ZZ��Uu��uf(q�S�#nq�6w<���:��uA���>�:�'�����Z3Ǘ��#�{���V�Ҍ�_�Q���`4P֋�@���¯�7�
�R3>L���r��04K�C��hFw�l-�^C�,3��xv������$�0�@�Ed�>t��C����'�b���E	���I%�w�� D�L��:U�A(B���'Й=xB���%Ų��?Z]1�>�J��Ku�t�2�Aa�C0Q1�8&uG��0�;:��ؐ�P)�:m�t���uf�>��)v���tF}h��}��c.��"�k� 1��i�����N��t׀G �Лh��Qv�qz_�G�%��{M;
� J���>���_]��dVM?6�E�#P�=�k�`��[TZ��3�#�:^�6x	-��Hq��[��'c������Uj���l3�'�:OS�(�	 ���\�C4Y>�!h|&jC��j*#�
Ɠ��;�4B���Ƃo��t��Y���V_�I'��C����83w�9��`��b:B�z��:XT`��|8U�]٫W���<ɀ��Lv�]��m��C���J���s�_���.������	�K�-���E��FN�_($^�����#�S�L��v$�������k�o����Ԛ�e���Ԗ���ڃd����j��gQE������0Z���9�f��$UJp?,�}i�+m����CtL�CU ���n��~�8�2�@���`Bcv
pK��BC�n�V�SMB_}�u�;{��F����4���`��테"%U֮�kj5�GB�U����5�H�O��Į�IsgK���z5`à��Ļ`���yjf+z�!�"D�(��c�|�.�9�p����&
��D�LR�{��ς}�t��ʽL1�W��F�&��x�;:��F�Q� g��*l�(�uC�7f>&9R,H�	{E�5���J��]�GR�����[�rW[�8wq��v��E�đ�"� e�����^ٮF��T��/m
��Y"��wVO�T���s��ߘ�$�6�i/p�%�����1���U�%.�,�\�� ����ߦ���\P���5�b�syqs��wW��J��i�Կ?���AH.�������X<*�:��͙Ao5޴�`�ۿܝ
�9^z#�Ml]�\�,@ !�v�Ib�꘮��R����[��3�0�h-���wK�i�2\XU��wE�HR���M�C��(�%�%s�r�yr�4�Q|@Z�Wr|C����Q��}.��@��X��n��xx;�ofb��J�{�[K2B���3������HN٘��ۤ2B7D	&��G_� �Qu.�#��~'xo�A�2�p��[Vh�ŝ�4o�`�(k%J���K�˟"����I憆���Dz�7�SE�
X�j�p�s௪"K��),�]:�Z9A&笷�E}�B�����&�[ʫ{���������ڃ!
޶�q���?s���Y�8���,���:���Gq̌�턷^39SS��M���Ϟ����}__�Լ�[�It��S��0�r�f��v�Ԕ��NV>�|��͗�VD�^]��nyD!�!���j��~�F� ��}�C"͈��3�J��y3���!^@������h��z��M��y�Z�R�a�ɗ�����U5�� �����\��YDr�D�,(�߉�����y����|+3�l�#u�-����#�*��=��C�
О�`[q7��(�8����ȳ�&�j�a�
.qر�{��-��i�n.'��4�3���D��,$z��NIi=�V'E+:XNR������f�y�)W����o�K)�/h��]z��c	z~���e!Ϥ���<�CZ��{ m��� 6��$=�{�҂f� w�0[i[�̳�kY$˴!��ǔcD^��������D4�Rti
�nC7A��n�������徢�'4��91���M�:�F����v�/ZQm�a%�.~YC7ܞ:<!���B&n����\0�����d����������f�����$ͱ޺*��ۆ�.�B/�����2:w��ї�J�{�Q&P��83�|V��p��e���f�hȽ[����V��s6�LZ3�C��t�)kS��7��^��I��2�����)��;U�ީ1e�ҍUl�{�{���*,��Jѱ3y��y���w�=P���j.�7�;3[}�)�����hE�и�<��u�b�,�tf�sr��f�Zh�v�
��ވZw��A��#@�IG���Z5rK�^ԯsG�vnIAAu"�r�+D�/�5�t�*\��T�P.3�]Ɂ�o�K��P\b-�X0i��p��,P��)��?�0k¸>��"���k��*�Σ�G��1II��_i\�n/^���M��9KұR �[d�Q l�:�?��MرL/�~��>��]�$r�t�ͅ=�@ǵ����4��<{�ۯ@U�k,<9�Л��W�Sv�[)�(oV&.�޹	Y�B��Xة ct��P��c�ʯ�}��C:$kj
:m*���׏ ��O=��* �H+��esl�5@<��
�A�����쒀���n�DU�r����������?Z����"R��d�Bgͫ&�~�����_i�Qim2_DN���VF��IU���C��D/V�޵�&R��iZ6<�{��oK��P�Gm�)g�A�N:��)��K~���
����&Y����p�2��dP�6 �/�L��Ry����T���yV&$+�F/¥�n�!f��h�#�dU�g��leԲe�=�`>`(��]F��2#�-���]�g��>�F�D\Q�
���I�\X��p@!�=�@+������c�A|P"��l�C~WD6"!�^?����͔R��t�Y3u�7�RfJ��A;��H��S*�����!b��c
�) 7�9�xb49��r��Nb-g8��9�w��o}!J��n�]�c��/Ѱɰ:�����P�c2�0�h��o����f_���9��/��l�E+�����N.�XԈ���jB��R1�n��adK ���z���SJD��dDŘ��Ly���t��n�{W�UW���9Sd	׹�3>8I����`*.�D�[�jEP�o�n����W&տx�${7;K��v\�#Nŗ�,�WA0���f���3�@�Y���:C��vI4�/��ټeޘ�F�+D&Xs��}7D����*�I
&?�Q��|j*+e�����.�
��/3]Ao��ַ2d놸�A��bm����fT�hx��Q|����x�	���#k�������Ȇ��3�yl�{���x*�D,%f�_dU�@�c��7�����O��gu��� �A�̻n«���-@%�P��f��bf��#�q�]���B���.��ؙ��7r�4d����x���4�\��.<�����O��2Cu�Qgg�p��?��[m�X{#%�9ˎ`�Sz�Ŋ!z�rd)eApD��&��U$�L�:��,�Z��z/jse!>���1ϧ��D�K�5�DRw�_G_�17ɘ�h��L�s�V��2;7��;��	�I��'_v�ۯ���R�rs����A ���>��cq����0���z5J~���-���EgYi�3�`��Q��������B���$�0�έd��x��A�2`|8�!1�ڗ�� ؾ�[�����Y���= �!O|���|[w���ΓO�?��,#xs�=@d��9���g�d������j7X�^�l��lf������k/����	.�<<��)c,�5��bUT2sC^�^?Kה��;��ǒ����C�F*M)Z3�{lzv���r*�?���U45� ]�kr�l�v0�З%(蝘�,xt`��
\��W�h�h�#':zn=�'qpM����ņ����T��x�L�P[
iF90��H�,�e��h\�X��C�AfZ������+�`5�%�3*�s���Ϲ����*��q/����t��b�rC[��Tf>5��KiD^|н����Wi������D7�h�JϨB���q}�J��'�E���T�u�i��ё���T�hH�JL�]緳wY��;�\u6e����A2��Y4.�����4"�����b�xV�4z:��kE)�����ς3#`���� !E�Z�������6=X����>c��&��x�:��B���r;,�+�>�tWz�=�W�^�/G��Rͱ�$v\���NΌ����XkJ��%�+��D&>�'r��Mc�0
P�9q���+����2���X^�5�i�T%}/�<��=)���-�ۣq-D�
T'{�����Y`E��o�?oX:J�Q�L�s޹�)���> +*ׂy��ւ�����ٷ�R�Q�t)��!����ͼ��m��٨G
V��A��|tt�Fn�����{�1}va��|����	��k�,o�{��٠�r��(/���{��B����.&�k���Y4y5pD�2�)��O���n-*UԪd��	˷�r�k�iW9�-'�h�/��e��
я#��e��ASޢ��Q����kYm6��Jҏ�۱���C<a��ɦ׬���GN���'g���ԖP���8�GN�P)Z\0g��ג#�A����O�_ُ� �x��|�䅩���u���q>���M�nԌ����rĹ0���r���!��"�N����!^�#�q�W���2��0���T���fI�*��F��n+����4B*Kx����\��f�-�|�]��џ��J��#��SU�u�~��d=���bIC��'�z��i�'k����|_|�*��
hZR�M���/F�7m�N�z�Sq��Td�`�VJ��
3��\�M��	FD�%�N\���Q�>Jhfb����=�8$�����u����j�7�6����5L=���)h�`�����t0�=�5��,����kT�R�����H�oP)��q��sX��VL��K�eCѩ:fe��EG[1�>��tM�Y�ؼ�]�9�k7*��I��HY_�|3�z�v~+��o�`ON�
��\���;�h���ZAUS9W6��,��w��V�<��L�.Ǯ�h�@�`�)"^��t�����b8����Frnd��,�\5kk^��G˹�+
�DLڃ��>������XqB��A�U%�� �Fآ���Tfu54V6��z�7�lsc��ˎk�u�����"O`����h�ca�%�!P�m�*��K<�ЯK��Lv���H>�э_}���`�}`�VEq�{��n7��ޥ��z�?�������`��z!�t���wm�Yo�
�D���Mx�����.���)<��[�6a2����!�M��뉪M�܄6Qޟ�������PF��LE��DD�$���2���,(n�{�c7uy�;(���qޖ2��"Ncp+}�GM�A��ať�s�5����#��H�_ri��sS��客���s�*��'��r���Y�����y!���_G����D�_�B�X�5Y�����59��T�0&x�s�A�cQج�	�F�"[`������D��
�xk1ļ�z�0p����v�����oփ�LW��aB5���=^���cd}7����s�.Y���Sh����J�K�����o&�1�b�h�믚\&r-�f��8��[�sBH Q6v�e�31a?�7� %�����7���&F�ܥS��O�C�~s���SVvX[iv���H�G����$���c�P�ZH�7ˬ��{�_#�P׳��z�?/�3���N
%z�B���\�����2{`��-�c�J��e����"�u?��1=��h�ʛ�2��p:��%���N�논��qca���(�Ɓ�g@e��WܯӞ�|�N���w(w>Y !��M�ŤD���"p�QSx%�?ayYp�~��ۢ��LtL�@�綅t ^ƭQ<��b�d�6�H]7��
aVw����k$����<f���J?^/�Wvq�DI"��\97b�<�|Xl�
3|�fG�TwԞ�_&\�iE�WWT�y��4*���:��N<����؜c�%ͪv���ٵ��y���C)�.��ɕ ��wR�����p���d��Do�@�����%�A	�$K��">ۓ9�j��0���-�7���ee�Z��F�W�QD�r��xY�/Q��%j&��5W�����fQ���W���2�sW ˨/���ԫ~����6�����<�u�=�C����һe�ޙ���IJ��y�Q��q��?lS@@T� ��Tk!jcm�w�tjO��C�l�ʰ��m�u?)������{�R��&?�*�z��CH�M�Z�B�$_���=^���Q��Ī\�3=f�[o�9�@}d!>�WC��@�A��S~�Y]��K����m�#�4N�e�Ħ�4�]W�)���w$�>5��}����g]�}p�=1a�}Y>�9)��Z)�rFw8����&)`tp4���ּ� �5��v�D��l+�;MZ,ߣ�с��$C��S����^�%��
��:��"��:�w��[�i!�e5��>���.H�3+$�G��??�ݍ3 {_p-Co2� )0T�I%���Y�]9"1�vP��,�w�:O$�3���<�Bfҫ���W�h��{�.z���(c�LU���k��8��7��3B	�Os'ί�����G�5��O+�����t�v�X��K~���5��a�j ��Z�zօ]t�-�J{�Fa�L�~�����&Z"�	��i;�*r�nӿ�e�����Wh�V�}(��!y�h%��k#ս|@� 0�2��Q��Q���܈|nʋ�l� �,6�m����.{R��QJ`�<��8�#�������*��
���].I$�>m6�֯�Y���>�	��R��BoJ�c�Ē���&�iz���F8��;O����@k�"#p��#Gs�)l��[�$)N)a�"���d�)�@��H0P�����;έ�v��k���Y�$_뢶Ӿ`��qyE��&
��ـ��^_�Ů��l
��z��L5�(�lE�?״nM��HX�D����Y::ha��b���#/i�:�J{�3Hf�ӈ<����������lhm�0�~�C�)�=-�[¿��E��_�a�LݼĒm$���ט��2�{i{ܻ�K�* s��t�>���߾c×�.uy׹�D��Ӏy�?s�F�����S�"�Y�.7K�0^�v9���Ő�⵽��e�9)�cA{/�3�{H��"�	�-%�Jx���$����^>�����_�X�<�X&9^~�)b_I?Y�Laq�GC�Pl�y�gP���Ԧz[�r�H7�S��Fƌ:]徠�9�@%�׷�?�l��9��OT>�a?2 �:l:������g��gţ�ET˒;|�������Z)k�,�Hs�P�ˠ�[qLC���&	ʛ���<�����-7
���)���z5jo�\��U@����W�񨢌US���͗�ޗ盿�xnJgn`�ڸ�}4�D`�������r���"�LV	�m[4?g�Z�F�w�=���ݫ?�α�`�fG��V��y�X�/��x������Thz51������4���|�u��X|��֟g�q����J�<�]]L�'|�:�Z�r�	̅�Me��l%�+J�w��o����l�`����S�]�N�J�T���Q�� ��&]Н�:���<v	����4T��&	�"��&�r�wF����y��yR���V��!7����p�⬺��1�Z̽+5��U<�K�[�=���n�h�`|EGN58�O��#>J��@B��,>�i�����D���<��B�#�xE|i�E����UxNU5�N8�)��u�L��r��lITj�hPQ
Rw�9�p�����i��B�#1�̉i�J�Jq���z��	 ��ޕ7�����J1����F���MG����/D�ՙ2���=��M߾�az
֏�1�p�g�=�D��L��י��~1/��x9���#�3���@�ǈu�m�V��$�,�p�F�5���1/�����%v���p,D1B����3G��K?�ǉ�o��t�EK�{"Y9uyQ!��gq��twG:Q�	d��BƑヺ�5��	
�E�h��'��O��@�Is
4���ٺ��N����{�P�@��h�S�*��s�ж�!��%��$��t�<ųM�������T�͝���{�N����M�?���&�C�6Ķ嗛�EV��IJ�-[�n���]Ҷv�R�Z�V'��&��ҷf�і�+�:��|��_ٓl���VYOi�)C�ċ1��T�i]?♪��`�L%��C�U��(Å�����_ؕ�I�m����3���`N�
O��yx 4�~5ɣe�-�j& m���'͏��,N#�eՋ��ga;8X��:�*�x-��%+���!��?��.��Id�"���˧��=a(�ڷ���7Bd7W�M��8Y."�+��E������f�6�C#�\!�o5;�E����� �]��5�v$o@.	a�Ơ�oD]Y�ȏ�'T�i <5����b L}�#�����Jӣf���qK%7d�����R$�V����򴆃D1}�A��~c�$3��B#u'�=�LO�t��h�hT<ZVz?�N�\h)��j��A��@f�!;}�x���������������ٛ�l���g��O&�����\`,@��ۑ��^0R�/u������xT�}��-���Eb�Ȗ�xY��ce�+�<�By�C��s�+D8N@XH*�&�E�M�}/�l�+�
���@E�5T\���.;�?/�P�C����;�u��5j��\��o�%Α�R�"�ʃ����A?F�W��j���{G�����m�,Gɑ�=7��~�`Xࡡ0+O��v��+��^��'�[��8�,uF�Sz�A�,�\Y��5=%�5�8�d�?/���xx��l��B�H!�b��4<>d����Y��Z+l[� l�-�ɐ7���������C�Cح��-��IH��QΗs

G���J&�ZH����$�v����GSD3x#.7P��9��3�
�Y
;ǹ�����!��z��
X*]��I���GƮ����؍�U)^������+��_d&W!�0~��J�قWsM�g	��/��+�d�w!������*�Q�Y��,*�C���t&��=	Y�A;��6im��`1<c{|���+JJ�T �a48Y�+#�����E+�=9�#3H��cuG�G[�Z3��=�ؠ"�/P�7'�h��Ѳ�^��
�yZê�YU�_{WI�s���~%6s �D�6%�Bn����(h�q�P���
<D��w��Xs����c�/̚�>��)���f�\�
`eߒk�x��?�����Ȍr����H�Z���!�~5{�����ꁈ^%zS�������6 ������WG�JuV�C\馈-��S�������,H!�}�$�\5�}ӑ��r���-���p!}��bf�D��^�yɅ��'��ډ��껶YV����Ptl/�o7O���-�o�A �TmU�x06��8j�ە�?NAT @f�2E+1	����&rr�TVx� �D����Ǝ2����U�5�6!cҒp��j�Y^�"�ߍb�{�,�/݁0�r� M��>]F&$��bgg��y�M�,�վ�8؅����������6��Ng����!� �ю�z�s��!�Xn�:�p~U
��C4$�~Ӗ)1.\�K���l�ǧ/�y�\7x7�n�B��X&���q���s0I&�`�}I�PG�;���m[ȑ�m�������w����Q�y�뷄O��ӎ7y��;6ؠrY>�iJ��x欢;���EU��E=)�L㬤�t����c�	���ˆ'4��9����4A㻫������>�/9�#z))�9�Cv����K���>w��S~*_6��B�p��v!g�f�4���ړ��2��T����p��oٰ-2�U�@ �d���O'&w;F)S������74���f�)���-г��;�>�W�	���@zZ|��w�Z�h�P`��Y���.��ER�e&$����]E�m}x
�E����p�ݩ]GІ�9c���%��у�������!�l1����
�^L�5e c�ز�)"�և2�W�:��L�������� ��wv��֥�����~!���Wz��O'��T%l�C%r�1��]A����~^�w2S�cҼ���Ո��_T+[F��as5����@�S��:�6vȔ�!���@��DΌκ�U c���%tYy��X-��i�"h���:]����`���l��y�^璉��7�����L'"��k���2�Ɯ��Su�o;�|�R0M�lP�(q�����K�M��0��`��?��{�?ߴ��(w�I�BO��F<9=d�h'�9�0�����qp�B�Y��<
C�P�'G0I@T��d�Y:<>|7�DC�N�BG�؇�łn;�Ō��;�S��F��_�=�����1q�i��Q�Ox��/���>��K���9ӊ2��%:r,��
�0
��h)�7�^Wj3mߠZV�ѮO�Q#NE֣C�>K�F�}/�|�hڇ�?�=0�+���;ك���7�tx\<���|^K-	|V�F����d&��
�!$��$b�)*�,Y$�Ā�7�y��L-�b�@}�`�B�6��h:S{�c
!�A�Dm�yJY`2.K���	a������盦�k�9�o9Ӹ�"sr!�8-���"gz�v���Lc�/��Q����k��yZ�7�g���a�v��Q!��F�8Z�p־u��>"���Nܑ��� E֗y�Z�*��U�ENZyG=������`�͇\(��AZ@�'�`Ү��I!
A�i+���2��k�����V����p���c������	����HǑr��p���l�Z�G�/�m��F��g��+4�-���v�$��y�:���K�kڝ����Ҕ��e�m~*0.�CuӲݾ�1%rc�q��3�r%G�`´+H���H�ӑh?:���lh]�PC�T��e!+ �D���}�P�_�Q�׻B���"�|g׉�0�	�N\H*4/v+\���t�Kۘp��ҧ��m���<ZNɢX?+�D�5bRl�(k��U��+ Un��* �NnZ�Pip�2��+kLM�H-�:�\~ߞ��l��#��"�����(���%9�^���EV��
G���b m[˙O��`�ZF�U�pj#U��˔����2��I�o�\��d���ߞPꞌ"�^���sV�*�;%Ԫ��&b�� n���N���
��y���"r��` �xN�%h�L [��opF���(J�T:�}������{�]$���R\�C-`��v. K5Υ��{�!{����B+�2@v0��^�W]�/�M�4M����G|��K��t��;�= ,CQ���鴋ZC����u&<������_�t�G�CU��� L tQ���Wv�Oq����h�Sl�m�t�+�X�Ad���o��U��!����y脲�d���(!��1aM� ��h\�����h<e�C�|�Ě�7^X����1��3�I*(�AG�����/҅��Sh���e$��jZ��K��p� ������YW��z��0�����f���a��n5E�\����jN ��O�����t�,{L��)��<�;50~��D!f�\��$��Vՠ��~c�T���+;�#�EW&��b��4 7}���;~�G�W�b�T}��y	���ӝ��\��,�{������pTm'�����	�����E�B��`:�l�Eσ_��cP�7M��t�� B�q;�
;�]VVh�6ӎ:�P\��êM�le&���y�^���w�km�?}�D[P��j�!�T�����-m�*�>����Q�������@%�U�/\gP�3�"
Omc_n^y-�}�(e�W�wl�&*�P��L�ٹL��>�e��ǥS�Ȑ`����p�莻@����v+�I�"ݼȋ)�ٜ-�l2�N��^�ڥ��J��1�C����CP��G����Y9���t�E��);�6���#��Ca��w\ 'd!�C`��G�v��؛R��rSzxu(���]�8+�CIU���+�mN9��0�A��T�ֆh|d=ct[�SBZ��r�>~e�kJ����|�C4+M���"P뱜JJ8�WA�C��c���\�ٗ�.��Y�h3����o8�x�9;`�Qq�-g�w�(N��{�|�>�͛?�u���w\K%��{����Uݨ��:�'��	EZ�S�h?��ݻ����+T��c3]�RIK����9+%{��y�Aţ��c��������kc�D�W�]Dٵ'�s�8������c�V��k�����O�tp�
�>Z����N@�V|������C��b8u{	�a�[L�\�ϱ+j�?4&�.��"/{��w�9k�ڀ7"q�eC�����{_gig/�M��P��?y2 <7=;��L��=ov�$�v������w��tٽ���}�Pww���K;�c��T#�-O��0uV`R"kǋ�Q{	�Q�I`Io}~<�Vr����[�i�(����7��V'G����(��"+�ƪ�k�Q���c�*n3��\єx լ*v�Y��Pg�n�>��-߳,�L�{Ɩ�r��M�k�8�L�%DYcf�gWp��Sh>�����T�ܜ���Qc�O�µ���e+e��1h�;��W�c;^��T1���t�6ɠ�QH�*��e���b<�g����d;�e~^�6�=%���;1�Kr|�w\�H�����,)�S��{--��g�fr���\
��m�?!#�+�ݧ�u�N���p�T-WY�+o�&E#С�0���/� K3�xJ���,�Ew q��<I?t_�` �%�`kdk_',�c���[��-�/A�Ci��g����w��y����� uB�Z:Sy��H<��&�4�qd���O�֐�k���ws3(t���(�5:����8o�E�
c�q�5�]~2)c��:�.� oI).MP�d*Ƶ:}_��z��.����o��^J�i<X���HǮf�x��3����O��A9;�ʆB���������P��ɕGPJ��F�iM}Z?�EQ?��P�l(pC�ϓ�&
��5}+{�ɥ�-*��fO}L�s�ni!Rm�Ɖn��J����~�j#��^�{���Be��U��