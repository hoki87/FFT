��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ����������]w���>�}�*�8E���Ǐ�36D_����D:�&Йu�%�BZ��cOR߃���>�k��&�A/U�oՁ�H�گqvD��|���H(r^%����}ȭ޲I	�����-�����t��l�Ǡ��l��(�J��������%Q��`�7^����*�2^6jW�I ��I6�#��#�^]vEN��D�m���S���fo��n�w�E�p98vg�7�1���IA��EϬc����&���z�/�Q{a�h1�/�� �{
ۥ��j�7�f�s�����_�.�9ྜྷɊ|�N�jz��^:�����9�oE2�`�� BD���;�]�N�#�@O�&4�_����h�L�Y-(�5�*l.�ֿ�`I���e�����ā漏��o�n�+R=8~ ����.��|�G;��D�o
?�^h��n�B.��t�� �>BX���?�W���5ARO@�J���R�pO��"h>����/���Y�� 9�0�{#+,k)�^欧���݋�{��{{�Te*)��"����j-��,�2��-�6y?�����~�
�!>�M�_��앳��+�J����.Ei���,�9���?^!V����t��~���)���
�X��g��7����|�䕕T�>;EA��3��Y�'�t�۞-H�Z׏���'C�N߉�����'AA��S�f��t��H�\D�������9�o��Jm[��^��t��3E�
�P;�:�hk��+
��E�M��(q#�\��E`T5� �U��H��M�m4;�ܴ.l�na�swe3�	�����UJ�o�Vx���Nq�����ݧ"D���;��*���9��LoO�i�C�!w,Y�bjȢ^|����h�E�{��.�M�p�(�AT�Q�Xl�[xU9DV��u�\��q�s�9ܦY ��[
�{B�k�5j�ׇC�5��'C��=Y��gG65�@L0u�����Щ>ֹ�P�Lʴ����_��"/e����@w�u��`�����in]d0/���^��$,�-W1�)<��VH�+�18Z�*������W�滖��t\���P�G�,:��+�9�V����\�*[w����uP��B��(󎞖�%�Ϣ"�^�{0~��;0_�tqY˓�?����a�t"&�w߇��}�E4:#Cْ�l��Y�X�t��������a1���)�,��@�\�j33'ٚzb��W�� �W.��y{��y4�䠍���$����Jj/���:� p�����i���x�$U�H$�����f�)�7"0L��mR,dT3��$s��LA+Z��r�\�}�+Sx�dp���wii�GK�x�e��qM��\�C�Ր[üԊP�k���/�����r�H!+``�}�Τ���e����0l,}/��kd��R�J�O��'��d�2�:N�~�7e
�������5c�iA��[�e��Z=���/#n�	@0����OK&�e�Y�J	�/��b2��/���Z> ~GL	 ����Êdy�l%	Hf���5����._��.y�����X�@?�a0��5�;ӎpA�k�4�iB͞����zkʰ�4ʁ\�������?�?X�����[��-���a�Ѻ�#6D�1�J�_��D�mv�L���q������l&
�|^Bru�gD�	��e��D�1y�`��s�-ʱ�N
���3K3����xX'�'{�Z��2
��
z���?xY��o'e����l<���V��$ \#π��PL'c$Ql��r����U:[;�C����"���{��s^i���xP9U�}�~;���,����C~�r�(��cE����9躿�*�`2c4�k"���!ɧ�����H�F����Fv�P�6+��"}���l�򞵶�T�@�W�+f'(lޯ-I�?�A%Jw���*���A3��P�PԘ�e�W�\��Ղ�F���N�8�\,p�m*y?���/�sIR����L���u�B���u�����!����~Zq�oT�u�ȉ��d*�5�����tМ��U�(F,��OS�?Q)����ḧg��#ڶ=(�I<��aw#J7����������3�����*i����/��l��ǻ�}bֲ���l�'0o�#8�@��n���쬞�\^��fIU��֙�xJ��n��scH"���)�r9����_X�Ԟ�"�

C�_�lv���_�R�Y��L���#��A��I�w(�� G��y��%�hRq��6����Xu(s�(������(���>H6�"�Z�.5cD^tY�/5�jE�NK��/w�q��%�
8h">�ǣn�*>?�p�K�0�y�̾�@�Z�`��+6�F�\�����f/�	�MB LEt�߇�����u���U23�W_謥LW͵1[6 ��326�����jn��%�����?ۧ�	s���܀�\%�s%ȱ q�B��8���h۔���hJF��q�oRǏ��-�z ��n�'��ˊ��!,t�y��o2!
�ʢ[W��v���M>N���ٷ��9�E|2)�Z2�ɏ!w�С_
��q7�qI�#�@��=��K+'�#Bk���2������o��h�.6��^-}�`�7X�754D�?��mIj7����WZ�l��ĭ���9�m_t��0J��B>�)�2)i�7fDQ�Eo�i� ������R�;0R�ה1�f�f���c��DF����ھ♑:i�]po}��+�}tk��s�{�(\�NU�Ñ:�~����t�j�%���)dnwx_&�'?jw�	R�B��D�l�K�]_	tW|�j����Oj2ʂ�oM�r���Q��:(a���7y��!���4�͞�N�X��u-62ŀʓq�K�3�������BS�x�Y�J�N�D�u�T����;ƨg��jA��FsA~������9��K"�oo��"G�>�x �;�~�A���P�ϓ��p�?uya�ب��w0˼��䰩Et�桻�A�e���-6d��r�&���O�f
޾}&z�v�Yn��hY%��擓��b����n�΅�w����nJ����w�o��y��쌸1c�]��4�?�r�Ú*=��B�D����jO���Ȭ��㙓w�x�f�ٙ�����Y�����P��m�O�/�M�r4��b�!A%�؇�����h]����/�J��i�yg���RӮ�2eh���XIx A68x�r|�R)-�͙>l��w���g�haЈ�Q��i$V�i�b�J�,|�rU �2�
7��������>��Ma�;�������ki�ϛ1��Z��!�&�UW����f�v �gƇ���3n-lM�����ȪY�6��>�n��ϝ��T&0ATo	K��\����`�R��3��Ķ��v����j�,�|+�`.�"�Є�/\?�j�k1�f�Á�՜�	n�ڌ�c�	�Q�$�o���U�
�<�u��
]�h�����?@�C����V�o0E���wz{�,3�����%%��������Ds�����cz<U�x;�����P�[��=;L�P�ӆ������#0	�{��=�{z��q_Y�X�W�ցԜ�%�ngY)�]B���{6�$��(�v�f�=Q~�	G��<:Vz�|�Y��LJ��l���F�>��q��w#O�Ī-�*�c>�f�UE㿂��C�qR��~`��{yn�خ�S5z�|�	F����sQA���4����^�p���Z_�.��XO ҝR��϶�̱�5<p���H��q�?�B�59?�	~�2�U����s@f���a� �0�pa#A#ty�a���C=��@�s��!�9� MEB�g� ]��#�6��!3W�E�?�T�>pc%�e�E�T���^�,�����r��<x�R����!@0�V�X�����Mf��ġ�>��H͜��_��_&
x"�*�ɣfo)l_��j#�>�_�]z�q�9�u�&*i�ٳ3�;6�Z���x�,���x�{b?�ª�F�����	O�g�����惕�r);�:Fِv��#�7j��E]u�u�t6���s�d!�L=K�G�)��*~8,���Q���?%�^������Ax6��IjG��F2��W%�K[�!0�L���Y�ڒ���E���^���b=���7�5�:TN��I�5.ڤb��B���|ulЖ�S�()��@�?�灒y��802�fٍ�ۃ��:fI��
 ���HkR��u�](��ح���>�Y���^b�Ɩ��9��E��\�o	j����a�7"�I��4��>.}^U� �e�֚"�҃쇴h��[v`������m��/.�A�i7i$b�
ď�ǈ�d��ث�qn��1t�C�J�����:�^��©
�&�3��Ti��n}�#�����ո�s�楌
��hn�݌,����S�3I�T�-i[��b%���U|�9�����"mޮF�����7>��[3u�H߇�Q3YO�Q���.��f�����������<d�ֵ��Ck��X`2�sn9�hU_�b��Fy����me��jz�R�_��;�6�� ��uQ�.a��F.VD�5�T�_����G)�v����]����\�g��+A����T�7q�JUz���t@ɤ����V� %�	�ha���U(!����/@B~�E��Sg�ڝ�y�>�a�cn����7ӟ��Y��C,��'��US(B{��|~z��n��³D8p��0I��i����4�I���p����=��W�4����i��$����lU46�����z�Tr5-l�ґ�^��Z�9:��	@���\2f~*�rZ/�v��
�;;Q`.+�-ޓ$��t�}3���VoYz��g�i��k�ThMu  �K��p�64��<(���v�&xn���*��^�m�_7E�%Ra����8qHБ/Vڕ����%��O�Dn�G[�N�q�3Jy� �_�K�ִh)tnE`!��{c�Jo(�:��;��P��"�j���-�SK���c$EV�@�!��
���^�+{=�1{��?J�g�B7���U����D��E���E���qj�x��:��H��%���Ԝ�9�{�0B��e(