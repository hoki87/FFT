��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�#&��#�<������M�&ӗ. ( ��:���n�$��j/N4����Y���;�{��p���&z��>-���Ν�A���E��&�;P��1qqzf����H<�����C� Vޕ���߆)��ڊ�U���|� ��_:5	���cx���,c%V켥l�r�Z�ؒ6�;E)˥���-X�����*�9']Y#���j��&�dclY�x`Z�rW��װԑn���]���q�&gNݩ�i�%3��=ճ��?-�U6����B2~�IY՟�8 ��FEH~��m9 !l"����\��e�X�۾IKI���f䚓h��-��>A^,���G�<~W����I.bP�pJ�pkfK��9.*�M�Qu�����wޭ�92�]�F~KS��T�y��4jq�Q��4R4�k��kt�g��I���kY<Z�*�
(����S�wM	�Yz�F��Ž����0o�1�/��N���2���8;"�`&l��� �		D��0({��l1���zLA��~�2	���2�m�QZ9��@���_]c����� ����b�|1>�䩓S��A��3�l��q�2�`���ļ���'�����+�D���@t2���J�f�p|�p�"���wv�y��%����YJ����5�����r�F'�T\��������v����r�Se�Q(�o��+��5�:�vG�� ���PW[H"���G��,�����D�20έ���J�D��_v�<��|X�y��ܵ�yA��m@���B����W��iȻ);1yd�+m����4?w����Q�\$��\�TQ5}RkI��.�!���xn��!�P�~�[�U[���GR��W���=�q�"74�[*z���xeF��"B�$��=�����tԣ���ÕF$M����1F	��'�R;M�k7)�Z�P�I��X�*"B$�.7�� Xk��",z=z���?��0�oj%@�ފ�Vm���^��(Z%�7ن۲'?�:�U��d��[�����ɤ2��Q7&�arY'����)	kڇ)��ک ��:ۉB,�j�pf=Fi@%�
n;Rdi����v�H����a�/�v��?���_=�*k�?��z� ��J9kG���Y����!Q~�)O�_w+��վ�]�0�"�bgzlC>�f/���lF��F�0������� ��B,��1J-"��E�v���N�.ܑq�G��7^���,{���w�r{~�T��n�ढ़�?F��S��Y��>u�M�c���ܒ�9�'��/��B�wJ�һ[���ԝ�@)�y��4h���3N��jX8�^�m��/�JOs@��Z��#�6t��A7��,D�M<,�'�cZ��F��ja�,}���fO-����'Y�	���x&Pz5$��u��y~ق�V�%u��@�0�M����k$��cP�m�2H�h����=�u1aB��9�ðw�{K�����_�G�g{S9�fo���4:@R��R����ު�2\����ut���k�14��"�m� ��S���1�%E�i(�ֽ�&��yzr�-�Lj!��SS���k��'�|���o&�l�j�������L����Up})�|�W,�y���Bz�s�r�����N�LWz�́b�s��)��L<��S�R���d����a�soO�>4}Q��l�Oe%h{3e������: k����)�!U�z�Q� �e��O�������=�]2[k�yGt���{X�sl�#j�U3�W8T�Vm��X��f�����벫�{~u����
��⃂���{�$)u��9*�:�<���Ty�+o6�て;)�5�(�Bj�	��ZӠ�\�����u�Z1��R�	6c7�[�����/�KYDU�j&��e^Å�*�G-_	�s��	:Vw|0���:>3���ۻ�+-ucq�J�M�b��� MM�%u���4���Z_8���c�5m��c&0ya~�Ӕ����6�X���ՙb��/�en �7�@���:wc+����J1 �ub5	6��Q�1C�Dmj��C�@�@���a-Y�
���*�H$�\�gi�]ױ$��N�:�M�,������������AZ���	���!/�����޷l���{K��T	mJvcj�"��F�����lD.�i�}d��i��eUL�ߍ3C��̇�v�s)�;��@���Wįר:p *�m�F*,Ii�����rm���neX��>Ԭ�飇��� X�L�<�0 ���S�B��X&��ث���f>��)�.
5���k�_ulծ�f���{t�1)̠]b,G0DUD(Us���x�!M�����`�2X��$���Xjc�d�bD���i>WB��*%M5�O?W`V|%-=�'A�i�x���lY��gV���_�<j��_��6~���b��i�Z>��&�m�M���Y�Wj���2�p]Q¡�z���\|]��k�,+���v�1���	r�x1(�:�cg�^a��42� �`8��W�h��s��_D��'_S�'h�+�8K6�:1�G\�:��9��o�%F\z��N{���񷗧�(bM�w�64�#����xi�H�ho�g�Xo9�:_IF|��Ǎ�HUXSX�f�=\�G�G��!i8�cf��0U�9%t����dW��Ex8ꀾ{��;0�<P��{	�&"�-���V0i#_2�D*`۳�D����=�5�2a�E�������s,���y��#@�X�>�u�}�.M�3*�Ƕx$�s!�E���v��)�����7��K^6�n�w�8	����tp+@�Dj�p� c��ν&���I<b�K�
%(�BRGB���c��BV��)�]L�U���仕���a]׀萃��s��;M���?YH�� ���.<�@��������)1��-@�)��|��0��&�����G���N��0F/�&ǀ܈X�:!oP��5\VJ�S�
o�f��Za���NՈ��A�9/C��=Zq�\�z��o���\��N��g�ʙ��e��|��6*�1�o&��X�j�˱�5�vE��D_�1mP��o��w�4�9�Fr�p�;��+&��xO��h˿��bW��c�;+�j��|A�K��ּ��p�X��|���v�L�╗�D���7������`4� ��@��T�I�/R�:���bj��͝�
\���=�
�;;�`�=zqm6�񛻥��q�t3�C2�][&�\
�@�g�C��f0�jA�SU���k�v�/�8껎�4{���� ���� IB���YIT�TB�ߴ1�|����ۄ1���q�A'.�Z�C>4U�SW�#�&�V&?Rox1�p�	�0}K�b8�n:�S8o+�1PUKw��9��|�PC3e����_��<(F�J[��h\��0�2b6�"U��	Z+��T��8��J�C���(�ڐFusox���1Y&�I�+j�L7�~����I�0���z~|!	�}C�=���e
RJ�"�:w�\�/gbPj=y5D�ō�R<E/������">� u"�d��`�m�:�̩1�w�Z��T��dʧvc�y;����/��"�x�r)K4)��f���������J��tl2��V�/\Z���<��A'��V/�ˣ{�^lFd�u\#�c�_<mW�h��@氥�#��&P�Z!�xGTzʅ�:^�u�H�Z��4��ZT�M�q/G��V?^m\�p�SmB��:�g�.�4���T����b��h@�S���"���?㥤Bw00��5>�ZD�-�iǵ��N M�\ä_"��j/�������h��,7�:���f�'�� 6m�Ւ-O,��E�v�:y8\�������]��D����҅����,�2���r�ckܨ�&�`fD5[nF��F�'֡Ƌ%x��C�B("��Ĝ�w,��s�,1sif��ک8��҈,��!�Np"s����ܵ���8ڌ0rV~:�n��N��<f�J,	KJW� 	J�]��Dy���*�@�t��_^��S��[�77��? ��M�[G�@�r\�kS��:���Tm����A9�(Rx����S
��9>������y6�Z��
��F�tę���e��!ޛGJ&��4���	p&%���f���"ZnI�3#Cb��ہZ�)��a�,�gV�e�f�%���zxUq0Tp�����J٫c?���/O��|�3,��t�B|Ԗp�=�f��֫1��p���Rr<d0U<Ӭ��֯��~{�8c����X���|IKg�ڷG��5I�-&�!�@�9�k����b�$��33���\e,Ө|(>i��G�b���N2O���BGf����e.�.}����9��)|7jz~x!E�9�Rӆ������ZzA{ِ�?^0����Z�(��asRܗޡu�꿉����d��hD�*$����5o�q� TRG_�ni��3��7&$�_e��Uu1��0��h�j���p�Bh\�	��f���]."Lӵqˉ4��r ��>�W��V2#Bs��aj�-����y{�M����f�e�J˜��3!��.Bo5iGO�ҵtƬ���k��ê��5Ć���?��)ʑ��>���j�03��݄k�m:F,��j��A/��1r�}t��LH�>�#�����&Tؐ's0�~6䰾��Ζ)4�2R�I|��v�����hKe+8ri&	�i��HC�Y�g]h�����hjNkE�^�4�?W2�D�K�~��Z� �G#�+Rt�����n+&|�xā���k�$I/�;7�O&B�����vv�H�#�Xؖ�xR"�&<�Z:������$�]��̃y������P����j�h�����P&Yrx6��]�� �48��Os��q�<C#$����4�b!��D��Z9�	jQ�@$����s[9#*�/��]w'��?�/ؕ������H�Y��UO��V���Okjҕ��6�}��/֟ @@�"��wG#�j�;B�RP��f�3?u�|#g�?Hl/)?4�����9��2�醲<��]Do§t����h��Jҳܣ�$D>2x��Uyt�ƫ@����R����^�gn~�� PI�x�\���Fn5�zp����}7D=�MF/����U��u���_�[�ʾV�;�iڲHQC�)����L��ڃ ���;���3ƶ��=�!M��a�D�Sb"F>��6-���R��&� �A��J�x��>1O�Hb��Z�S�
�oH&H�o����1�^ī��]D���h� �