��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#���������l��U�~�׏O����j9�PY���`T���x���s����uí������P��"��b%>�1eτy�<�gܰ�N�Y�	� {��I�ɍL�ݫ�G�R�k��Q�!E	�5E��.��:�͂2��y�m�-�.E��i�����YS�
��@�H�ۼ��nD��Y�l"BU�.TԊ�=�-�����q���Ǹ��j��ԋ����tr�a�ٵ�]�b	��%�ɔe�)rYOjX5;V��R�������M\�	D��ҏ����9c=�Vͼu��Ro�P�Jf�tRvsY��c�"n�XO��	3g���Q���^�Bʹ�7gQ+Г���$�-��t�8�����A���<����l-��*�|d���5#�z�{{�����aA���]7e7?(U��Am��\��?-�J���*14�6?��tt��0�"j���1���*���i�i��ϧf���(�E[6Q ���ԛ���̘=��]3���c��J�|���nA6K�D$^�To��_�ꢧ#-?(9i"�N�������9��X94��^�T*v�b:�t2�q�f�\�s��j�1�?(�AA�y΋�6��j��Rt�Vr3�j��-�RBܙ�(�J�X�c�&�&�ͼ�Y�X�{��Q�og��	dw���]=��>��3s��BB*w�:^,���w\�}�mn��U�.e�d��(�b�@�rD_p�w�H�=�e��2w�Y�R�M:��d�I�-�����t���=�9_9����l�H/r��~����� ¯��X��s7S�hӳ ]��wI�	vo��o%l�D�+���Q���%��|�o���ζzi&�$�|�X< ��Xְ�����v��0�ӟ>����AHg�d��0i'�ٜ����Ԍ����zQC�d!�F�m|8�Tc�A� �H)La���6>�9X�U�>^�W2�d�7��D@��5��\@G~х!<3Y���]�V3�kPPj�&X��3���u�~Q��+��.K�z?�����'\�$���R0e����y)O�t��;S�p�{�^����i�P����H��R�ʁ�~m�X�<K;@�2!�$��1���%��,Q�+�B���0���|ٶ��<��wRW�.��5��[�,�;Z3����i沅կ��Q�1V=��X��@|����)�P`[� �6��A���hnxKq�%Ш>�k ӷ�Tz�l��Q[�V(l��'����7jH��(�B��C�3Ǧ�*!��D�f��`iwd[N������k~	����SLX�LY�G�Ά�ȵSf����w�b+-���9kg��x|zA����"Ȑ�hӂ��lI�����=��V~�S� ���I&�����$k�y��>]BD����/�M`�qז@��a�Y��)ǡ�Ԍ�a�c��?������4AX�.Ϊ�1
�[����C;=l���b�eZE�d9y�j�/�����K;^̿��L�t6�R "��x�|�q�z"H�x�cL:6q�+(��s>�W��Q�ڝc1��w�G.�4���Zt��匏�U�)-M x4�l�u溕If)9Ȁ"��
�M��el���P+�&a� �P�E�P�&Z�KOo�]��j��r�ሦP�cT�P�a~Y�H.�����_�6̅�����Ə_�"V������4h�P����Y-��=]K\��vVeuOl��U����6��ț+������U�.a׬�}lsJa�~n��K4�Y m>�eY(7�3j-M��8T-��/��Ip�gSYO;�W�����j?8�.G��e��g���o�Ñϭ�ፌ����n���3|��7P�@\�?��%���dW��K�L��z%G��u7�
i�_�8YUD)��"��1o���z��a��3�L�J�D�I'�l-mY�;�_)��`���7��5�8eh��$����>�/�ױ�լ��oF�H�˱��o�����]��.�Y ]'~=I�U���X�&e���>�i ��&�^*ʘ��M��gB���L+�:T����i���oA�gi���(�\$Z
�ϊ0i�r�A����53�oE%�*� �hshb��<����(���S7L�%��v/cة�I:ŀ��A�Z�"����U�ѓLvN��њ%ڈ�	>�	�"�~����S�Ml�)��� }�zT0��?���ں��K�����2oi�2~�m�x�R�g���Φ��vew���Wڗ�YN��'}�.�z-���T��=�r�W+�XEm ���=ޡ�R���ʞ�rh1�	�5o"�B��E�݄�}�|���';�+8����o�U���-}*�+"�;	GpOG/�If�F�9��9��dK�f���dk��^|�_��8.���׭���� ~��
Ix9�u����)*��4�8(�#�j��n��=����Z#$��������rl���.� ��>���Y����R4$��_�S�|[5y�qu��7KK�2n��^�Qg�i`<�1�i{|��3K7.�� 
�K�8}X�F���c��H�%��LK�5�s�����'ʄj����f"����6�3�G�����5:=Ҏ��q��}�K$"MkM�&N�����ͱ�65���1~E?�\gǉ����l'��5>��ɀ���Kmu��8Y���U�q4'i�&��Y��i���	F�?��;3�]R���#�2�T�o��G��dP������U`��	9�����8k�$'S^1����G��SDw�~+���ς=���قݓ�ӜE����w��E�E�A�3���h�3d5��+�؎�!7	-�z���N��3��Ed���K>+�n�_/6���6�ЋGp4�{!T�Cy9t���������u�%��he�dRQ��_�{�ЋF�g�]�]{aMe'F���v�$;��Z����z}�>��\�A��/\c<!n�s�R>6�h�l�����X<�s<��/;[�ne2���~?D��(g�M����b��JI�2&4�ϫ�ó�"�D(LS
�-�_z \F��+�M'{V����$��Dʾx���w�������~�7��n_�h.��6��_���/���z��$nV�_n�l�+>�2 ���p���8��K߁|`VL*Z�f����Cziua�L�χĹ���n���������R�+�ԃ[�=�y������?Yg��I��h���!�o�Q�3Ө��LoSgڪ�K�Vc<V���"Z	L�7TfE�#?�m,j�n8Q�r���[�')D�}�Pͱ�>�Mn��u��ڷ}ۈ~G^���l�E�é�c_	���IB��)rsA�nq��lċ�O^�F�>���u�g7����.�,K7/���=+�=C�����in�>R�;i*�y�����C���:�,���Jȍ��
��T���#��E����1&��>�"~CnټH����$Cʲ��y�65l��V����=�s��2 ��o���W�lU d�,C�"�������K�,X��^aDD�����1�h|,[^�w�%��Fu5����v�TR�2��E�G�*�7��z����ǌ\�;~yQ�
�L~�ȔqB%�ד �#F��R����u[��xh���#p�RqO�˟��ǉ��W�5'���u:RA��g�҅��*��a�)��#�ƀ9n���Hlp���.y�����ZVi�jO�q� ��-?rb=$i-��kw�8oB�?HJX��i6�z�T������&��U��P�b;-�u���i�R�H���q�����z��}C�U���t~�����t�Q��hޜ�m�e�_��=R���=WD��({���'���v� -�~r�뙃�	ѵ���g�L�>�OuRq��j"9��\�4J_�Z�yqe
��'�v���t-ob��a�P�lx��UζYCS��,�Mu�J���r9U��;��ͫ�A���;�x爏'����qw/�־�*N��@��.�;�{���`<�i͛�����v�!��pF���`]�!��/QW���F�@�N1}Y�:(�&��:l��R�"�h�8{������f^zQȧǺ��`=h�4�S`�ΝU(�������Q�D'A��װA��0& ��K8����[F*w��C;J�YPz��@ےGc�ޫ�ZU����!�
�l˗�*��CӸ���P40�L�Y�$\�����[r-�-�W��/��d'��{֞Gϑ���n (b؎�?���:�=w8���z�kN�DlK�	������t$�MP�,�9���YԬ�gc��;ʏ��et�L9����M����q�'}�t������|&MPt@��?F�:d�c���U�3c�V�������6���;�jt)/�j4^R���`˨9[�G���"s��d Z� ��^@KӶ?�c/�S� `B�)X>$�~CaQ���Bj��0D����[I����DÒ�r��Y�ͧb��!���qJ]Tu��A�i��uJaX��d�
Б�r�`�z
�ۆ5����<ON�ⰲ��C�V2"��&��oH���uuli�:������V�I!��7����_6f����W�m�"���i��!��g6�w���.�W���{�DE����[[�@�=���Np��y(!5��G=BI0�X7����_���$�=�#	�o���ȅ&���E�tX���*�z`Ĭ`���^r�.D|P)�V2�	ܛ���u;��Bv@�(d΂N)��@����y[�bI�N7��/�u	a���7�h��m:� ����]�_�.�\�1k�D򅤰�/5 p\]� o#t.̗�40�N<����W@�� %��L�'{�`Dy8�s�Fk��뒀�F��#$�#�ӱd3��F��y#O.����z�!L�*�M�w���^�ݝ���v<�>Z�j�cA��§/��w�V|J��y�~I�ţ�nVg�5z,]�B�#�q����sH�����(��ߎI?v��KXCϼ�1����S�{Kܶb�K3��	�̖�B����^����k����֞z������9A����c�c��ӑ;
��xmd[Qne�*�q�ݓc;�;/z�P�j�����{��g�
��*w�
xQe��"�5�8Н�w��2 N�#�2r�M|&���
S+�,�xʴ;3��
��`$���J�;2ԕ�����4=$��M�M��AU:���S��;!�l�2��m�bF{o�	���G	�p�w�I=��S���s'k>���&�BS�!c�}�j#�wz��D-��2�u��lȳ�Jh����r�1'��lH||;�^=^O���jm�[�ÓIؠ��?���L������Ka�8����qahD})����+r?��izI21�|	L�ƌ�� q¾��o �g	��O��@@ou:7���?������7*C6�U�ض떑�f�bs2?yZ���
�O�h��h��H7BL�&l@�j�f��[Pٔb���j|U���Ue�B7���/�.��"��\q
�}z�|*p�}�� �� &������m��̬g��?4a���y���^�|�t���Ps��?AIN�$Ej��[<i���O �q,���O���}"L�2qý��T>dT�S��:�A���ɬ28	�����Bf@8�1��d�BȊ_�l�T�΄�s���Ow���_�ݽ������>r�F��Uv�;r9��k���{ s�$휿��S PZ�o� ��*�x�I����px[lp�É�/4����V�[�9)�"#��MM���	�������s�bʙ���+K߃F1p�,1=���v�Ji��C{�=C���I6. 3=�]Ϊ��&[���,)Y��>ՔC�L�T�y�o�,XA�I����/~/��J��Y���s�t��O j�r�E�`��YbзD�.@l9Q�K�����=e�'����+[�F^�V���
^��rf��Y��d��}�@ ��������45!<�W�k�$� ��l����"_X���ِ�HyL�S��΋A�XG�/%Ǌ��2�M.���V9ޓq��lohh[|�-rq�y�bHi��h֝с�x�亳?�z���h/z�f��SG���R2�as��X�_@a@i@��) ӦR��ft#�_q��$�i����6O�
�	�Ƕ�}�!�����9<��T�F����:�e��j���5-z��J�d�|��&BR�/CS�U8t�SG[)�g:fv���!?�E1g��,�⼥]��(1�xXg�8)t���
����2D������B�H�ReZ��
b9{�"u��2ؕ��� ��Ò�8c�|�5mqieڼ�gFm��s)w�kH+��.�z�,1���M���ڎ� ]�L�{�G����]���Ԧ��]�Q�Յ�?��y����5�ԅ�A�?�|H�D��ҵͩTJ���o��r��Yҋ�(9�پ]���^:X7%�XM�$����E�qLT2��?��d�@�o�.�жj)b.�Y&����

����w�Go����S���(Ā������3^�pw�9�VF�j�ڏ���#9(5ku�ϲ�_�_����q�6�_`˝�e�S��ɞ��hD�ܿ^7,�	CШ7$����~V�NF6"��8�㽍�_�����Ԯ�w��|�b��0����~5�����`������3�v���)c\�����V v��,H�^�|(��;�No����s���/ț��+T�?�n�Ʈ��ױ8�O��-~��W{Qްĝ��F>I��*na5��4A�c���x^<Jp$��K��@��M���ȶqx����;� ��tSQ�IykR�:�:��*PX���dW���w��ME�ٸ���ǔ�4'�gQy3�$�F�C[P�w�w�;r�(Κ�!R_-&�fM�7n��}�5>,�����N����a� Б(�I���7��Zm��p���(:�o⚽[��G��rh�%��PWf��@P
��C�/��w;�o?�~|�_��C����~%�@r�u�v�ƌoň��5M���=����)�O*�m�ϙ1���Q�������
��nc�Q����~�5����������B �^˕��:)T�oxg��A�/>�X�RC����}�'Am?�k�e�����}�쫦�}<(��e�v�� rq���G�ᄍ�D"��B��h��n�y�Ԁ۫Sd>*BP���,g�3�,;#9-1҂F���>�BȐz�,������u��W����fDI��!1��29�3����� =�Vp�U�,�O�(ھ��?Fظ��_��7ޠDΠ�������W�K��͡�P���1���A�]B61\���RW�Ƒ��xΘl	*&�I�bX`�v:$e��4LF���L�N��S���KK�� ������l\�
�i�F/�s��r�����p���L����AS�M9Uwp��]�3,�)�V����T�*�i *7k厫����#�['�I\\B援�j�j9��Q,�TȨ״׿P<�*�=��3�����"BE��O���c�6��$:!f�N��2���+�Kg L���Y��A8�һvd�0�K�1��ɮ����9�>��'%�#wA�1���NU>��|ISE�����YQiePۿ�!��i!~�0�>�LPGb��L4�6��f�KxO�oj]`Z.P�q/��0�������¬�ʏrV�LX�d��<U^���#<���dV,S�-�����R�dr%���D�i��!� y�	1�� e�A�-�,jOV�I%���ߘ"���*���olR�<iz�I'N��Ғ��{a7 *���~�GA!	g�
׶tʢ���J��
����D�j�d'��H�!�?<3P`���: �) Bj��[��|@�HtP�#�nJ��f/ Ç�,=�Yt��8�(�����e��*:�ybC1m�%��7)�e�}<���>@��ֳB�OKạ�>L��#��|auBL\~�t3��faBM�xN�@�yq��-��D�7�Mו��>Ƌ��h��!�����˯��V$��%��Bi4	�ei�
�NS���_pQ���7���#���ف�-����Y�+�=<b(��Н�*z�,`�2�~�;Ot�O4K��r�˲%5�O��]����z��-��Ǌ�Y�c^�S���$�P�M[�Ϗ��pQQ �;��P���u�� ǿv"��v�k��G������{^���y<��ج�sϕxC���F�1���$�r�G�^#�."��?2c�Y�j�@�؝�N�uc˷Z��J���K����9��Q�u���(glu/�$U$��ڋ;�V%.��X�/7�w6h�K��}n����_� w|Ŵ���٭Ŗ��.���+���2Dy��4�qX��)Vw�;�����'��uQ����6r���}Tw�F���p�����Z�1>u�	�l.q��&���|u�J��ч-�,�@�a�������X-�A739-�=q���ekx6����Z���\Z8)TL����a� R���փ#-�b�lR���OI�%���kx�K7C��R!"Y�]�,�j0M��8�G@l�;j`�#T�^��W M�8�jud5(>���܂ J�k��#dq2�ݝ�s|��X"拹$��jU��L]�'��">[�'���� �P�d4&����C>�K��HH���~�鱫�A�PQ�;��-I���<�zy�*l]�Y)o�3�l?_a
 ��X��
 �c��_�(�8���G�&{���Xq�(yC����ǋ���;̖��LA�ސ�Р�`h��,����J��H�dP۸w�0xA_=�w�ֳ���T_��v���˳� ��j�g����S��@�E�.�J�����)H�+O#��S��r!���Z]��&��"A�����V�8ؤqE��i�G6�@$�ث��G�r��F�7���my~~�`O�U��|}*���w�3|#�I��U����Z!0��aS���d\�)��6}�0���]W��ꬻ�I3_��i�P��D�Q�׏�H��"��
\R>KbO�j� ��b�u,Zvڠ�gYƏ�;I>
/����Y�@���2��� &㐯����/���;Ƀ,��e:�#ԉ�:��6����6���<�m��<�zF���D|W��2<��)5���z5E)CD,��Dέ���ն�X����L8��k#p��D���T%����;G��ۜ/!m �U�������R�j��7~����MH����?\OY����=�����?ߏw6��\����H�ڝqj�zjĴa����~���q�O[3�Y]9���,H��8�K��༾�����{Ep�Ci���	�օ��}{�O���}�1�u���&���*����[��j>P��y�M�m�L�[�\��TfV,	vm�-���{3%���E/	�Z�����I��+p��M�受B���-�'8J�������qj�^U�����-��r���ך�՟b.�g���m���Re_��4��.��x+�Gd���f����u�'ֻ�*��7o�D_,(�Y�7E�&n��!j�(��
��4-��@ǏT��'#g]$��Q��U�G�Uϧ0g���6�pV�$��QL�:�
��[��(]�Ӹ�2.k⏭S�BW�'�b��[J��6�\��03�N<�������_�m�5�WN��ku�,��$W��`� �T({8�M�63�//Y��� �����'��?�Z���'�h�v���}?��������1������#�3����5%��$�2E��ڄ5�յ�Px�u+��+�mb����qj����Rm\G���F�6�߸��n�^� >����6���1�;9�tE�4]��HԲ`' ���$1�6-�x�eΛ����$�~��$�)[�yU�A�Q(���9{�B�.�0i�(��a����T�ް���@\���[��[��p�	s�ǯ�Y�����4�$�B7�`�������2ͪ�=�/{�Rj@�����Oȸ�y>�3����فHU��r�)�����9Q^���PfK�JUФIП��Z���VN$mO����G�� "��L@�м>Y�Hm1�B����<��j#�j:�羉��3�dH�{؂ "��q6 �	���a��}�My#�M��c���I�7=�!�ڦ�3����šF�<������}�B���gA8>` ~08�y�����(�9�.����"@Xxx@B�o���,�Z h�}=oo��"�F[�o�S��$'�Ө$A���Ag�Ͽ�4&־�D�J��N��W\b�U,޹8�>aj�S�0�p�[�
q���w�t6��eY���m�fRe6,����P�_��?�CS��>��x������m�F�e���#I1�,���>I���8<���_7o9 ��fн$Q�/;��\��?]��!�����ǩ<D5�o�no��#�7��uġ�Um�x��PL/2�	M��Sb�#(i8P4��Y 8�,�# �,n�C���k����.��t~��?^��<-πhcc���	���U��L���|7ӎo�]*�Ԟ:�.^2�r�7U�~^Ișc����X_()��a�-�CV٧����'P9�|�ʶL�6��ڱ@Uۓ�P��5�ª��Yq�Kܖ�0�<�<{u@�X���{ �ψ��	�wK��E���B6F�5j�v 
�N�#{�p��^=���V�-�B���MpK�v� �-Y-�T4��Uf��N���%��#�U|N4ʝ0g�uOǼR����Mkl0�>M��D0��K�j�)�IJ�d�14����I9�ҷ>����^�I�K�6�;c�k�c�~�$�NA퓻�*�����ڈ8.�):�*L���л��]�N�T��0uo�*����Y%�|��	D8W�-�ǐC�M�z�ԪC,���J�{��u�:�o�ˑ��^,�G�j)�i�g_|���~e�t�Iuo:x��|������$k�����6��j��LXŠ]@��4O(��w�9{�8��K����9#	K[E�6uE�ҧ0<I���>��}�b�x4@��F^*ǧ�B�����UiK��}��`�)\�@i(�*zQWڛ���u˂D����o�և��v��A�Uy���E�H,j�!�B+�3R����1�ts7�
|����t���n�.���,�v�u��-A�<<��%�NѾ<�Fi8�۰���zC:��lu��Y�T�n�ݜtd<�j�YgoA.>솫��8$c���A������$k6v��g�1���Ld�׼�1���"	5�����O��9�zG��J�����t��k�kU�úb]��l� �v����v�q7��e�h�/vy� ��� ��� 4�����0激۠ESj�*P������q��xf��|�/w]���`o�f�W�h0w�u��<�w��T��zX0�	��	>���w{E�������a��:�^��Ի�*�RK��e��#��%T�AYh�!�+��#��кJhP�ɹ��T�j�-6�6o�T�N�`[��U!.Ȧ��ɘ�Vlͥ�z�%���4�T�^��m��Ͱ���r�M��Ѹ`~��8q|겮�Iڻ���Oi�Ɯjm��f󔲪R~�2|�'���u�4�¦��2H�u�&`4#�S�k���6-�#�.ŖyI ���z/�a�'+ H�P%�E��8ȳ�|�L�y��� s�'�*xb7���w�@>'ʹ�^O�z�0��W�AN� �O�gLB���8�����Q��m5�hb�N@"��8�η[ ���(�`�!�P��v K��ń,���
�=^˜��aA��9�\�f_�[/�V���?�!�E�O�1ژ�����
��,�v�g�kB����������7�ZN|���&Э+���l���d!�B��;�a<�a���NW���b�َ%�;ڶ&f#?�C���8�/�4�'���)�}L3N@�B�P%��T��~��Q�J�q�J|�v�o�v���t?�o�s�MK�CF[�q��΀D	�,��Ƭ��4�k�j��K� P�[��o����:b�61$Dj�:m#r�������Q���o&���EJn���};���������P%��=�\F��w�!4﷩�TH�u0o������zD+2]&tB�i4T<�<W�{x�\���A+$|ͦ��Qs���*���[�m0��K�x-f �)�(��qGx������&���*X�)<����2<g*��/>܌�]�(�99k��VN �v���u�*�]<V��V��G����u�Ch���E��R�T�se��u)�S)# �!iB"m�Ӂ�Fk!��6):Fč���&i/�6�hC�ON��!�"�+p:d��NZx����V��3<���TTs�*e+��.R꧶7"�Ar
�u .�9����<�U'��
nb��N�4�ׇ�C�{�49��y�*n:uI����� 
���/y��+@*כ�r�iE]J�;�M����V	��ݐ�X�l�l�t�J@���\]��&�(�]d	�K-���i���H���1#����E:��K��Ϗ�/h�+�����F��wF���go��7�"�&�Y�Jj������RP�r���ۛ�w����R���Q�#�'%�C���nMu����Y�6w�m��2:Pl�R�N��7y���LA�&?����;U���44�����J-]�����̯��N�,��^(�~E�A���wDL�+lD�ĝ�BZ�_W�be�Z��0Ϙu�����m\��ˮA5h =`�O�U���J��u1���S.k��I7�,1A�A<��҃aj7��rŭxy0XW�-��W��s8�B�.�}&�Z�	�_�x�q�<��\���lG���Pw�i��x��
�)�p@W�"�Y�=�9m�"�����g���IIfD����y�rc��R�mc3�۸�(����X �Bvዽ���c"b�`��r(��9i��0c[��C���g���cۨ~?���s&�j��D���Z����������@y�-�]m�}�lq'2R��#j�NT�Z�%�8����ŤL8�	k@H�_Ch�Jd��٣�wYA�<�۽����a��rA��,��A'����\Z-)�B���ȇ'���nh�ڿ