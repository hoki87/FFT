��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�#&��#�<����胸i�J�y-�(��*�U1�OA�7�-��/��it�Y�Mv�}˽�L�:�^G�U��/�y�
�[fz������ �G A9�+҆���
�-����2$�6>�#�̼wC���W�^���D�|{����˷�0��KɠnBf2�3Yc���6�i�f�5��?,O����3�ƞR��rM{ӽ_�W��{d��Hi��Z[X��P���J�Q�=3��jɦf���8Ou� !�1��B^+��I���J�m����t�U�Oth@ަ����d�R�0�w6���惐�⎫V�ˉKӘ'�TtU�c���I�y3'�,��?%�'���V���*,���<pA��c#����ۉ�W��I|r�亘%�%�"�`8�%�?�o.��´�&�!�<�Ӱ�E�y��G�b�R��p�`��]0�<%@7o|�y{�Ђ�H�b�NLz�{4��	�T��t�lm�U� �;�X2�ǐ@`��l_9�=+q�-��k,j�L�[Ǭ��ەEz[h�z*oo�p]����=w6.��.P�F/{J��ޢ�k[#�p����PlL�+��}H@��GeSU��=�F|0�Ϲ�S��ҽ��ӓ0�0�⼅��ad��͢�!��P�[X��J,h��I���d�2)�*���u'(˓�;����@�QZ>�r�=�x��	��b0%�Ԥ�����Z`	����T�wZ�����n�u���{�.�vޜ.��Jmx�%�.���i3g4�O�=��B鉦,�)�)���o���Jʍ2Re���5���ji��8%�Ţjq"��y~�c^�:?{�,^�D�jv<]���*�r�i� L�| ���q�X��)֌��|[�L�b"����<x��s|��p���;�֨�x�����Q�_ܳdC�_Z�V��f�5���'��D3`�w��G�4S�g��JYkO�$���M�R�/��!��`a��mjg��H��gO^_E�>s��.)B������д�����Ŋ�{bh�bMq�&��/ j���9�u;�a�빲���۷���f�g�6M�C?��\��0"�E���3�h���˙)�{x��g�$xX6h��߬����zPm-s�Ծ�d�I{?'ܔ����1����(�/�Lj��"�\�1o�Y`'	���Ǝ��7��ޡ1s������N�a�L�� ��!��D�mu=�GڠA�/���n��#���""a��/���<��^��APS<:�6�~;���q-ص�N��H�k'+�؎"������ �x�F�o�U�'��̟����k&��y>�2D�׿��qh?Q\	�J�>�v�],�Ջ�_J�_{A����^kM��<���l�Z[B)"�y�����g���s�I�S�0`�9c��z-!Țw[\��{e��nՀ0 ��3�����s[��w,�(]�.�-�]5\y�{�u��n��u=K�4�'����Q�
^rӲg��+�D�Z_��s����x�c�9�Dϲ��&�&h��v���<�3m~�����ik�2+���|(��C�`�7��~~��TJY�0,Y���Km�G9�M��.*���w?3��]��*�C�ݐ�8cu �8$�Y��]us��Њw!|R�+Zoi�*�^�#�m{�\��6=��y��I����nֶA�7.��9B0�+վ��\F��.��Ws	94	�CX'D]�>����Za.��E�1�]/s�⏕f�a�P�fL�n՘����v`},�&�Lo+_�״�9�h+h�����3�${�rR��x�B�D�	���x�:��g�v�V�<7>�Ӡ��MW[�6��bTn6e�����R�[�>��/�u��>0/���s���v|��7�l8z�&������U5!2�%VG��>>�J��d女i����W�XWa��8��qN�WķA��������ѩ�4 5��A*���4�
��@c���`V��̯���`�w�{'v\1�p@�~�����|�նH�ʷ68d�Jh�Im��켧U�����n�'��~@u�<�W��dS#k+�fw˄�طYZ�U��4��z����{_�(JP�Q�ˇ^>o'���Dr�cDΰxü�o����/��y�Q�S���d�jwu���R�|�V�
�.�x$��x[9J�w] RA�<XE��H�L5��I��7X��@��(��8Q����QP���EP\�p&�5Y�7���X����M��v��`R.�����
5���F��m��?fG��uD���_�aU3b��Cr�h 1V���MM�YB�`"F��叺����z�LB���/���΢�!��_�@H��kƞE��k�QH���iuOP��<�3����~��V��mӼT]�e�H�ʡ��ȎS����<�T]��ޒ��e�kj���AH[`;�}���(�A/���*Eg0� �<:>���M��� �+'.�0/^;_�R?'��?��]WmMp�� �1���mT��W~���m%s�^Y��	�}��6�t��S�g(��V=���M&���8�a��	�q�/�I*���2�3��Z�8���-+}�|ēkJ�8���I(��
�ձ��߰j/�<����V�Z{��M�X�7��{f���R���1 B�sT�*�'
K���.�X>ߊ��I�]M��#���@��kQ�f�९ȵ|����᭗$ֹ����m�p�Fu�][K=N �h�m��TL4\]�]�گkm8W	���zd[���Od�:�H�ܐ��@��0��fb�ࡓ����}��r�Z�W���(N�)%$��4�8%X{P��E��2���%/1�]wt,3��	7�?�� U��h��>=�f�0d����Q U�.���'A��w?�1}�b--�󬄥b,}�{	���합��*6�
 ��I�H���'�3�Q�dd{v��_��.�R^��A8�#��0��[�[��vx���\�i(fP���C8�=�ˢ1��<���k^�ىj��-��>?�F�P�i�Eh_�V����>Uk-m��qը�c����6KIя:/�G�帻�ַ���Уst]	8�g��XW)7�ܥ��t����C�b�c8�R'^q R̟XT�j�:��I���L|�x!���v��'�ni�B��'K_���>��uc���o�,�i�Eՠ�XNKΚJU	��0Dȅ�#{�C[u���ऺ �����3_�s��<�A���iq
��4s��1��w�YS�<M"�����Ai0+�*�K���!'��Y�=3Z|Uq~r>�N:�̀堨���u��'d��L�]���2��8;ȗ�q��Z�����t��,�N'����RI�/�b��P�ńŠ�#�U��S�a�n�ydÌ~�3ܹ!�q1��N�QN����D�>�g��]O�C�Ը���6�Qʴ#� u������R @ikݑ��i���i���p1��vP��@I��g`��$�&��ͣT��l�M���{j�+�㋗̮��$���f�N��P��R�*@`-���Yݦ_�X�5�������eP�rk���2�O"��܇*