��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#���������l��U�~�׏O����j9�PY���`T���x���s����uí������P��"��b%>�1eτy�<�gܰ�N�Y�	� {��I�ɍL�ݫ�G�R�k��Q�!E	�5E��.��:�͂2��y�m�-�.E��i�����YS�
��@�H�ۼ��nD��Y�l"BU�.TԊ�=�-�����q���Ǹ��j��ԋ����tr�a�ٵ�]�b	��%�ɔe�)rYOjX5;V��R�������M\�	D��ҏ����9c=�Vͼu��Ro�P�Jf�tRvsY��c�"n�XO��	3g���Q���^�Bʹ�7gQ+Г���$�-��t�8�����A���<����l-��*�|d�!�&�J1l����9^��V�| ���a=3�^Y3�C�@�#�l�Q�����I���"�Ap���-l4d��,�������8�Ո-z���#�����JD�C)�*�ߠ��)�5+�,t7���|��O�_�%�V�o�,E��U�r\�ken6�k���u�Wc�_��:sd�J��URm��{�;޽�Æ=@�l����:I��
+qH9, $�h��:1�S�:�^�bmes�_>��e	��t�RH�r�{� Pl.�fkĤ�l~Vr{2j�jL�~��l��f�w�j}L�fb�7݈���n� *B	*(�s��^���H��C�:"�HTi��� �Uu7K:�{�jN�I�狖6�M���1�N�=w�OR��s��X�In��A=
,�
�/?�_����hC����ȥ�t�
�:�]�`^��(Q�����'��.�Sm`��O���ōȔ�Ge����ۿ�Xh4�E/s��N�ߊ�}>%�3�TE�� �4�,����L�&d��}���o��8��4����6j�y�$�h����2��s`,1�p,�||f�Mf�`��~ڹ���^��C�J̪�+ODB�܊���2��+P^�]�j�HM2C�|_�� ���8M��).�~��[���K���E�.��fo��C�]�"�w�'�����L����dIdR���B�}9mUԧ	�����FU�_���y���y���4�.�j��1�r@,��[���s�*I�S�C��K=�E���*�({:}!}�����\OF�zj����07��p�PW��u�3�-O0�1���6�ڡ.\_��м���[k4̂�G�W��$�0�K"�Օ�1_��?����*#�R�k��3� �{[ƨ�B	���]�4�zp�����@�T�����p���>�������J� �����t� ٿ�9?�dI�-6I�Eϼ�HlY���W�Û�K��ba�g���M��� �[a7�m��+�_���Z�ʗ�N9������8��װ��?�^���d�ϼR�N>�a��K�=�bw�)HȒ��Ss:�4,��r�R0�U33�U��&<���+gZ�縸��k� !(Yug'N�Ju� h�B.�Y�{�>�Z��19�X�>��b�&Ҋ�ƭ�4G�<���wY��|>�|��7k�I�5��y$�㆏�;�.	���r��ކk�`��&J)G��;R��;�|EKĦ�����D�q){A��g��?%�n�S"�t�#��fm��r�c�H�����0��N�	�9 WC��\�	
�= ��ι_�)	;e���
OP��W5>Ih�����C�/J-��s_�C�P��o:�)f^��#N8�L���Y߯�+P:q`�����I�*� �FJ���i��o����G�Ow����G4��`{���獳<^���������70%r��*>��n�M�KT����.t�g��4HƜ\���VB���>1���=�ѩ4o!��Yq[.�4+�I��с�3p���AT�W�)��>X�@���\�I3���5wYBג�~��|�>S������ EhqG�?���**����H�)�#���vK��iiSܝ�:8�Y.r=&�)�G3���5D=}�+�����C@�m�)���$#��'�_Ҟ��4A
�޸v������A3mZQ��-�ca��Ƌ����S������Ʉং5��%%���r%  �6d��@>z�8^%�S�� 4�Qxeo��T�L��b�M��&���9��"�Jc��[�p�w�@� (�Z��v���^^��O����2��E}hv����b<2k�P�F)��u����1?A���HC�ұ� ���m&>�sF���˨ڰ�bjYFjC:�ր��k�����(w$BGH���+����`k�i��d�5X\`n��~��J���;Ԣ���G�6�54k�AE}!)ű������MK����F�
RZ�yJQOZ`a}�`���� I�;"�َ�{-QɄ}��k�}?�q��{����)��,sln�@/�E������(��iBځ���|9\�&��
A��66��xW���d�o�k/�m-G00�:�qf0���-���)�U���R�&��aP��G��3/���#LQ��^ tK�
x����r$o��,R&_@�z�J�#Rn��d�O��?���AN�T�X�я���e��m�_��F��iW=o)����J����Zx|���f{��)��0yù�����LK A�:�o�r>���EƜb���`k�Ǎ��!�j�ѥݢz��s�"�2����;A�I��R��lx)�[v���Z���W0���DUc�r.yU�YXvG���iU��/�7��mb�?����I�*,O[b�۫:׳1W��m]�}
G��$���	�����זn�#�*5��1�J����4��y�w	*�ݸ��h�|�[Y 
.о��u�a$�����s�/-˟E��[
ڗ�,V
C3����bK����2@=d��PВ�0�t�+V�"�����R-��X��'v�����NBs"λi`�����7NhQ�43�R��jW�`�WS�i���A֎�y��D��&��(��4`�qf3�m�"�Tq�,�H�iK���to��H���n0��*��1�8��:i��3�+ ��Jus��h�������ϱ�ȞX�4p���Q�뺄�q1CdB���G}�A������sy����/f�9�/�=��kg�(Z� 9��j�!X�A)�^�G�p���r��&����"�z��o��_�1��j��Ը<�8�����Vj��e`g!��ΐ(�ّ�y\�N�0&�6H ��+u-M󙉡��/M{��׸tBǥr�K�FeA}w�t�r�>D��p�l�G.Q_>��m�lp3Q;b&P�m]������ �lg<g�+��J�����"�w�5�}�����&X� '&x���-m��C'9[,��֢H,��+����{=g0I�،8m�8v.�4�9�;@��A����Η���8)�3�f�;�f�ĉ�d���t:�q(��@ ��LO�%�����OD��v���Tr�02W��:8mҍⷀm�4�PM]�:5H	���С�(���f�o���W�љf�KAIf��L��?q#��n��Tz��
����2�3�IJk�w�q��7Ox���Eo�������Y����iJ�l��0�\�+~@�=F���8q�c昴��W��z�눾�:;]1���=$S韋z��MW�Ƙ5�σ����鵀��`V8�Z������0ι�ƪ���\��,N)�2�0�S��^g�I`Z�X$�=$�8��-v�����ux��,�n���K���?��-U<�`]+�L���X�;3��%dظ~�(�o���U�/1��@<��kn�^��7^�-��\�Mi�%i�o@����ߴF����9�Z�Ѡ-�<*=�o�y8�R��G�����E> U-�$>g{.��3�O�M'�a�T����ڂy�����~*i�{�Ǿ��4�XdPG��Hx�Ԇ�*��&Mؔ|�7�-N��P^IX�e��؟�t�eY�d�>���f�H6�.ҙ1����7��S鯧�ɖ�&*ny�L�v _���j���2C�,��9����y�<�tU=Dh�e�9VU�T���f�CE�Eų.Fw����T�;<Z@j�5P͔Ӡ����^��[���X3s�1�4pI����� �'�WR��b#�wO��i<OiB�l�vi�O��};Y�w0#I����,q�9a�k.d�����N��#�2���xx�vA����_#m���\�	��13B��Sw�>J8@�!e ���hod�:q=���<i�Z���+�67�I$T&-�q8a���ZkF,������⭕D�y3%󶊙�����kƨ��˛р�3O��ң��x|g��n��<p�!L�e�`/W5ad�q04+�q�e� a����|��"�U�",���[�{��swoUUy6$�VL�6!S�U"ֹT����(�m�ڵoN\͊�V�C�q{e�����ly�gFL�
�5I��@ �d�=�S�F ǩT����@�!�^�\�FF�,h�!��`-�#�b2<�/����,�ޚ}��'͏�b��5frߋ���Wה�}�/���ޤt��Jː�Mo"��ѭ���xU^9%�MTv�g�g#GrO,j\���K�-�P����wg��**�՘�S3�-5���/e��i�^(�q��^�a�Ұ�@\�])�O�*���N�+P��<���ë:�ćQ���Y}�H�r�pI���&T.#"'�r��R/�ma����F�����R�@ıD����#�(8p���Fe}�IXRB[��衷�,��
v݋�,�t~��/^�~�vG�B�ڋ�ϛ/s�˄�H��M���e�"�R����%�Q }��ou���S߯���WG
�:��5f/��h/����j1����WW����5��!�@�<I_����Sݙ :� ������3�n$+Gf4��nC����CئG�#U_�ey�ӱ�X��I�i���q�R�:\Q���N1���+�5����s��
���//��*$s�;5��yi�Z���n�]���砨��O_��ʢ.�dvi{Ͷ���Q��P�4ls50�0�~��#;E�k/�����/Ux����q|��/Q�Ef�q�R�L�(}���7�o��[��kd
X2�>�Z�;[2�Z�<���I��9�Kl��b����^@����HR�İ�I�o�<���3fA^ v�����'����N%� �Rqvq���n� ����p���%���V�����5�h�¡c<�	��)E�茒2��mit3o�p�*e�?��N���SQ���4��u]&��X/���Z����f;-�Bw�yj���O��k�2��L�!�hwڴ^fP����&U��'ȮG:e�/�H�y9/!�h���3��S(�Th�洐^��lj�@*B�ِY�H�b29�0��߲��@xRH���V��l�CY�;��5�9{�7�%��d�u}���nT}���-�b�ޤP��K���O,�5e̥��J.cn��Q������m�f����(M �ߐ�BJ�}j+�}�te�sz��P���Bmq�dM���A���T����q��JW�������f�͟]#I.���_�]�Y8qGތ�n��"Sn�[�dv����J���%n "�����w˦N�[t���>������G"�`����[�(?s�sP	x���v�Lf�o�0���Ԋ�ύ+��u� Ye��ˋ�z#�;,<�7�.�*��8ʼ@Q����]rCf��J!���}����M���j����b�Ms[!Q����q�3��[I��j�o���!r�8�ˆgnx�қ}���]�u��$.��o(���P�I:��#�`J����|�Hdo��"S��<b*r_�6���\�|_��|dι�v�(8�t���''|3#6�f*⁜w�9e����$M�� ~���~N��I�Gn\�y�2��:3�c�n���o�.mV�I{����F,f��w�#���W!Z�z,_�0a�����*�iVc�	N������hkeg��6$;,̯t��$A�Ed�Xܴ/��*�Gb�ߺK;�Io� ����IZ�;l"�u�{��K���~I@vg�BiZj6	ē� +ω����ôi �:����YY�_��{fJ;�Ҝ�V����1��f��!�$2�v�2���vW�z�[�8���f=q7���5_�(�c��6��+��MQAn%&	�������b�H��Q��d�
a9�L1����W�s������$�Hii;%p<*���߫Icv����[� �;V��
���֯n�("�A�2T5'�I9����	���v�T7����B-���� O�S΂��C`�ཙg���Yݔ�]#��AY��]�%/�P=�)�N�|�	��Q�7.��pQTv����D�!B�.��������y��Rf|��<-���t���!`#\,�kQ�3�N��&+>
2�3�Ew�3�TÿtH�tn~#������U����?�Al�\(chmqJ�}Ub�AC|nQ(^�J߄N[�a���2ӡ$>)7��|��jC�k�.��'4i��j#�[�s��Tٍ%퐁�(���I�튴�<t����ǰ#AT�pU��܎�(�/�@+���C�h����2*�.���x��~p�}z�D���������/���9^U:�zG���I������yLDw����/ޟ���d��ߣ9�̆+[}W�5X>mR�N����'E/��Kea/�A�ZR��s�*.4k�����B�Rwo!��f�=�2��	ܱ�R�@��Ru���������1{__;���N��y����U���%�|.	�=P�l�F��&�=Z��ۖ<�v�RJ�0DρwRMq
'R��F=`2���̙�r!�i=�A��_e�+��%��x�����G�SD��>Ϩ�2�x�|L?_x�Ţs.��*�-He�����<���L���'~��,��F�6��/7\B8�p��z=,��5*^��^�2coK��TInyz�E��mg���)3g҉$�ɑL������t�$h����
���D�qm��fDVI])n����h#�G�]������[vY���%D��k�&Q����9��٣F6�C�V�m �3��?��e�q\kX�U�]q�̦*�pro��x>��QB��/����٪����D%#}	���5ٿ��1F;>N�ߙ.'���^y'�f)\����X�C�~1��2�8�� ;���4q�
�Ib���9 �ƍ�����@��b��ɹ#;?��w�tJ��V��#�-�4����>�o������s�����P(�6t�eq������R.�ܩ����U5sg���	D'�Ͳa��\ܗ��|a��_��1�0G�W"��������wK8���X���ct���e�r����6{̀�����8�M�y28�o���ڽ����[d����zR�a�|$G�_b�x�Cci����J4y֬:ͤ%����/�]2�q�K0��?��)�Sp�K��e;�>C���ޑ��t��d������JO�/R