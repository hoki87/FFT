��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ��������튢V��@��3tv�x]P8�^��#W�-�D���L���s9i�
��8��N�mF�<̭x�f&B�Ɯ�� S��w��zǘ��!頾�U�ov��] ~�	e�|�"�mo��8T�M��j�</;�
�H��u����f<�XC��y��d�F����������x��<4 �����{ҩ+��RF��avQ��#��Թ��2kZ��t�l懻�ޱ�/f�4>���FU/;�f�h����kɩ>�gt-�j�Æ�SɔCV�:��2�(����2�Za���GWX����v՝Y8k�C��Zv���g �[����&m������sN�:vūEƗ\C^d4�0if4QT��X���p��Xm������ �
u��cdX>1ލ];M�W91Oa��q�� 
�y=W}��V��)z�� m�D
RR����[�o㸕;�,���2�t�/�^�sźD[Ʒ���.�s@G�A����2�mbu���y��|��5-��ډ
Ũ��'�+�b�w��I����Fr�~�բt;��
D��
��0��QEu�8l��r'Q��PW�N�M��h�b	�$ܛ`UJ&�<=H��9!�65ğ��|�(n�g�Ө�r!P77�w����ruC�1�6�>D[@#��~�Ɛ���&��h/��sL�Jk�ԧ.�_�p���,��O�##26R$�:}�	ԫu6>x�rl;���Wd%{62��Fh[$sm�AH�+i:P��UZ7z��u�0bΒ�;-��p���pŴx;�AO.�wl�m�$��0D�����-���z#�*�G�7jW9B�>����Y� /09ڝ�puQ�=��D!j5�D#�cJ��^��@���~� �L���+~��_�a�ֈ�
�0C��&��k%�u��x|Xp�%� 烼�h�aOu����ϥ:ץn��?�⦢A;�
�Du�X8��A�Z��q��1��Y�T��Y}���d�) ��)*p_ʦ�W�c]�l�{x�QK��i���	/! q�OO�e��0��o��/��S���uga�*��S���Y��C��7zL�9�����D�"��M+�a�	��Q
02��!�>�BSn��㯿y���.�>��P���w�_`�04������[{Ų�`s&k�@K}{�S9qXAVh	���ii���m_u�����R�- �ޖv�c��������ֵ�?��'��la-�p_0���r%�9��V�{1܎��z��b0�f���1,�߃Ѫ�KA�hF6��J�Jm��Z�+�j)<�i���\�_A���<��>�첏�m��j��!��EC}���l[��`�<��74d�i�(f��x�6O�`�^�:X�2��u?G\<�h��oBE�ƍ�osQff�3>���Ƨ�7���qc�3s�����N��ȯd���Onp��V�i�],���#�u�Uz��-`�G{�;Dd� Z��@��d3��;���Iʢ���A�P(~��	vm�8"�{�Ni@��탤�٩Lzg�ngt�R���:p�`-���ib9�`�M������2kn2��n��:-��o�-�r�k{u�����WN��JR|f���"�\�<�@�KF�we��������:�PG���b�Os>�=�Џ�D G�~@W�6!Όwy�G�W�鵳mzܱ��BE�\ϺA����=��n$,���V�Epyɉ����=��RdU �QN���x�F]�#��f�����d��ΚǏ��p���~� ��Vn���o�$��U�cni��Щ!<}�m�T�<Ek��/��~)��G��s׸S#�@@󀕚�^&�&�j�y���fe�;����� ?�Hԏ�rHuf����c��o�	���x�~�m�Ѕܨ0����@�#r�� ��SF3����?e�!d׸���]0W<��4L�0���7���ۇTzֺ���^ç7-���PsWD�y�Huv�V�c�?����]��6�mX�v�/2�aM2<o?���>&3rG�-B��n������Pr�u��L�]�k����Ӌ3�2�(�rX��k�d��\�2�^�w�~�D ���,K���'�hڛ́�1���Int��s���Ė��+���9j
s��:o\�'M�YC/_+�� ���T��g��u�޺�6�	�쀕�dveh��UԕO���kv:�Eɠ�џ�3ah*Cc	���to\�\������TSB[���0�jL�#�R�Av��ȫ\6���0FS��W��[PKk/cS !��������{Z�k�f7(|F7�8�v�E,���d��¸��+-�by/�h6���Y-�k(g����^���<1�k��"�X _	wY���'-�ZI�y����%FxUʴ����g��`�B��		��M��3�vagԥj�R���\��n�7!�����NRm�z�����"�b�|��������I�DViP��mX��sr[��̭������D�{n��9��Ʋ��~׵�������;�'^�ưڅLF�<���?�*�s�%�O��Q<б hh�k#���ǯ���-�m��b7'$�`���M �$u=C+�dX�+	}��Y#\�c�֐݅����wYU�1�E�UT?�q�oЁ��DU=���YK��N�ߦ]X:�,����v�2������#��g�1�oV>���vÛU��+Z��]3`j�洴L%E����\�:��o��=��5��W�O��PI�{}���ȡJ�G�2ք�zaG�b�g|O!��>���o�@bB���In���.���
;9i�6i)�1v�SR�5C	�Ç�z�}U�V� �MŊۢR ���}�/�|�z�9.}�;/=��di��P���+N��N@g�����t�a]=רar�AS��Q��X,[�x�E=����s�p�~���,�z�.�ڲ�Qܝż/�f�4�rJA9z�ΐ)hx�Vw�O����w:K�M�	m�ŧƾ�<G�*�!�R<q�}�e�-��6Ƈ#
/�ok�X+�Z�+k�'ق�����޾P�X~IV!}1W:���K/�F���������4��O��WYs�ـt�Xz)�� ���%�f�Ҕ�`�@����:Q�] �4C��ںi�{"��nͦh>[_�'O��Ku�8���ɥ�����i�"O�t�����������K#ҽ(0<�K�M*O\-؃	w�@0���)MK��+�)q�	m3��������#"��]P��4�mҸ���\�ƈ��ܪ�k���VUB��mC/��~.����o��kC��m\����oYŸ0�'�H!�r�bb�R��
��_��NUGx��O����:f����]��r�� fP�5:n�,P!cd8�p�d��~�eiJ���.��>��7�4�v��V�&��m�!I(��~���J�Z,e�,��'?���4����4���h��_��qF՚�Y�
jx�'�Yd@q�[�Z7����_xC[�rU�"�)�(m��4˧�(G�sTZG�)�r[J�c�R�'e��
�'	��fWTV	b}����F89���oﶿ��Sة�z~֬�R/��4�Frñ\����i�4�1/;�S��:�FM��]3���T���	@��(�W�](�j�Y�p5�ʆ|��"4��B���v�G������#*nDd ���*�����8�z"�Di�#�*��a�mMn�Y䨷�xy���؅�4[�+ۛ�X ��$?�ƩF�ǐ��ގ��� � 6��ݗ�!f19Â�N6[�>?��Q��w�f|<Ft:d�@�����ݷj�{e�>p_�$M|���̔���t@&�� �U.��D?6�H��p>(^k�5ũY�E����������Q����z&c�.?�*?`��
!�#�/���\N BB`؂F����5�Y�p$�����4�T,�,��I^R�\�l廗��I�ʎ�S��W�:Xa�w����	H��ܑ�.���꣥BĠ28��	������� ��)�ߤ�]IƓ)���	�Ff�����{�M2*��I^�$|��9�-��6XJKjXk��
XBғ,�+$I�����J�Ŧ��P���{��`��]13��X�:Ɓod�/*�?|W��QԢ�*�U��d�B/��!�}&����ݱ �I������?�dp-{�--*Ec�l�k�/������s���7e�:4H��|�v�?"�ڝ��6f54/eM�*�ݘ~f���H��{�'���P ���C��A/� WH���T�j��qtH����}�c������w2��eֻ�C_K*���1փ��+^N�?��7m��i��]��8����j�Q�)#�ܹ�[�#�͙Ke,� @*�:0�����(u݉�hv"�$H��ء����0%@��"t<Pw���פ�]��y�ݺA�2YNu���t�Y�)f����9�ZU+���f�s��GG�@�$��1�6e�������q����N�WVX0��s�y�]qn��cin��E��6�WīD9�phR×d���vN�D&�P������a�����7��9Y����Q�yy��7����y��=�ǔW����(k�̩��$�[M�~G��_�OE{ V5�0kU�������P;)j�ZL�O�Cz��' �!�����ղ������V�4����w��-�Þ�B�G���u��������������(z`�K��$+F"?Td!-C��Wƿ)C�ܸ�M����q2���)�C��n��D��6� �Ѳ�F�YP�%�ʣDLZ6��w���E~�Z~zL�ӎ�go]��k��E��䰣_N�|���!ܣ����G���O^33�?b"�T`�¼{��W䣠N8	E^���虽��`�:ڤ�_�%E5H G�VnWX�Xg�$�^��s8-:�,���t��C�.�~�KMeX����Q��N�d�\�ȡ�Ǉ����'i!R/o�nz����	q����*(�H�/�z��F�yϓ�څ�{����D��R�(&����y����'$����Ī�?΂�K�~~4)f@����/6�48��[�H��fsU$_�N�z.��?�d9"j�j�H�א�g���PR��B�w�� 
���������"ض�݉��9�Kdԧ@�I���ژ�e��O�zp�I�f*B��Yj�  �>��wj��?�Y�7A7g�_s�)�)�"��J����Zk��� �~t�d�23M�j��
�u�f��%a���Z"��0�%?�1���G]iy�P�%�57 ��'Ɩ�X��jIA�֕��y�R(�<�/��	�wn�<�
,^�<�m`\��6�
PF����^ı��T�i@�K��v�t��U�>�`����|pj:ڲu�B��s����ciж8xj?�&� ��|��``}��4����l%�X��p�{� �E�+b4::��_�?�j`��+�I&���U���fg'0|1��g5���	�
OQWKʬ�ǩ1#�Ѹ8X�b���w�u)�!N�M=���j�O.����~��G�K� &I�2 *L�֙�&iNF2O0d��B8��J/�C�hڙ��?��%W!͸dET�Є�>�˞S���cP���|��O�e��,�$�/�'�� �H��FՂ�`���a]w��R�U���}U��|`�؂`z�֝�+q_���žeoz�}<�}��)��m��z
��V����.l|7t�{}����&c݇� Ж	v�pi�pw���y*�
�C�k��Ë\ݗ�՗D,>�K�+� D_�1:r0�U6)��oO��d�;t8�2#,����:	T˧%�R�w���ZXIjء�6f�[��B۴3�'RQ���b���g\5�AU��o��� (���Z���g�h��������1��|��1e]��	�$��)2X'#R,(����r�I��Uz�;o��"�J�L䨶�!qԃ�)�*�<h\��V�Z.���\�$p|�y@#.�ݙ.�m��ӡf�i��:�31���ߵP�Ǉ�F�����t��eB�I������!=����,����wU���C��v1a�o��k��-���|�r��'�(�C��.Z���B{�S���c���i�S�^�7`	���Z�OP��)j�E4æ,a��Q�
S���HH��1�[&�W��Z�_���
��-O5�V�g0�g�J��-C�e����.�Ⱦkj��W�B������3�$-R�j�p2����*��"��2��\I
L�x6��վ0�:5�3$����X���%
a��U����_rOHA�� �u�`�x&�ռ�t�#��Z��2ZtH��'#�0	������-����F^�K{
�.	H��y��R̢כj�$B�v���Z�Ē�8"տ�\2^u)�j�A/�9�7�ͯ=L�1<w}���^������%�3��چ�(3sgX	�I���e���0���t�C5NC;�
pP�"�Oݒf��I�����byܩ�ۈ��5�eCg��YΙ��):�1B����Wg�t�:�o�#���Y��ͦ^�wm j=�0��(ח�&l�Q\(�{�d}��Ӣ�Hj�s����L�
U�H>�!�k��:�!��*�U�n�5S|�&V���������Z��f)
Byǂ�1Y��ehb�����!h*��'���H���d�j�P��^���4^m�8��B ��\�*
�2�Պx=X7H��EA��{	���5M5�-�	
�]�%5����RX53hR�}�cǟ�Z�gD����*��U�f�*��'fa�^�E�z�;�\�����\W���i=N@��\�)����̎�O���T���K��z-
���-���e��/��U��"�l��"̊F���d���]�<��l�=��i,B:%����&i��,��	�2ţ�r��e���0�7- h�\�V-q۾��'�c��=����?-�n��}魜�C��r�^���"����0�ԉ������*Dg�R!	�T�BɪC���޵U�K)���Z�[u����`�Z`7�bm��r�+�s2��۴��ŀeS�����p�g�]h�nԄT���>��Z3��3�L��|J
����5M:L���Wb�L��#[#�WJ�?��^VkJX;$�3+�{>l�����J�(pu뢹.�	�e�	CEOα��FFOUa�<3�3�Kl*4C(�g�<D�+���W���a\|�*kT��t���e�Se$�����щxz绳�Tm]k��������&x��"�j�/8i�h��>Y� .}jA;.c�4�^�m���r��-��;
��~c<xx���Ћ5���^^���.*`��W���0
pd� ���n��p����flR�]�K�T����~�����BU�A��whS�S ex�m�R�I�`��L��"�TK��ݨ�5d�|2N�ioZ �Ց�5\l��U5V-�?�-�oߞ��uO����*<�@���6ezv�u6+�������A�Cd�'`!�O#<<u���6���3l�"�LA�V�~o b����ڼOE]�=_Tǆ���h%������_����ԉ��=,s�a9l�7�u��b&qY�k���􍍢�)�۱�h�X�5��2����`<rnC��E��� 2�k_�]� ֽ�V�ͱV~���?ࢮIM,%�Ɲ����Q[����W}�}�A�Q5�}���@�-^��z��������Q��!'���3�|�of��Q+9s��?�υܭc�A�z��0�*��JEkoB-s����b�2�Ź��h���✮��L�'��"���k��nQ�>�A�{j�LD���ա�d� �lŵ�A&�䣛�D��jWaJwҭ�Z
7�3kwp�V�����'���Q��Yh]����*�,�ǜ��������p
��^ce.��'Iz�?�P��2�n���,�qi09�E:�@>���)޼E���ᔾ�	5�q�pG������u!��o����9�����]]}(�f�����wz�u��R��I*u��pYڌ\Ҭ̍AF�u�����}GZH"��&�(�:_�2���Q	b�`h�s�Q=R�hÞ�D[6�LN���[z${+��9�$tte(������Ip+��΅v�Ì�B�k��������N�#�\�Q�9�C<ay�^O��*d$鸖͐�	[��5��Ocч��Rs$���}���*8u�S	='⩍���M{����8��
��أ�l�� ǒJ�F�q�5��!�lc�����	��c��.��#A8�aR*G�<���kNh�Z��
��������PƵ�@s����4Z<�ʓ��*
��q]؛����19ߐ���=�&mf��U޴Cҁ�{{�Ƴ�Hf(F����Zr�at}RfSmt˚��ݹ��HE�6Y�Kmm�s)(W%`!#�U��q�+��e-���	�b�?-Qq�-!
��EZ����Y:������C��l2ء�(�{O�>�@���XŸϼ]�~�
�U�����_8�	:.x1E%�3C��@TL;T�FG�g�F!F�h�kp������D�x�N���I����S��'��p�_���e��V�M|[��&a_�'!�Y�E�%��;xgl}���w��&��r5�ĳX�9�tzR���4,�-#f���Qڢ��H�ZFS��ֳIv=ɹ�3��"{���]�U�pC�!*Eߥ몁I������D��`�i�m2wL�����{J�����/�sD8�6��D��O:�t��ʘ�LP�(��I�<��d�ϼ��6_�w_���7�6o;`��N�>2%p��I�E���t�dJ�.�S|N�yvBX��cj�6����4�N�tt9��68�B��Eϛhz�̗nf�s<�<�ˡ0�t7�}�
��e �?�z̤vf{+^dS����Gf�J��.:.��O����o�R�&���_j+���zb���zvc=�q�
��&?�E�k#S�n
�l��[��rW��x�n�H�2��ѝJ�#���i/Kk�~�Ц�[��	{8�[��EE�+��?vg�	����0�6e��8i�mk'
��[2�-�M�T��;�r2���t��s^颫�+�{���9}���Ȝ샄�����]*Ƀ�_R�~F�7�K>S����m�0@W��lʮSSx9E��q3���_��fڞ�-Z������!�>r��M��V���\M��rDy"�2�OW W�,f��j����.�窩Q�^�ˬ��9�ԏ2�KԧY�ͺ0��2��!�艅������W�4��Ӥ.�\z/yg���Ւ��P��X�u	Y���%�t-��L���I-���s=�X-�ʸQ1��d�ç��+6�=L&���ղ�gbk��/!���_N��j~Af>�*�W��!�j���p�a���_�4��1��$\�xO��|%�ʐ��^�|��I��q!O����k�Ӄ�_3��b���ҟdx���^�0����ӽ<#ە����M(Y@��G�f�Pc�8�ĥ��"�X2��.�8�o�S��k�KۿOf	)�PvF��K��&Q�9�D�K��=����\36�w,NH��a(�*�c�]p6�M%n�φ�5�3e�G���U7 ��a�54���D��,����;%e��/����!��`�SqXզ~�k')o{�l(�ҏ-|!�;k�ˎ����oX&ڛZ'�3���k-�~�ESg7h$�)m) �th�����ĸ�0�7z1-�B���aė��Les�	�|J�*�HÆj��p؃<�3�x�1��p|<^Z�}o�H���O����N�;���x_���Ս�;g'�i�0�����DH�L*�?`P*��-���]dZ��-x�=>�>��]��W�.�?�����1�ᴤ����#�W.��"
�A�,�؅Q��p;G5���.&z���v!7+�E�<�U|����Xc�3���)��Ł~�{����0�xl�ZFw�4����	���w	�}�NiqMv��x'r7�)�Ĥ�<��2;@�R���,�=ۧ4�թb����+�b���/Q�E�NM���aq,�3Uw��G��h��2RQ,'Ψ�>P�0�m�Tf����?� *w��C�1l
�;���ď�� (9���A5M?���)�˛��[�+$濰!�������D��&p4�`\� ��w*޻���{�p�u4��	eJ)��«�xQs�k�ӝO*Dр�<����藊o�ʥ���
Qאs�o���z:�����h��NE�q�qm�%M_Q���':���k��=m����Gŕ����]T�2p���f=6pY�0z����|�z`�]D_T$�����T��f��[�a)U؉Γ-��j�X ��PQtLCK���)�s�s)����0M29g�Ju�:EÖ��p�v{x2ɜi�wWS�X0^L��:b��Y