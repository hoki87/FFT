��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ���������,C2Gz��K�^�F�E�D�ir�Q����;(�h�Z����l��xA�C��2�ṗ�A�5�j!����~~	C��X$I�Q-�����E1*q(��1��&�Luj�J�'�����.!6�A�4�@l�iw햧�cv�ρ���g�%@d~�ʖX\^�j�s�3��6�Z�b�D�!z	�-��}����/�Dfs#ŧl�q��%�
r˩�]����n�*rTj�$Lkd��cq<!��q'z���WJ�3�{A�Aq@M�)㋊��U���:��"�ɖtaMR{ۜL{��)X��'u
>#�����[���-�Ɠ5�#
���G��J���A��[�*`h>ʍ����{>�����膙Lnܩ��=I�DWO�����!�;�Ս;]�>g�:�P<��A^��7�nX�C� ��X�VKlSK��$Qcb�ʀH� K,@�����g�c��,�B�D����J;U����;�٥#�|�ľ:r*�������@��i6p�v�lc�~��Π��H��!����N�yKc_��M+�%s泔A@���3ov�v'���K)O�!���s�������d�^�Σ�3s ���:�Hi_5��+��ջ]��r���)�iƇ˥���o��m,�@�z�����N>̛�F�q	�`�I�
�f����IBz�g��v� "O��9�����Z��\���,C_)4���	��/V�3��u��:�
`,|2��%���<#~�^d�_��i����E���Ǫ�q��L3��W�[�90���F�];h�Y��yu��
�}E�D#���7d�>1��R��Ï.%�`6'u�g�Y��)�~vÓ� *������1=�2^���������$,�y��)0�	���wX�N�oy&���6J�V�h�U�ӎQq'ģWPw��G���Յs��f�������q�a.?f��f�B�.�)���������O�q;57�w*�A�סG����!
��xRW'�8�j�i.���\ع�.hkjR�i�=M���������9uκ��teA���nC�<�B|9�,��HPx�U¬�N��3(��2?<�!;�
�J�E�Y�"и�윾��Ʋ�/.����0�/�XF��`�{�~�$4v3f�R�WA��k�J�D �q
;�q
 W�⩁��W�wmi�o����%�QA�0@Q��,��;�g�m�����ᖸ�z��"ӄa:�N"D~)�����Z����p5���;�vV��!Kf �]��Z�=_`�tֺ���bH�ސav�Z����Ud)�V����>WB
P/>�n~��u��� x�V���R�[�e�X����5{u�{XL:)U�D]:З��ޤ(T8��5h|^8���fs B�ӎ���V^�Ƭ��T]G�GvN�c����\���K�Z-t�K���z�Έ�
��U�ÿ���=^ 
��@2.Z���㍡���K;�>�/�Ң�{��E���A4o�"s���J��z�$�����@V��9��XW* ��<��n?��2M��v��;��`��\&y�
+��?w�G���cu������01��ގ�1�Ñ�!!�z��n�$��!�͸ �ZQ���Ƈg�z+=�ޭ�T��cջ��b���������n���*}�����b���=,���N�zv�ȭ%��\&�j�8���q��gKU��R:;���k���&6[�u��.D�Jij'HW��*d��<��o��+X�8��� ��}�C����0�b,��Ɂ=��h`��Os���ܚ}�����������D�}�	��_ɏ<���0`��³��686�YB��#\p(�y��c�C�̩@��)���F�'s�i0A��c�U��ּ@$�^z�ϻ}��p���/������2
���}@]�*�im*�I�`�16�R��2t^|i��������բ��]���fv�w��Pe0�pM>����G����'��"���H�*k/!h���f�Q� �5v�"�">H�~�C���'�F�}P믤�O����e��j�C$��$T�z_��?���4]�o��5�vKX�ȫ�Iq ������a�6��`�
S3�b�x?w'x�Yk--�N��S��%KCe�)%�+�3T=]�K��e�rWg���a�����\祥�*N��|�9�Y�	����OK4�K��Xf�v���7�Y��A�r�,�T��F(b�~��c�I��w��2�*L�6��b��9�=���̺��?-3:��ۺ��ʵ,Z'�.81�(�0�M=r=�9�~��`|���� }e\y r!�P1�j?���4�e"���CHM	�A��'�?d����L��IEH�D�{#'�Q@�������+�M/���Y�J�Q�p�)8��j�ZI�C �,N]�ζY�v��Л��n��[�v�s�,+�>'q�aZ>X�ʃ+'��������H����s�i�~m�x����]o��P��X������qL� �MO�y��$>[	<\��࿔y�*��~�6�Q��jW�o;+�N���F�lb�KS�}j񚄨����R��W(�f��4=�WHV�~�m��ܮX�m'�� L����/%�l2�>ߋ�]JN~oq��hM?�.t��>��c}�B8�B�<vHiX��cԊr��5xh��_0����"&8�Ԋ�̉IM�����.xeRNn��#�,y����B<RZrr��)��h��Ao�X#����:�I����w渖&t���nW�e���UOckg�j�IL0�ެP�?Pk2�?����DI�H�,SZ�&X3�ˠ�!~VjΈFE�0��]z�������4����;T_�����ÄYџn�����Ѫ?�8��Y��A5���7�tG�Zq�հo��x<����0W/��`�'t�wV������g��+�2ߢn�R��^W�Z��q�U&��&I�����ppv�0���p��1w�vIfm&��c�3ݨp͝x%v��M�����5�A�K���+Vn�B����i�EL��
��3@�_����0�c|�'�,49���Ȅ��O�Z�-��|
��B���6��L�8�5NB	����������G�l*��$}i8f�N���9��*�>�I��Q�U�d)N�S�Vu��.���A�̃���X����NBnXY֊�"I���U̟Xu!���A�J{9i�	�$A�lǏ�P��q㷛ws3�J�x�3(�@�����`PU
'R�� E�ox<բ�Xm%z|o0'��k}�T�2�]4+�v�	�*�t��'��sB/#��U
�(`��s���Lȯ+,�ƶ%��Y� 8=��F9`~A���x�J�	�=��d[��"��?��RG_���>/�zS��]`�3ӊA�Ot�&< {��a�\6�ǵ�W�EFO����d�=�G�Y���N�ѣ(BR�VܛN��By�Z���Cw�L��q�L�$��vXa(� �r��>9fqΕ3�	)w�`S��Oc��p�7㍯�'^%{5ċ����=Oq?���x�3�&��@b�K�v�2e9���U��6]�`��C��n��n��eMn�/�j���k�>��P�|�A�4�6=X��t�x�4����Rû4YV�/�u+�<���}e�t����uń�h&�M��B�&h��� [ڪ�뭌��h�	>����/�2d���������h�?�z����A\wn2���fF�p��	M����ߵ�� v
H.�ˬ��s��t����}4��|�8�M�7.%�:��`�c�h��d��W�gd� XL�2��z��r�*s�Vn��*��'��R�X	��M3��P�!E�|F��+&}i����N2�m&�q�0�����aj�X���,1b�qY��/Y�|� �0 �4[�T�5������)9+�@��󘞼��A�D-
/��6�!�w�δ�\�hk��{P���K>\;O��Wq��1;�E2���^�@' ��L3�V�
P��V��]�Kێe��[?j��L���n�����Ћ�W�9�˲�M3H8��V)����D�� ��2^��q��(�)����T��|Y�܂Y����yH�KZIpfu��ˊ�������{��m���NPch�w���|���ƙUT� ��S"Sʛ�ed���wmX�{.��P���u��̒κ�O��!�k��>$�|5��ίg��F�wm��+}�ߕ=!vFfU"�궏w9����� 1m�ڬH��A6��+�m��cv�Z�?�ȿ��r���1�젽}d�o��lYe��>P	����Q��1V�s��I�}�9��g~�I�i��Ɨ�~A����E�]�'�З�c=0#����Ub�7�|���a"�( ���{�&
����u�:�����d��Ff�Cp �:ա�&�4x@�Ran�.�z����->e��t���FW.	��|"`���8�a�Z�͛SQ.�s���Ct�p3�׌���s��@�$W�7����k���(�L����#<�u����]_՘�բ�Ȳ�r}%T����j������������Ai�E�O�/)u�q�����⭹��>9����ۢL� l��N���aF3C�5Ī�ٓH���\�68r �\?���,���]���	r?���e�X�$��׸F ��~\�mb·ON�>�ՠ>D@[.�Ѓ��)�E᜕ᮞ�ʙ�
�����I�_�ړm��<6�,E�\MG<�sb�aB�����M�$�p��r]�>���i�����L��lo�q�!]/�lo�.��O�e��� �3	�׹'4��?��m�7 @�`ս�Rnn��z�����(ٺn��
�,���0��J^�E��sEd�?W&�� Ѳ���QQƭ�
�P�v�z.N�N3>(��M$�N�j�s x��ޖ�{NՂ�0�Z[�\���%[ހ 	��X�ݑ�Q{ɽ������)��d�mCF� 4��1��먫�\BP�yY.���# ���;O4ס����2�Y��"�d�X���0j�S��X����&�/H~|���-��f��zǿQ몥�ߍ��@����֛�.���X�3	t�[�E_vj�K�;��q���8�l�q9�|'FA��]3��XR�FZg����M���*�L������/H	�f��/\o�4_(��'�7/AM�c��hiv�3��
�ubL��	<��'��1��視���KJi���Jjm�Y�M�h�*ᲊB��c����'��'�o�i�}��'����a��>1�c$Ƃ6Cw�
t�w㼁��N���������j =?��^�[RD�{8[�	�gҍ�<��jf��������R�<�JRl���T X%��
ϋw6_���kIO\�ԭ��0�7U�jԚ�f�k�A����6MmV��~�u�!� ��y�6X�u*���l�AA� ��xuՉ�e����k�*3���S��{Ix���E�8��<pm���=�E��>������R%,T����y�y!NxGV�������1����ek6=���ϻ�ֽ��U��x�-O�/M���Q��}�(B�}����'Τ�D+�������[M�$��]�Y��E�y�B{j�Fh��m�濕��e�QM8�N���n�!H��t.' ���:������d�O�t��2hx�\��m��5=IH�.4��O(F���rf�Yv�Ʒ�}�3"�8�!4�q��ӵ03�:Slԕ�w_��n����U�tLkֶ�s��9<W	I�=Fy��ZFt��"�xI=�v�"�lh'�P{�mm�C�P���f�ed)�+�,G��`M��K�flH[<�1K&����Y���3��-�r$]��|��������\/�#'+A�������i�����h^����:!O�k�36�D�"�W.�A��Z�n�VϕblL���켎v ��Ơ�4�E:j<�᳠E6��~��>�<0�P�'��[���怉�-�a�p�\,8�O`C�� �0���Oz��ޛ����[��k���l�� �?�!��Q��	DI��F���*Ⱦ�r��5@KEe��n����
�#V� ����U"�h���0��5S�)���t���4^3r"���	9�-B^<*�4�����(A�9�^��gН3��4��lH��uc�C�u��� XA��tT��`����{���-2=�QA"2����`ٵh�M�!:�$�Ѫ����{�2�A�Z��/��p�M��L>����Jw�ȃ"O�G�&ZӚ�ahz��9!tff��A�
Y<Bw��Ħ���������j�a��ɱn(�&4KH��-g��&-���E�]Cvp���Y�	��>�:�u��ϲ�=*Xb�t�=9�ѵp�����;E��X��/1C��[|��kطk
}Z��b5Q]|rܞK��9,e�4�6l1I�������{[aK��F�wF%M�\x�e)�d�ea�u��|�vz��3�k��"��R��J�U�" �yS�@'G��*��ЮLbX&%�liY�Ɩe�(�4�%� ��i�/�t�g��^7���E�u�9��]�Vw�-F�=8�� �H���E9ZPć[=#�Q�&'L�3%�+��׶�7@����IY5i#�r|�1k��󨱱?=p|P�"�F�s/RY�~ȿ�	���M����``2�D��s��mz��w�.��;UK��N,��e�><ŕ(���<�,e�cP�����<C��`D'�)g�- y��&ig�^�	��������'�O��~����Fk�G$9`��ƥ8�o�T�aW�����7"�md�K,n�R(�|;��l0®K��`�<C����ذ���>o�)����',��;g��6l~�[_LК�G�r<����&)��Cx������]j�Y�/@������\ n�MӲ�1�ꊭ�+M�w*+Oo��`��(�zq5uVXs����aV�.G3`2����iCGn�Ko���RK����%ϊ�	 �m�E�^�p�eR��QM�d����I�u~��"֝\^�F#�T�|��[z6wt��������P�L�z����,S�(���|��k��e��¿����²�B�{�T "L3F[��3��|�h}�%�?��DB������^`S7I�%��5���7�)�?��)�� %���X���%]�ʉTe ��#�WQ?�'��k��G��t\!����?e��������X:m%�q<�M��?v��g\�g���'�빎fC8��$>M������cU�s�;DʩC4��8�N
�BR%�l����b.ё;���4�ldN�����R1�1Qs�g� i.�wqz��F�/�%�m0�=�-����$"���U��@��Cf�H���4�s����g!�7	���� >s�_�]���m;6Z����n�I%�w�����#[���.sk�"Պ�e��l�:���R|�U	��9�ҳ3,&�\9y_���������d_
L���o��5m�PdZ��$�`�!���HP^cT%$�I�XmYR�6B1���z�oN� C�zL�i�
Ku5�5r����5��~�!Ƃ�Ǧ���y8��E]la��+9�L�����4
����z�q�25����ry]������@̾\u���
F�� ��(`�0N�.����Q�¢U]�{K�JSSb	[�ɞ��Yk��$�\d�%̶���5.jM�^�4��\�k�Jn8�-�Aveߑ�l�K�̩�~�2���̓�V�����&@:�{'��[_tq����|q�$�"�aΞ�5dB���{����)�<��F���Ç�SVr�����uE�F��WK����?���7���8�������Ԁπ�*���on��-o�i|���u�ۻ��/&&d�v#��c'�?��q��<��Ԡ�G9���� #|����ܨ���UT��႘'Z�;�0�!�lb�2��[�"Z�d�r�[7��ݽ�rw)�s��D�U�X�_�3'�䝐��N��=\�z�E�\7N�[�W�3`��2�����/�/���9L��I�L�7PD7��g��G~��
����I�TU�k�6 5��6�g�l�Vaf:��ˋ�O�
��e�Br�Z�kU��4=h�&W��0|&LYb�h���6�ș�y�6"�X�o^-ǁ�����>�!V���c$lW�"�es,�p�(�n[�^W�qB�Ӵ�C��nB���s�T᮵�Jq�*פ�^]�~n2 e+�[�vS��y��`ۼ)>Ȑl�85y�1��W��5}��7.аG	`�$p��������
��|9A��勻����pI��k�?���y��3�f��%@���J�����&��: ����ah�����2�y�����^+��K�j&!Xc�?Vޭ;Ɓ�^b`m(Pyʽ9���1�;���5�������U[%l�&��F�g��qfۙA�X�F�={+�OSJ:{�b�Б�����h�\�0O�_oʑ��>�k=W���^L&}f��[+(������ۂ��Њ��;��Y\���y�5*�:iv�K�|�Y���I��mD�m+Q�T
O��yV�Z[Nv6�i}63o����:���cޱ���ft �н><�6�rr-l����P�&����0@��>��bCW�Y��pdL%q����[u	�n���M��8�2#��0J1����vA���؜i��Ҙ�;�6ЪF ��9s���|"�F��L���&%���V ��8�Ũ�Xy#D\�P�vm���,����Q�k$�@���4Z��㗢�[UcR?@X/!K]{t�2$^'%laO�{��!��wj�]��	�Ri^o��:+ĤDKL���,��Џz��s����˽�Ѐ�av����Z<I���lI0?��*=Y8С�sf��v0Mˮ5O|/;�/4B�v���+q���o!�<!Xկ� "J����I�f�����X���iP��|��1u<R󁛀��]���i�H��[b0r���.^o�h�S���R�ulv�*N++κ���ښc��^���� ����Q,<c��)��:P'~�f/�S����d�S,ܗ�ٵ���e,�%o�n
�`��u�8������ǜ"�::�����C�c���*L+���Dx8�
�UP'Xu�N��3�!�:��i�/M,I���I2բ�]����i�-��@9���4M�Fz\�d�P���N�1�ga,�9�t�kAp�.f���S�@L�*��M�P�#�cy��t�p�p����F�Td��~J�@�NX~�W$�l��d^;�n�[5�Lh0�2�	bx�@���Bt�u� �^NLԝ]n���-��Y#�����_�2�Ւ��*w�g �ݑ_��w��$k�!_�r�< ə:�8ᑮ�.i�@�5	������f�	��/Y���f���m5�4;���C��)I4KP!6�9��^rF+&�2�鶥QU~���Uw@,�k5s�<��D/D�kֽH��l1.s��:�7iUk̾���$���pKG�������0+� ��޳~����������IQ�9���8�J�n���L�u
�A+����D����>%;C�o8�M;�c���v�Tm�l�G���O��d4��Fl�u�ʀ)�*��F�Y��ؼ;@wǛ[���Ia���3Ë�i�@��ٚ�s,�%�(�!]܈��aZ`ӎ�a��_9`-�w��I
쌟�;
 z��XN���4�˰s�ď��Ms:~�R�O��\3J��ۈ<s	���Ҵ�ϮW�
��9e�.Κ��W �*�WUEm�5�WYr�����e���O>�@��6I�W~��6�3� ���C�E��[#m�{��d_��GH�5uv
��j�����k��.��r��JQinDy��������y���d��7n֕	� ��:�K,2rכo���[y�L���V������}9�G!䠗�6��>��w�p���+�3�
>��\�D���4�r�ҺK���?� ~�ZF���n_W�١O��[F$0��i]��@�=YbqDƭ��AcX�'�iW���δ�>Q
Z�/�A��������]/g�1�nHJ�t3�6vSg��}��,|�{������S]�9�a㳎��)+|A2ӰFN��a��r���ӿ���ٗ��, �5FĤS��z�:�ŉEȀ���O����	���$w	1���؇�!@ؼ�εSQ��L���3.��rE��`ӹ�j�(�\L����V��9M@�nQL3�/�	����n���x�Zq"��H�O�R��bu�f�iY�����xs4e�S�:�B�v��s����A��=��F�R��Ah��������%��*B�N��
P���%$��v���/�x9��5�Lݛ�|�iBK�����x�>�&�b4��V�!�͌�#�G������+��,q���h�����i�a;`�ֲ1`nM�B?n�[�e!O����	��χ��ir3��D^v2��5[[����I��3ܒF��
��g��Jʫ�qA%/���Nj2aio�g�g��T�Q��&,2%�~P�$��z�
 PG]*QѬ9fG?'�kN8���w��Sdb�����9U�t��9Ak4U�w���t,���3B�©�b�;�b�\AYŝs�㧱u��������
����$0���W_a��?Qx�5��S��~�	D�Ӻ�BF*HO$!4�v�����V�1�����>=�X�R�0�a���dJD}4��^�+�L/R�Թ�4S�Qb9�O���.�4�"�'	*a��|3�_���N%J-)ػ���N���Jdu{ؽ���xՒ$V����M<x\L6��.L�ݼy�s_�F (�t�僋.\�{sBD�����i���S���|�8��� ���i��jW��y����dS��Y�@i,�����)�ߑn�C�dD���Yo8�f賃����';Q�O?޺Fv�0��f�gK�mQH�m�Q#1J�3E���-�v�Tu�XX����?���pn�*q���G��W��ҚЫ�R2lQ�����c%�����{�y�y��1�[��[���x*ԁ�ьÝ�把�n�:ࡌM�`�u���1����ňm������&I����&�"�e�t����5_Rm!�X:/�����y*:���VuE�k��C^�*���|�d�7p7�jQ���ⰾ1Z�j����D#�"Υz̒��E	�پG�4p&H=�/xk��.2���	�y�����jdڀ �x�"C�ZLC3��:�O�;�53;��Ϲ
,AIuᾐ���^m�P����[�����J��3V���P��]-f��g����R���!���i��޿��'���$	�]v7�5a+��w[�y�yvW���Q>��V��w?��ϣd\N$��uB�x�f��q�
�ҭ,�:��.'QFc�q1ь� �WᚎU�"*�qZ d ���/���OH�%�����z�²j~Ƌ�kN�'ac�?+��R0�ӆ���Բʧ͞)*,��
�X��k4��@�$l�$z��	�w��NV�X�9ˀ��ùq�SQa�3��ϗJü��<�y�V&�XQ����Oxd)���&F���r��=8����^���o?FTsK�5������np��ǽ����������(`�;r��R+�H9�8���M;/�Ͱ���`���#�P��ς\䯝��<��n���>���|Y��dde���P�CO����"�!?4��1�&�e�p#�GtX�� ���ھ|�q���H��M&��ƍ��F�51;9�9<��a��aДIh�&��r�����)�e�#!�+ځ˨b��^C�P|ٚ�	u�Yp�#�a�MJ���+��+~D�;�`�A¤�)n:����3�j����x�LaP��ռ�K0�����9f���r������M4u"V�;����EPU0���u��ŅQA�e5gk>��@)��tf���������;���f<���g2�>u�Y� Q*�2�ݓ���xbko�eBB�f-8����N-���Рʰ�b�%����L�|��|�{�F'?��d��Etoyw� ��
~�cޡ��������2�!1���x�؃ur����4:�L��H��8��.֎�Ye�2ӎ{��im������S�d5fקb�MA=��V�,i"�s���u�ݖ�#��?R���?��Y��q�s��A�4/�6��6�Ȍ�Q®}kKfm�WxZ9����~J�o ㍲�	��K˺�g��E�[�|�H��dw�ǦzL����~������5��!]�}�âAQ�u���������=�h�v$����Z�/�Gh�%����ʕCTB�.���㟐i��!ҋԖ˙���D�M���D����H?�[�5�ck.�X!��1���2���u��SGOc �݌���}޿B���5b����<�
�e����S&̏��ƜuH��1��6�g� ^�������͌������o�R5�-��>P$�fMK5r����Y�n����q��K`�Ca���z_#l"�Y��Q�A��%�t��,*�7{��c��h�c��c3z)!���q�/����2���&�54���>��USǠ��Ƭ�.D��i/�2RbXGؠ,�N*�~py�МRJ�A�F�eq��b\��@?��r�S�8@�I�ـ򇣭y_:���^t��V� Z杝�wD��	��F��\/(���(�|��@���>�i�Ʒ�_1k�(�m�4T�9�)j�^����9wA�z��ܪ'���\m��+��,P�b����ꃟt�_��1X���DgX��=`�Al�`x�(�~��=9]�ȁPJ%�$+49��n�: *.	�ۄGN�>*�X���GǤ Fhl��:b�t��}X�ORN�O!�F0 ��f���'#�	�|�h��^�����o|ds��T8,� ���vX��|F�6��cl�;�]��@�A�&�@#�S	DTmUòI��$-
4�k�@w���͡���5O�P	������ؑ�@W4�~��oB�-�>�,������1�g��d�2��9a"��~98s����iξN�X��·p�*E�YKjV�ėyw?y?N7��t����З���{�V�Չ�Ȅ&E�ٟ��i�]�a��Y���j��և�H�2�[6���O�6�^��e����9u���d���lt
z�6�BĪL�ù��]v'��p����Ss��Ƿ��X0w*�H��!��������6���T���H�5ոai �u�G����fh�ËaGgV�X��~v�>͙8�V���ot�wv6
JW�"f7�h|�9 �8�	�"����f��U�7���w�(�����{����C 7�=����"Tn�䚥,�$�Rӛ�����Y����I�x�E����`bl����O�!E+�W��߹(�����&D;��*�x^f̽�LY��bL��S��4-&MG��Ǖ�Ģ$oR���/c\0ɤ��6_`�0���?	A�?;��'x��2#/ap���G�$�mEz�b�Z���M.2i6���~b_����N�dӮ�u�0�H��YC�1Hy��HS\��d�KH�s@������;�P���>׾�&�%�g#��'���\��GK�xY����,�H,�-$(\V̍�8�	�c`jN����	��X�#tI�wd+�)���e���9ud��5������
bK;���*�0��S��@'o�O��Kt�{A$�w��w;{1>ˠĚ�7���LrT^� �a�82D7$��&�eNq�e ��ȔĊM�s�;�։�k*��B�Lm��V��|�wzH>�-�Ug/D56��^:��9:�ؐ��먆�s� i�� _V�P�l��5.:9���6�Ǹ�-3�t�Y���X��@�6V4L1q�e]qX��c�^�=wk&�'E@7�]����W�.k`Q�g��=R�ʅB��EMrQ��U|Ԇ^`����P�ף��)����H�<��u��C0�5-������~hEx��.�96��F8S"�Jf�M�l�t��uA�52���.��c�ĞV��jZO��9|�����\^���1Ͼn�H"���?���:���1@C�dg���;M�Sw/�������9 LRQ�u7^��}����iD�(܅Ƌ�\�����>��:vdM�y�5��~鎱�޺���w�h����O�I�҈��AP�3�j4��:���,���)̡�-1�!"�p���0�E)C��!-��3p ����1c���H�ן�������tnK�ߝ���,X��bq����So|�����İ?#�㤃�T��*��ʣkS�(��~=�@x�\�ٴ�KFy��0�_V���'ɱh�L�mm�mcL��S���tw��㨩�(�e��:�}��~���Q �%ɺOX������u�?��\_� �}��q'Y��M8�լ00�g�DX�s�wn���庌iH鑝��8�u&�P.R���p��/F�FQR����r�_��"�]��&�ݺuPe*:��OU�5��Z�x_E'"����"p�C�9`��{��L��%��;�n�1`O	
�M�%�
�"_m�jϴFMu�r�^4^I�k ��D�����K�F��O���02��mzk_�8M)��2>R�oR�����3{`���L)�W/�o��'�c)>4���O�5�"�cۛ`O&��iL�S�9��}���98�9�0�ʂ���w2V%�c���l�'K�.\!N$�f��*4�\�?��Bf�v?��)��,�r��\�Y��{dw��u�^��\�����z^Y4�T"��>������2h�1���C����Y6��|�g���6�Rݑu*(�?�[�w��.�Pj=�z$bM����e�����-�	!���oC�����p�����I9e�4�ӄ��&�X��/ꈧ���f��
g�ʹ&~�l�%_��mď &�n�j����"p�4 <.�L�����<z6-M_�p�L�ڙUw[�#���P�[������L�"R�Az�ڴ��.z�1ʹ�����P,�cR'b� <��*���Q`%��ȁ�G�$�3�s�b!�e�/�/-fOPC�R�	b�4t��{�����r
�>=v{���]WlM]�R�h؁LkErC�WL3|��g0�xǉF,52�|�]}K��b���1�"Ñ��̘��gS��>��tF�BszU�zm��������jo�j]��b*B](Aƕ�o���L��ʭC�_r"[b/
�֏|�+��co�����i����̹K�Y  ��:V�޼�?	�c_h�H��s���W�|S�O����o�hPu�^6K8��t��ig�����ȞfK`
���9��j�1�8�NDKF��R^��]ྐ�@��lBzڧ�:���(`�ы�SRS�+�!�[~�U�Эrk���\W��V>�G�խ@�K�;���6Y�f��X3�ml^l,���Y�j�kj��uȉ�h2�S8Z!����E���b~�0�S�agt�VG�w��|S8�彇��^,�{O�흹U�_(ǅ!G/�*J^{ń��^���C �Ԥ�8ݱ�,J�Y������N� lԋE��� y@��#9*�R�v�f�����d����Β�����9HV��l�i3ҡ�-�ӏ�+fSZ�lIO~vB�2I_^���c��&��*���k]�����ݔf�,@0&F�����`���ikA'�?-ǖj���e�_�;�|6Q|GBR�� ��#AV��ee��{0�G�16�~������@���"��,	(��tQ��D��T�R*@�&���Eh�K48g˶)�,�""z p�>���=N�^��0��,��./'x�&v�#�]�Y&�!����5�-�r��ւ���$3`�V�=5ǝ[�xp���N[��0n�x�+
���V6v�m)�$�M�.+GՎ��5�ЦM��Ԅ]��Cc���`f���po�D3��)?-�K���$���2�8�%0��WRH��mǏ�y�v}7�0�~�e\��V+���eM2����U��F.��^N2��#��?���gyr�D{rCf��so�ʟw���.�]]�|PS��S��_u��F�pA�{0��]���?\�~��z?���1�g�Ĩ�y���Ż�.I7��0Oj {��D:?� ��Vj��'�XnW��ǂ�y�ۣ���:�� �ܖ���z8�����nkea��ˎ���z+�Tj� ;Yk�z������O�N��D2�a����m/���A^�gv�n LGK)h|黎�eԃ|���x�m8 2sH�}u^\@�dS������T�`$�8J?��T��ְ��1����v*\�x�N_�o&�j��i4S��Ƒ��������`�Bʳ	'�}�~A�T������n�W��Q�1�Cز��=6� o�Ch�����5�п6�ejC����bR
���aQq�u"��O�u<�Tf������q=
;x^�}�ڈ}�Y%��B^F1k��w��#��kI��:DD�7���l	d2279�'�SX	f�e�"�73�'.��Q����)`{	^�*�I�yGW(��Z�l�I�Tn�&���m�IBJ��a��'�^�ܒ6�m�i��h�v[���	�!U��_7�B��V����Mܬ]Rf�1���;� �FD��7�|"�.�w�?t �"2��O����b���pUz{��5�M������XZ��E�f	>Ҹ�n6����Z���C��Zwտ�������	B��`�����h�#srz�@��m�Us�Q�[�ђA^��f���uٿ��A��HT�hǈ�&��Qy;!�k�D��a$,�n�pָ���@�C���~���F��-��7�[���Ņt�i��ν*��2����_%��@d�����F��HTu&U�������W���р��H�-͘���hJ�/���R��=��������--�v8z�aV��I'�@���:��Ibt�'��o���D�jt��v�� ��Fq�К�eP�̢9���+A����ނ��ьܟ�G�����T��T���e�+�2�ٛ�`?\J#�:V��D�)�b�Z�;��)
���e�⑗���gc3t<��Z�`Y�ڵW`}�����?��⦳��$����&$5��X6A�/)�٨���U[���I��հr�"��Qǉ,wR?N�TZ2ٿ+<;Qw��©�z*�i�0����5������V�
5�=Ź�5��=A�󿕲'��iS��G�{�4�N����GR����}&���EQ��  �E|
��%N�z���c��0��E��v:�1�F��"nቺǀ#	�k��� ��B"�<z�?l�&P�!҂6����!����V�<C'L�ka-~{B:Wq�W��ҝ/)p��@��O���S<٩������o�&1v��܃��� 
]�)Q�0�KaC]�������ZE�>
Q�m���)�?e�:ț�#%�髄b`�[9���� ��~�����q�c��;{I
�j��~5�B��M�5!F�f�[&b�Zթ-�+ʤ�_����2c�lKFP����ƿ��O ��U/,�S��ڇ%��Ax��od��;\3�ݟO��(6{��o8���	�!ŷQ�y%��c�P�@!bN�cHI ��n�j����B,	�G���W�-H�7�י?��AU؁�����+�[�&�p�]5�j�:��ы�n�>�*������i�+�25s;��/� \��ޥMz�hؾ��<�y�Q������@�Z⧆.������3Mt#d8sUY�Ǳ��k�b��_��a���r�/�S��y����{Y���@�.�R��j�]P(l�cAr��5���E^�ߔ�E�n/.��9�8�����l(��>=���q���1	
��> ��5�;ة[�V� �D�FJ�(_-ׄ�4��l�HDnc���TMH}��^�6����vһ��G��T�,�[�e��y��KM��xi�l3K��~c�*�[a���A�h�j����T�(_�";�.,�I�a����]LW���s��z��υ��"�~Q$*v(��P"���0���*Z�×w�BB2����"�_����eWJ�KU��%#|�ͦ�Lcu��&b4����EQ\NHį{��Ժ(��0�$"Y1v�l�)	jPw..D:^5��j�t�P��Ff�'~ov��7�s`|������A��l�A�K��	Ն��X�Ȳr�pq�٬�v�u�zK��q��p*ҝ����^�����3
�(�I��>���IڃH7�QF����th���f�"A�z�9E�_�gpJ7�����7�!� ������i\�ܼ����WD2�b���h"�`Y3�*G.&���*��yx"��\�Ml�Y�%I��/Bj&Ɩ��0��_�P-\I��.�M�~p��?#�:�3Z�/i���[����wg#u�QY���t�;�Y��v�p����b��1(��J��ywr��y���fl��{O���vI{Uq��J�����υd�s���\��H@
%5�Y�Vl~�BZ�)�|��=��D��c �m�8��˿t�;���	" ���=�m<��'�w5I�d��	���vW��y�8�$W]�g���[w1�&e�=��e���z/��a�Yο�ho%��Eb��f���sc:��������&�7T�
��'�O�z�z&�u1���
n�`�ި�:54��LJ'SE����&^X6��[~�'�L�E-K~��ܑΚ�,
�(*y=n��Y�?t`��wG(�(H{%pCsH�	���M�`P�`�N��sϬc��|4I�+���h�����=�]c2������L�f��pr��ҷ=L��v�VYU�r_�Lg�aZ����<o6�S
�!'2t�����9�a>�'f:�W) .���^�"K��l�����Pp�o����3���(����S��f�&������A���i���̀�W1�0�_&`�G,+d)���nMJu������?�C=�?<�rx>Ŏ5����2�X�5�u.��l)IG՛�R[K?�WW�ω8�r.��y�{�?��__Ē�����+���B���M��ھ�B���˫��8�U�Ky=�px-"r��i�|@+v�bZ|���H�{��n��(V��6ըL��h:^ҝ^�sq�k������b�*0�!u���e����0L����[�\�?r�ģ%t�h�k�j�hK*kEVπ�[������%O�3��B\W� >�l�|��+�X^MR1+T#��z@���V+�1��>�/0���h�:Ǧ�{����p�|���f��o��Ų��N'ִ2SyF�sMɊ32��M�<f�+
]� �/H��[�nl3!�S��ã{��[F�%a�l�������Z�$����8�֔'"v�+�a:t�#|"�j�z �؄�q�n�KŸ�����%��Q��xE��b��7��u�S�p����!�m��k:��x�#Ȯ�Iԝ����	��Ǽ�$~9���ϐCdJ�k�����!Rv�mpI[��y�6�*l3>�*�F�Ԛ@�SN�t�������W�'�C�
&g��C��R��.a�1k�
�k�A�����{�W�4׶����xk�$��V��������S:p4fYV&�Fj_{��n�>'2�eRi����P�p�B� -h,*<�LSt1����~�r7Ƹ��U�(�[���v��wƽ��|��E�O>�� ̘�u?�/�@S-9PQ�>?����|\��i�~��(�9���������wۜ���3��cZu����O�h���7�}�J��%e6�Υ�!���%O�Bw2� �%��q��`0�z �9�>J
)z �X��� >�A�+�
��H�L�̌���!<0�7 ~��H8kW��$��YͨPS�G��d�c���<̲3G�ʃ"��{�~��p4*ݩ6���=}2�N'%�vD9��>
�tgȜ@������h��5D�G+R�My(z�rb��p����(�&��	贇Dr�˸���|ɿ?����`���c��O�/FWR|�\'��x葦�����ɴE�^^Cza�e�I53 ��fȪ��7���,Т ��_�^# ��*���R��ߣ��s�n��#����ki�&�>b���`}a���m��TX؆u�꫌�7u��`2X�bng��h�uq|��'1Mɝvk.�~z��[��0g�μ����A�(H�X���^�c&����۵OMW����zB��&s�^`j�+�����ǲ����JL��2��[�A������lg5� �iU� E݊�f���p���|��BT��W�޹�p�b�Ԋ�QU�1���W�Y���});��F�uD�}i�\��r���:�HFʂ�(�K�8�	��yg5w0���My@'�j����JV���	�y�_U�@t!qJ�v�[����d�#�{�훊:߄Q2vլN��eX����_S���`��{���QBX?B�����h�Y�e��֗��\��M,ƌ� �f���7�� ���S�IˏTQ��u�`�j���u�-�{ܠ�U�g�Pö/nb���ɬ����Z���"81[R��i����O�- r�<���Ǘ�B�㫧�Z�x�6��ꉈR���fE���=��qhh����y���6=�G�M�6 Aa ���g���f���.�66���ծݤh���N�:B�T��&��+_�gcJ�A-]�}�!tS�BT$���5=���(
�%�䃺���*w�7�.��� I�%?�l4�K�� ����:0�ԍQ^4e���2�?LrǙs;%��Q�Q?O�@k��)��h�B���u�t���(��쮠A�%J$x2�c��g �Q{0�+ ��y�#L�8.>���x�
��W)�2�&��k�l�h'6fA1H|U��R?�L��0J���D�
���E���wI��B�&BI �Idz� �kV!�Q�GS���_��i�(��_�ܑ��9�>=��v� EO�zT����er6
51�𨽺�EId�c���}r�}~4�p;��\�E"�Z	�,L59��(h�B8M�a`aR��V�<< ����@�ܬ��`T�ҶpT�i�&��&�������¶���A��6%�<x����T?g��dT�JJ��L|DL>�[	`E �)�z,K�y�b�Ja��z�&��´Y���D��ѠMT�:��R��U�qa��ՍK��c�O��jw�U�dP�eXU蠒c=��ىz��O�][î��~��n����|iM��#�_ǂc��_G:|s?��z�8�p����a��R�X�M5�dj���~J��gep��C8҂����UVf�;�# �B��x�[�����`_����MV�{Y�i�H��u��"�6����coZ}x��t��l�{�T�7�z<gVpK叴z�Y�=�mʂ�YR��-���[쨇���7�; x���f�Y�C6�b�q�*YP)�&�$�yE)Eo����<��n|�)#�Z7�����sN`Dcy��L�@.E��U� ����m�U]��87_t�������OõZ}�16�B����+�
��fZ����o���bN@)\'�(�{n)	�	$�:�+L�����ʘ~����ɝ��1�.q.i����a�g��An�>���ti�H� H�h	ì]d���ެ7>ҕ�\�e!��g-�Vg�bz;_w[LxbnX�H��G�0�:�Vu��>1���P�3~Nڹ޻��U?/
jx,չRZ��_�i�\֎��m(u8�N��v�׿�*�K�(�#�1����:��S��]b����H�WX�2��N���OrR-�a�RpOX�E��H����1��O�z�X3!T��`���,e��#�'3�ޢFBK��~����e1��M:�;3�|`�Կ�K9}de���;�z�8���W�Zg�W�N�L�~C���uE`���5HU�Z�;o�&$̔ed>�R&b���4�y��CT���0��H���^XW��Yaƒ�6�ͮ%����Dj%o� ���II\�r��7��ʷ�a55|���[[~6c%��4��d�Qp�բ�S4˜�:���uH�gE9�?��T�d����*��"�1 ��j���bǋ�.D��j�\�.��m�F���Ķ��v�K�Ӷn��ʣ��^�&j�ڎ���e^�t����!`��:�	f��8�	IXQG������ v�O����g���m����o�-.�`�*����������闩�5/����zP�T�r���䰴V����3�-��9^=hRQ�i"4P�{PFۇ^��6F��#xz�3c�o��^K�����U5�A$��V348o�����K� ���/0��*y~�pMoEc O����l�%���Ĥm��}#���Yx���wD"̹ p�&P� G�)W]�ؤ1��q�O�����)32���V��'�;S�������JE /)��˝J�{0��]b� hKܗ/6j���/�PN#�X���cTp� ���K;ɣ��.�.)�
c�������3��M`��{[sAjk\zh�n�IٯZp)!L������g>��ƭ��I�,EOHdN}0�1����*^���+���R@����A/�3����*���!�{S�3���S�rլ42ɯ����M@+���$��3���{�7⩡L����J���z��qI��y蝸�dL��u�|�&��/�7�QiSo��T��j{�=���_'�aՂaE���Nm��yE�(d�׃84���;a��܏bCY�EԤ,�< H�Uv�\"��?>5�a�����S�����U�yA��0S����rX��}{�
���Ǵ���դ����m�D�*���m���&���<� ������W�L���ȥ�M�n�F3�������Ml�i򇹕��?2�!�9z`�֎��){�̼mj�#�'��m������4T�a�	�n��5HESR$ƦŘ?�F�5d�0�6�z0,;jɳ[�̺��D��P_�����F(N�Q��2����><|˃�ҍ��qw�0WVq���oz8S�M��{������,�}��=�9�(#su)Jy�S^Ps�}]��e2Д�RU|Ȭ����"��fd��n_}Z�{E����>7A�{����^m����䪁�)��^�޸O�������`�}홪��g�y/���&N6�5O��AV7	dG���)���~s�/�{�㱔`�, dϢ	��>1��+��l����x�K(`b�S��_7GF������d�Q�l�4:{y_�ڡ)�6j�益�ٳ�C���R�̐Ij�45S�	 ��Us(��t��jOR�t��ٚbr������]�V��e�����E��W����A6\3s������F�D���R/�*�=$Y�v��w{� U�Qn��.�Ň=g���V�-���!C�}���2���dm?�XɃê$�i�.�p�1y%!�M��AOJ[�@��2���`��)b82hL�]ђ��0�p�ы`�)8,L�ue	O�>�@g���5��Y�f��ˈl�1������ �9�`�6�f� 0M	�`��/�����N Z濙:��ef.Y��a�1�!�$b��t^�G�DC�\�LJK����.)q��dyN�6��+7c�( �b
=�j��zz����T�������ej��u����t�H�3�-dd�u
WQ���$A���B���J)����>Wzy(U��|��~�|"������^ >?���oM�Ga]aQ���E1pG�1��L,Q�5��<�3�ǯt� CgJ/^ďz"\V4"�!"�dfGwC׫��6����m�i�v`��m���m�[L<`���[�1�xiY����ֶ/�y�p젽��������ް.U���P��[�!: �rbs
t�jo��5�@7��T�H�D���m*��4ʻ=��,a���T����y�o��J� �J7��/����i��}{�R-T��<f�n[�!������z��$A�}UgJ]M{A�9�H�	�Ǎ�w��i�2����%�ٝ��Gp(�"��o���O��(��r�VwF�;��؞��gp��+�6Ӎ1�	�8�P���zB�{Y��y.��)��������Ie&�����9�7!*o4o1��'��|"=P�j�/�l��#���^1���v|��7+y&$\=o'ct)d�+�����ݨV�Z�\�I޹�n�)�r@k�<��l|r6*��gD�#�u]��Us�$��Y
�G*[�FvL��v�н���C���M�����2�ck<�Fb��*��mEP^g0y�@�3ӷf��z	&t
I#NL�@2��.4�C*��|t�������&�U-�wn)�Թ�n��S�g���8�5�|89�l1խ@gY��wg5�"�^������)��TnJ���n�M�`�:P�Lv�<�,��л>�����p�B���LHX��!\��
c�/�_ȥ�R��}�[u���Q�]���H��2��u2�b���wR|sK�C�ꇐ H� �����E{�Q�3�rocl�g[���̽Ke��ٽ���0:�w�ؖ
Ӯ���(�U���{�Ւ9�Q�=�a��Z��P�q�%��Km���ʼ��CNY����M�)��7�2p�'�)�x~���U�7��6Ʊf��b$4��k��$.���N��H�}(���q�l�n�/��a�������r
��2�xg��ݮV��
���p�v���~z��ש��tC��y5��,��r0��&�7fu�d��	7�qsCm�#i:�t_�S���>dF%?o��+��	_��o	��S%U�&���	��ܔ����/�r�b��aH�˜��}JG5���ń}����P�z|^�(�캀���e��W��Ь�\3��R�#}ǷV��Ά�����dG�	#���E��sw(F�Z{��A������(I3g���l��,��B5V��3_|S����|'�nt0�5��>�Uaݟ��tw�]�2��XR���5J8:��~���\�a��8*�����'�T�����l�-���1��jp^�NJϜ��۰��Ă������\p�bA���V���aS�Y 7�p�b��_��~�y�4��*��R�z��n	y��@O��џ|z��b�l�xbs�9O03���;VC���b�:3I���wf)�p�:�8�)p�_ؿ
�\�l*��C�3E���^��+̯7�쒮�NYɻ7��W�B�pLw1UmR�y�VY�3��-[�^��*�2���t3|�Z�p���o�QB��x� !L
�\�� ���g��Z�h��(q�E�6J�K=�ެ �vl	�z]�U��,�g�D�7�i��|9� N��,E�P��6�}]tX��#G�Z���M��N�!t��D�1gvzw}��D�#3��O��p�[Q�b��N�J��g�_73_v;��eM�Á|$����`& D[F�GlJ1fi�8��G$ÔW�7���"����u����ɷ��. ?�fK7q$� !�jM�=C�e��+�t|����⤃�E����d������3։IĮ��3M{�<�E�k���Dxt��gC��;�W��p��f'/3x�F�<&ve��KV��6M�^s��w�t���ٳقh�t�T�f�>S�v�b��m��M�79�/,�s�J\It��T������0��MH�#�ۂx���I�#g��墢ʪ�(�@A�w-YQ��e<�sч/a�y���}*�o��M(ۊ�ġ�� .�)�_���;]Oߪ%��QS3�E�J>�E��=)d���X ���Z[�U��r<O�& �`�u4�Y��?��a�oRW��2�K����T���1��ج�7�v�숹_����"��wy�gG)���z��j��Llt]lA���}�����'���l��~���x�1��~��;MPY� G{����>�B���;��}����vB{*�8�b��2k�H
"�|(��29��s�����̮�5������MT�����f�8qG���L� �`������yAn[r���P'
v��OEcax���l�I�]��!�e+D��Z��ܗ�.���Ʃw_�&]T����G�'3pS��_~��zԕ�K�i�߯���yɚ����!��GOU�'���Y��<̳Z 3���3�N��1S�0�o*=y�V�L��o ����?�e������Ww���� *��y?M�&��K�Mq1��SA��y�w�Ҍ�6۪E{�5�����5��w[�������/���oyv�/� ����ٷ1���2sĳǡ7֨���b|�vG�ؤgd��Tq�ՅM������B�b7�ty4���>�F4���Ulc�K��Ĳ��'�O.���j��H�I��&,�8�p���F��tp}Y�$Vi�/ _��P���C��Q ǁU��OI�_�R�"�)�t�3�*��@4p�	�Yp��ɛh4��f|���x�
�k���=։��%�_�'�U�n���_��7ʃe�
����(��rx�8w��1��Jr0�#k����s��������q��Ayl��Vgc!2�|�6�U\���l�Dd>�(�|A^��ښD��7�2E�3����+ ��h�e�H"ЃV���.�;�r�:����nu�]��3i�����q�4z������V2?��LMD	� �}�&;�2��6���C���{T��C�k'��y0���L����g�L�L;�NR��5�83WR7��K��)�(���R��z���#o`)�@"���/���G�z;~���A���Bn��<���O��s(�D���cANE?��c޽ ��oq;�Ū���6��/X��#�Q��^.���J[�au5 I��&�C=}�M���1�AѠ}t��N~Pk�WׂǟtbG��FYdv��C���P�J�!�[u�q������+[�gbWT�{��Ԋ����S�i�k��� �G��Ķv&(��> =�Ǟ%&�S�r����}Ӻ�[?�Clk�$���~�g��ॊ�N�P�Ӕ������P��q(L��N���XԳ3(j�Ug��D��{�xWt��}e��Zu�Ԙ���~����`�����K�O'�=��*���l#��b ���b�HR6wƣ�<�0]��*�� |	���L�Ap���Q��oRk��R��3}u�e���Ȫ'�+�o&y���]�(de�o�/���9�dqGl����-Ӯ5�������!G25�S�Q�(eb#6�n(g�*ݶ<ʠ�l��@D�����S$�"k���׋v���U�Y���h�����ъ؀bP�B�b/a�JT})	�?�N��),(�4x��JC4�ZM���;5���W��4�7�t�)���}E-�6��1_�S��aM�Qd|�~׭6���*UV�Z��ߺ>�q��k�Tﴓ@��\ت�9��?E�]a]�x�ԋĥ~H$!��y�%^
��<^�c�`[�\��%���{DҐ�N򮈷*�Ï/��)各 K����,���*�ʧ��VA�L�{���0�#2vC|�*6	���a6�9d�Fk����1*�b�22��=&=��z^6��~x@+�t`�<��M��\�"Fa����u����T�(!��FL��ݟ�
��c�U1������X���}��^)ikTm��8j<hִ�4���C�K�Fj9�- �9n��Og$��G"b!!���a9�A`�s����b���Q���,Q�ϻzXci�|�-�W�U��:	�\�UY%9�7�T8׾��$�n?���S+�%��kO�+A�ݾ�{yz���H�+$�UZ�,�����u�U��#|z�4 �H�-�����v[fZ⳩�^����/�7Z�uV�g�a�.��֋�4���q���g��<84�����ͪ�X$�]<��-�����uC���f����%0*�� �I���Rw�B�DE���GO�Oj3y��_��Q�ySN��g�u�M�e)aN���C\��ڬ3�t|�&[��*���E샍Θ��%I��-a�,��p*���Ɠ�k`�`�'���J���0�P�4iMCxQ܁Vz��JB��|s�q�y/F�*�[{y��@�-������$}2�x�?�b&}��Y�h���R:u���mgUg��l9�g��k�` ���3�d$�^�/s',iW�DgD����0O���ˬx8�4��)�	�c��'å��3�Ӂ��tR����x7���t���� ��<�SLp�_��z��34��a�ľN8��~p�VȒ[�r��]�9e�UO��<a%�]k4��w�-�Vcq�-�?4�؈���I���}��a~��i�(Gb�b���n�V� o���e�jC�����(��;�f��QΗ	����Y�~xR��5�2~99�+���r��P��x-VFP�di�Uʜ�NX76�E�S�hf#/��9Z:3|Dx��:ܩ�84;9��Yl{Z�����7r�(�y�x<�]�������/��& �:��+����GAUh�՟�R�k3i&#�`�)���\`���-|'�}�ߛFI�<VN��Jaa�d�D1��W|.��-4<��ܥ�E�VU�T�.`3:D��ʂ���|VP�	�5��1M�KY��-g�{�@�O�k2��Z�B?��6�4�<Fۼr�"��m�7���	J�i�%���	꧅[1֏L �&��h��UȴJ�畯�F�<S��L$1�rN_D�S/�'�O�I&-sF����Mt��K�S�p���|0Zt��v}�QX��I���d�h����E���W_AzvT#rlG�몶��h�=�pok��Eú6���z`i�ԝ�4/"4��x��I�=\Sv�H}+Q���Bv���5��CM�6����-�hf�&�_�ՈBUe��㴣�\�D�,���|mR��T9�;9��,�J��jyw35o��L�X3!d�\
9�u5�6��z����_QzҨ����,�_@��8�ʪ^������b��i��kW������j匁s��0y�zbЀ�"���"�?~	9��^�������fKb�%�Bq��.�����8��y�y��Y�c0!��<_��B�/��R���]M��#t���B#x�
@>��Lm���cX��D��:#��Q�]�EB�;�d6?w����N
Gi<i�Q���u'�紲���q�:`����Pf��'����P�a�e�H�ꘖ�au^��,	�����R°����T��-�]���P	#���a^�[O1kCm:�r���	~AF"�ꮣ������FWsǗ���?� �1�~t�@,;��#��T��F��hd���DM �d��C�������>LEr������ƔE~�b���K�V`H����4����5����pQ׭�R��4�F���A%�a����;�(My�;�����B��'3��rtr#�gc�Y-aZOl�q��%ktrQ
�]6�4e��3�Pd�!p)��,���q�A[�<1��;���j�,f�y3(9��<��Q�&,Y?�/W�ή�6��Ӊ	MS�1���{����Q�	��e�Ej�1_�66d����H����:�t)�5�֔�W�T4���������ؑ�Ew�'�o��i0���f��i���!��ia��.�(��L���t�+Ҙ/[B�e�ױ���zz��'jZ�PAp�i_6\�ɛ���5����V�_KۘD�̻^ԏ���9#��S������=��K,�\��ȃ��(�2� �P�j|�0^-��+x�)���o=ph��u>u�Ҥ���x^i�v���wK�}G�B��kȎ��^Y�܅��K06,�A5a�$�����6�<�y�p_^���A_�N�8$Y�֥��-�g�����M�7�����M>�]����Z��E>x<�e�$�N�^v�ze��G�����,�Κ^�����*6V���ə�]�9��w��T[v[��S�%ZC0�@�ٳa'נs5H��%�ʞ�}�,��<a^rw����Z��q1��m�e�Y��kN�?`��2ſ�nnˢ.��y���ԧPsU%�#R|J2�0�%�#�ĭQ/�$d�~`�� �/P�b���5�B�Hɉ�6n�SX����)`�U�������$�-`^`k�;�R�}�`�+WkM�v�8���[�
ꃞ()vȥ�o��-��pX���l��kX��3�����x��n��I+C���H���qa����(RI�-����tt�ʋі�Z5L{�Z���}�m⬚o�n�c	w�;3Y�M+Rvsk;��	{0�T}g>�U���Wa^9��E�!�����E8��2��g�ph\�{�(xO�)�*A2]�iFPB�G��=��[�7bO|.4z��Xʹ�=�*�k=aש��Q&^Y@r�)`�����Χ�&�Q氊h7� i��������.W�O�?��jn��N�خU���ƾ��?��A�di�E`E*X\93�G�!�|�H��^�f�o!�J����'`;��R�W(��+�R����>��Gf>9喋�,��| iR\P�3�1������wg��/4"��Kf����]���%8���w*0�Mţ��Ƕ;�MD�x�J�ʾ�TNe��H*�i�:�Q'��W|8�k�c�"�C���d�a��E�7��HN؜-�k��A�m՟҃c��M��9���L�E�	["L��,�pԧ]\AsR49�^��l?�4h>����~��eK�:S�ዑ�J��٦d�-�ǘ-�(p���S�(S�r}K�,��.CD�sQ�����28�|���i#m��J]�/���q�O�=�zm�B�����@�2��O����*8i��R�Bcf
���˛�;���)ݱ��APz�o^ د��v��^���|I��Ԟ?�'B���Zy^��v�ݺ�C�����)�ڱۻ�`���WT��˵ۉ��y�.v���4�m�ݥ��O(%pP��o��϶�+6�H�YP��	w��(SF���9�2��nn�c�Z%�m�.x��#X�{��R�=J�?�f�"J��
!F��^�� ���c�`�$�ߺh*�ݭ�y^����J�g��m���̾P�z���אw���fe~̡������,�	����/@ƭm.���@X�z� �L�I������	�Z_�?q���zX���/���Q�Ҍ��0̾5t���sč�E�"V��pJ��i���ct�ah2+����l[�2�������$�m��b�f���O'nT��<����D'�-��j��c�#ƈ��7��F퇺Ѿ��.��}=@��1��7�O�_k��+�wcO�O�u� [���ȩ���Mq��I?	����&:�-�<�Y�]�ZN̯�|so��`�^���M*=��(4�D�8\+��@���_s�!��]B��+�Ċ?��2q~�ߦϜ]�"� �h�=��3��>�.��������[����L�h!U�҅���wJ��ik�'�� ��@����O*Ds��� x�,��.Sk�[�o(;{U��e ����-ny2�s6 _��}1�*+.��iG�X�l��~t��z0���-V(W}��Q�\���蛺���� ���8��zPro�U��I�`2S�~��h�(�����X���f�Tt���C<���E��2�{4൩Y��+�� /n��)�v�R�<Y��z.9ܠ�k��68}�֦Y�{�yEn;��]�/��_N[�
e|���XW+��Nc��J�*HPu���?�s����5Ϊ�@�����p�)ݓCP1��X:硈ozwfetĊ�aO���YH�D�q�õ��<4��Ĺ�0v]�ƍ���.'���C&��(%v)��ϞqV��2�z���y�}LFIQ�y��un=�V���1a�]ս�s8m�*2���-SGLx*��K8�ZŸ�q�ĵ�=��2��#����&Ke�!�"�[�3i�G�#r��#�Ԟ%�yY�u,���dk��O<f��M ���ݞ�8��M�u��~�8�)X��JN)SG�p���u1��� ���І��zILjuj �Y�lK�x���@�+ ̶��g�4���G�X�f�L�«�B��"�xi��Ԥ�k�x�2V}_$m� /��
�|㧃�B�g���}��1O�!IJ$q�R4O9�&_:Ma�g�R /�����~l��u��M��\��;�bD��k����p �&mm�%��X��p�A��"��=�4ojݨ6�Tx�b��#G?^�)@�}���nuR S�h�LT����s�..�)��Si@�M�+��cixH�rH�F'��u�w�r���;DG�F1��݅��8Ki�����o
�&g��fC�v@:QLr
Ğ�//��F�۸bj�@��4�ࠥ%����k�Ws ���`p������߶�$�' >E�g{�+ՎF�N��B�K�@�G���)��!�7k�ړtl8���]�j��	1���1}��Lɨw ������ӅH^M�s�y�b�e!�d�'��Q�"�}ܙ�&!����b�'T��6/0��F):?mq%�_X�ڜ�t�F~ ��j��tF�Ҏf<�D%&N`���q��Vَ��������ߔ�ͩ:k��ɺc�y�[,�CJD1[W?GH�CP{tL�hB�XH@��[�]G��K���6���ta)���=�Pg��ʐ����͆�m��ך��B1��t`�kD�ˏׄ�@4�ŋ�mp�oq^���%�v�*��~k�^��L)�������[P�,��H5>�Ҹ3��n�'��q��G���s����J�x�4�C�f�>Ԍ����Ta�[�K�kb>��U�Ek��T�~2�Xr����ME��QL�@e�!�������N�0��=`d<_�B�H�Ie�
�P)`�ٽ�O������H�%0��!�UM�,W���Qq��DE�~�m���'E����9���bj����e���,Z�]�&�e�>�5OXp��=[a��'�ky�/fK�r�  4�X�ݨ]@{}�wl���Ɖ=���/h;b�65uU�я	|Gc�Y�x�Y�Ct�\�;dL�����z;PK�a��G.ωx��8�MnSq.(�v��~�Cb����E|��4���P�=�;HKG�B@!N��߭y4���I�O��R{��ߞ��y��/��]ľ���ghm�&�<b�(�#��h�
�E7��Z]����/W�'B��R���\�P�ew�P��%�+sFkDޅ�ϯ�F{ޞJ, >O ��*Pk�;����o�Uѵow�*���"9hD�s�j<�?�-�@G�T�\�~2������pVD��qu�"74}T�δ���I6���^GW��-t{��:Hy�xm���ť0:6f�b�W�E"��/[VvU��A/�<�Y�g�[j-�/xIGK�ȄrU�S�)J��;Q8�p��C�b��d!+�Q�ф~y\FH����Z@���0�^@�����[
D�
ȧ_n2�ϵ��Z]���k?Py��9��g.��2Y��x{/@A�6b�74�T��Z�a��ie��ϷWb?��)/
D�!7��Brb���+���%�u�1I��s�j��d&g�ʖ%N(9��u��Uv����������]ya}�K�.{��"�@�.}%�gHX�c���(4< �&�������4抦���D��;��4��m�:�N+#�!��v��.�3��F�R�W{T�AG�	�������0����W$��~@cFEO!5��ZA�\k�3��:x"��p�\6ꝴM�-�1�����?V�5�E�<Ł�u�sW-:g���=� f�cƁ���H C0?W�3km>����QN ������[�յ��6��w�ϑ�-��O�Qg��#��=|$� B2Ҫ�[�r��.�#^
�U��吋�+PԸ��Aiv�7�Ϋ�EL��ǿ��\��2�P�Ew�(��˲���;a�]y ɒ�S5T��5�#��c�ДN�4�+����T'����Uj.Ϡ�,��ry�~�e�I:C�^I��g>�ϙI+�`�B�X��ّ�S� Z��*:E˦��V��6*�4�^��?v�ȋ
�27 ��7m �'f��~�����JťCœ�<CEj�狂-��	�6�E# �a��X<�aX�B|P[�D�lt����Dex% ����f~7~A.'�F����GZ!��VTA��e�o6�_��,�\'�#���u?�*�c�!	@�v��$��O�W��#H v�g1P�����)hY���)�kU!�J(���m�ܡ$�S}�c��s���yA�Ϸ(�^sdS��*q�;�����j�i�jt���D���u~�$�'-��'mZ�ܱ�z�0,N+��%��8#^�q��5y�R�f�E��I���C�?i�E��J58ԉc��-��b�b�\j��[�
�����>�ekI�G�!t�6(��υ�})�H��hD���`�"E�ָd��5۔�ö��Q�F��?���᠑p����E�p����I=V�:��!�,���6OA��:Zw�j��� �'n������Ҹ��"Z��t��q��I~cRyW�0���y�㠚���>��J��g�V��S_��K�T��?��MZd����8�C���z<Ze�� �
v���t/���JLDf5t��Zl�.�'r$�7��U/]�'�����#�'	�O9Ԙ*,�~ĿY��n!��^�� k�J����t窄�T�ȱl(u��I��D*"������� r@̤���p��p�g7b�N6�QM'�8@��Gl��m\:	����Y��lrR�_��cR��sC��]P1p��xdg��Ξ=����p�$+$�<p��/����lF��"ᡋE�}�d���"h�M�	�)�@������������h\�B`�;�?Ѧ1�Bۘk_�vW���q���]���� ���h��R	<�B]��������vi8�J+��[��6�>�V�y���If�q���S���׺��*X}@	��� �4 �~�zd��k���+�y�.���6�f=rذ�(LʜG����uٰ�v</��y'#ҎU��+^{���/�P^e�.!�k��o�������c�"�g�6��x?����bM�uFL�ִ�DG�� PO��B2�������՜w��#mݛya.��`D��'�*���B �\ �Ea�[SF��ۭ��K8&���*1R'3�^#�Ap��v�?v0N
��vh2؇��8��9��_�ϭ��ɦl���>Z���I�%lJ��aVk|�_*Z_�w�EZ��P�Gu�ÿ�N1_{N���"����L�q�D���%�����`Y���]���b�qG#9���y��r
#@!#��ɮC�E��k�W�Z�X��S�bq���5%�'W���m��C�7�uL2���ے<�~�첎ܔޯ�\�0�+�9O�>��)B��+Zo鎥:)*�ɾ���;
��?���ص��W{د�����z�Ʒ��HI1��òy]�G�Ņt��8�gqs��c�Vz��w��Lb���V�Cws���smÍv�S�̘��� ڧ�Byz��!0�U3�)�ؕh�@�ׇ-�������,�����*��o/�"ɍ洠�����;�W�g�n�z L*�|a4}%���	� ��G�Fp�q7�C!E��=�b�b���1�}T?�٭3<�K��@v]��5dm�d�K�*�´W �k�Z��V�Q5�#���M��$�A��#�[��B�C�K�%�d�d҅d�T*��-�VH.��.U;CX��������AO��'��f�����EV�G��I�p�s���0���D�p���{s��Pnf�L����*yraz�|Ʉ�x.mk$���GƞBb����\�3�x���)��U�xzG�X:I����(���]��k�O�bn�cn�v��,�۹I�)��F�ܻ]������9�x��(څY(2/��^�q��i�F��,(~ńG�ͮ5�	)�����G1U�6(t|��RHb�L'���7��4$~Y�k	���M㭃�̜~ne)q�e�3GN+��0 G]�V�tV8�B=swwQ�u�
�4/�
�36مO��%����;������x%{��E=H���7+�lX�9)���i�ȗQ��\J�eP#㷔���	W���*��d�zq"��w� ����0�'SA�[��1��ǅt²���XƮX�U�aL}���'�:��� �HB��P9�1�2[���b�u��β�����_�hA98u�K����Lj1����N�e�|�&Z���Ǩ�`��7{4���DB�b�Fne��٪��r�[j�7�mۢ�xS&25YP��83���kɷ�5�z����u
<�g��tt=��,�ӯ
	�V��n_ MS�	\�9���;�kb�Iy�+3��7���+8��R��fC��B�K��nY�4�&
;�>�ד!X�#��������]����o���YLߒ��Y��%͏�WPd3�m�3��^�SAK���6��r)ɝ|�t%|���0�{3�j3sY0P���i���q�r.P����7��ya�^�#R)r�gDZ��6��:e��c����U]s�|�q%��#�&�o����T��
J�?�T�������Q)Y��k���o�:p���jx�� n��q8��B+'QJYp�7�0Zx���G���?���6�*�Xΰ�%}T����R�gy	���e��Ȱg04��E�jH�}���+f��u ��I�=;� ]��9ۘ�r��=&�����#0tܠ�>E��u���a��c�Y~�CymSN�Q"����K(�Sc�v/����-=#e~�R+u���K�Gݭ��G/�7����&u&�t1�V����*��"�l��h��}4�'I6��
�
��flq­\�
Q��3a��I��4�����_��>Ɯ�F�>lBôy�������>6�쟖�;*;�F�P:{��V����ļ��%�Wv��	�:K4fb:�S�>:듁לT��h�Di`�KhD K�cF��~��:��h���.C�{8��$Vͪ*D?��ʑ�فE�.�-ጼ����L���j��w��k��s�&�:�H�ʟ���U��rw�)��������M�S.�qj���Q��`�ۭZ%R#e5���V�v�yѐ��T��m`2��}��R���:($8�>. R�	��*� S�^�%�)�B����vܲ�^w:1�������}�	����f����;�*�)���:��Ȕ�����mC�N��[�x���e`b�'3�3�V�8Ү��-��A���q2�.��FA˅��j�EEp$e1)��}�&����-u�� P�bo�9�-^����_�pL?V[c�g�Hz��J߸;Mp&��"��p6�`���=�6 