��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#���������l��U�~�׏O����j9�PY���`T���x���s����uí������P��"��b%>�1eτy�<�gܰ�N�Y�	� {��I�ɍL�ݫ�G�R�k��Q�!E	�5E��.��:�͂2��y�m�-�.E��i�����YS�
��@�H�ۼ��nD��Y�l"BU�.TԊ�=�-�����q���Ǹ��j��ԋ����tr�a�ٵ�]�b	��%�ɔe�)rYOjX5;V��R�������M\�	D��ҏ����9c=�Vͼu��Ro�P�Jf�tRvsY��c�"n�XO��	3g���Q���^�Bʹ�7gQ+Г���$�-��t�8�����A���<����l-��*�|d�n�~��ʙ��z�A��L`�5RT�	}qC������ލL�82h�7�v\���ۺߔHs�sc���R
����K�\�}C��k����5ϩ�� ��k���|�/��*T
���
5�U��䤲�@urQ���V!�+�1Ee<���H M��[�]�x5~}����/�n�=�v"�Eb5y��JM�n�&X�'_��m�*jC�F53V$.��vm�o7Wf^I]����J��xR����2\�8��p�uz����Q�E�W$B�X=�>O���FI|d��/�6���&q�x��2�+1�8�e�m����Ut�6����Uv�*�A�yAǺ�������Ŭ�n��� ��o�6�/��������U���S΀-w쾫�-2�u�Xo��C�[ ���i��ɖՉ�
�U;�!���*(��W\eL��Fώdc$Y<S�,e:�'�
i�F�a,���cݚ@U�{<Σ0���yK�������
cM����R;�ܮ(f6Ln�Cb������-����P��2��P�%J��*-թ)1{�/�#h�ֿ�0��:��p��vu/� ��U'��0u�v��5���K��zZ�s�L�p�i�n�Z������YV����j�я#�.K�U}����Ӱ�!z8��[���O�d�S�p�W��l��(��ɱAZ#��U��"��Wu.s��< �����FAP����t�f2�z2�CUm���yS˙�a���k�k����z-
rS�<���I��T�' *�~)����v����/qf�UX�+S�%��������3m
fm�5S3�ѱ����}n���X��k�t3�����X7K��]J�WV����zԵ�-S����'g�,�C��b}��kC�geNp ��0E���㖆׾��A�&��	��SN����@d�9$
SF�j�&T؊=��@��Ϊc�z{>����mÁji.	��	d�2�l6�!����};~l6�������gW�_�f{�uA�!�J�LҤ>R�0����_� �ꑨԩ��8��6'jjd�6�N��&��W��:�I�h٪��F
W�I��WN8�c���&�K1�D�_^�닞�
4�Q���N�YgHX/�=��9��ؼ��w�-�FL_ҋQ��>�VSo&�Wz)���b7�����۽C��:Ǡ�$��� ~Ry��a��8�+�����r��,��cl����ۜ���e�/�e��+g-�x&&�9A+�J̞w���`����@f�q�k* �K_s=�J�~��#8(�X�8=��H���Ƹ���G����c��6t�RE�L4���NB_"��$\:P �E!.�U2�A댃����f0v\x�2a��y��
`0E!���t�wVk6�=�G�AD�1q9����p�v0�R�K󔪶h�s����0o��Q�@q ��)e���W��ͱq7C��g<���Y�Ý�O�~�	'��8eV��;��d�^�f���F�C��J��]��)���Ć� v��ɸ!��n;0����u٦�e�����+�"ԁ _
fA���t���פ㲎��PG�h�RI<t������2�N��s�`�2,�74j1�>~")[���Vq���Vة�M��p��S>���{]�7�S>��BB��KUF���#�w$�Z�w�����{�o��חS�[J�N<���$>�2d�i�D�?bȄϸ1w
����.�R|�ҽ��N��͇L	�E�n�Ǫ/���)��3�#Kk3����֭�|��h5g�e�+␈�f��
 �^�(�6�$BK)�t	͙��5קx�8K���Ё@S��h���C��/69����$k/b�v�Q���<�^(~hB���� 2\� Ǉ��3!c/ٹ5 :�}�B�,_���λ�[�#Hs��e��3�4(&��P�i�h�3?��WD�{�4��)�H�"&����c^�l����ܖ/oI-���f����|j�Q�2���#<��N(��Q��7(��	Dr�O�ȯ�G�a1���hu_�!>�Aj$(k�3�+A�f���6\~Lo�t�L�g���N8Dթণ��`]�{"q�?Q�'\\@�y��gTN��C���8	��Z;�Im�3i�����i��A�D?�XY�������w�Ĺ�Fa�*2䥿�\���:�׺�z���דV�	S΋�(��y�$����1y2t� %�&g�����v�^��U��)t\�p��>A�����&���%�(2K&�Չ^�V��:+��9���j�_������+�@<��~���ǆh��-�J�	wFN�	��W?+�߶��~��~֪�R�k(MY�Ӄ�}����̡nG���y���!39��VϹ:ơ@^m���
+D�wݗ�kk�ωP/w~���eB����<X�WbTV�����#�4 �s�[���������F3^4�NA��v�N���j�e���<W>H��o�9��^�M�ذI��s��=�#؟ף/��lG���}��C`�׏�gJ�bu��P��7��(T�q���k��Wڭʘ���h`���S^���0��=���?��"U��2]��S[���9-����l��@��~Q�Fڲk-���;�5w`9��d�O����M�v�c�xJ�Z�?�E�n��DN���zŝ[�1y�Ⱦ"��2���������[tV0 ��A�ֿ8��y�
U�� �z�Tvlp��*���#k�.~��(棕����8��'a�8XЂt$�B:|����`��(���]���@1���kd����L?�����jOX��;�n�~MM��䄧|�'	9�8+�0��@�˺t\ mȎd��HLF"��Y��4�~3	
-
��r�v�r���I��E���������l{b���N�b$6��
m�֬o2V\Oj)M1�~�p�?��%�v5�{Cq^0��玑�]�D}�xq8mA#������I�UD͆�Ϥ���-
�ȕ���9S�s���/O�T���?���m�Q��Gm��� 5���?��r���\�1�evx��z��?m�p�k�
����T����H@k��n'&��x9�������2U��[����<�1Ex�Sg��Y�W�5�+���M-�~��"�iA�!F-�~pxB�#E�~�t����O��8��wݴ��-'�[�-���d� %u1��o�f�Ԯ�=A���� Er�#���c���r/b��*� ��!.���[�;�'}�ڠ
,> ��Q�Хw}t"9C�-]�5�J�0��t���Q�c
�Z��Cz��c�gnf��� ��*)�qf��6l���
�]�ݩ���K�4��% ��Ye�x�膗I��1��B��jk/���rrD�fy��������x�-^y�m����z�Ǜ�@�h�������[��3�:�~?���0�Ѵy�7en%\�uk�'э0-��-�R(��H	rE��7�]�g�:�M� S�Fū����/X�׽r��c\���d�˺klM��b�4j��˝p�1���<�~\��.�A��3^-�����FIn�5���r�*���{XΏ����{� �
������~���Y���Ћ�2?��S�A�_b�m�"<�"Z)�O�'��5�n`'~�v���i����c4maFB���wj�V�{-��G�K�d�lh�(�����4���e}{c�q��llN��ڭ��ˀ�(X�s�%�<Ca�z@6S��[>�`y���v���g�aLvn�F_Jt�D|�!`2g�{G��f����<G����~oW^�2�m�'9��S�6F��/sѽ~�ٷ
��ߞ�#��[K�Zm�Ě��䀇���>�S�ϙ��A{�|���!��3g�5��4��P��c��k���jyڥɒ�k���p���ftyG�����_��
Qz��')"N`-G�T�?���6>�mZ5S,j刱�Nb�zs8��F������~}��bCG >N�0=�m  �!�9��%�ڲ=���"��)aa�%�TN�Z�5�Ke�l���f��<ώ}t�����jj�;r�wy5W+�C�֙�8Z9�������r�D�����An�#����
���'<AW�6���A	��NH܊1�S�c})�����$��[��W#,H�5N ÈNgt*���s����֎ީE6�ѱ�E*	����_D�ș|���R~º#�z���j��$��"��~���П��w����7������N�j�;�-��)Y+p��G�K����'n�����e�6���g��?��^~��:�`?[&�c:`�b�\��&����#��9���b�.qd�+l0�N�f�b�O�ȝ�)h���6[�~I9��A�� U�Ӛ����ȔȘFˀ]ҭ�.�Q���\�D
K�B�x�.D��*�
XLu]��\R5q�	��]��<0X:�M��ҝ�P�*���J5���E;x6�3�3E���Jw�d��Vs�6.zկ'Jl�D�خR&�����o���Ԝq���@��f+���'U��p�ĒmM1����!�t���X��(0�(y\��`5��}Px�ILPZD�1��>j���N��_�ڮq�h��Ѯ~sօeE�;���OM�֡3(c�MN1|��g,\��?RC�����.���d�2AbuZ������Jt��鲆�T����i��!��ÕG������;FD-�2��BF�����u�I�Oć�$��L[�|�7.mc�W؄3����'� {�WA�Us�Md�u(�T�=��,N��ǖF�S�un�r��>>Wٕ|�4�!f�(�a��cZK޵Ui6*sM������m��v��$Jy���R4(p�l]6Ә�yf�Ѹr�l�S� �B-˩��4ELt��PH����xRk&����:� ��X�PK�bH��P޴����
��:g��(��78;���\nT*(�G�t`C�<T��$�k[����:]��V��
r��Vi�!�����9���!hj�'�3��޺R��������mL���꩒»���'S�Q�� ,~�w#a����l+���7*L�"Q2�<���]����^�h�$£ �8�|�EIlDI�% 	�����$y��Y����W�U��; ����9�\���
N���������YDߠت�G����s���>#��,�?_��I~���\c�TeN�Zg���8�-�����p�� ��t�8��J=sͻ������df��ؑ�/6���	�����[���g �퉹�����	U�x�!�f��0���D�[����*�u����G�2��%a2M�K_WҦU��<M�cw.�#����gb1������޶9���1�4ךƺ�K�̗�G����ú̍l��A��H(F�#�4'L4s����Lە�p.�N����g��\���S%��:?�U�U�:R�L���cPF�qY�t��Y����ƊZiH,��y�~��Q�ԡ�N���U�
(
c�sˁ�z��u�X�h@u?<;�4���呓�Efz{i:���nE�4�1�d\�8+a����~1��n7�?��[tm�h��O,��,w;Q4J�r��t�LD�D��L�!�.H�+��t/��t�bU#r��d	�r*��;�l�iU���3���h�4���o���H�T;�Ե�8�=��O"PC�?h�t�D����c0,���#�gh�2U'�U>�k�a��%f��U䙗�թL)�a��[�oũ���zB}S9x�(�-Y�&�`a�ك�[�B���O=>�q³�p��S}x����1�#F"�m@�Gx�����w���b_����r&n���Ƒ�"-�pjLw}J
2�g|�gUT�L�3��^�y\�Up����-������,X�1eL�E��������_��!��������z�����cS����[��d&�z
��k�Ц�&���������6G������k<���:�p|���
8ms�"n#��u}X��m��;���g�E�Vi��Sa���K�����+3�)��Oa�0�5E-��	��5`�����4�0h!��'T/ʖ���ǖ,1'DԜaKG�V���t�H����N�V��s�G������b�2��o�Ŵ�O�Xm5��r�����F91z�OL��������m�������U����@� ��9 �`�����ϣ������6P��s�`�㐵���&Z3� �ȍ�Տ�b_p��F�����˪UhK�yH��Q�F�[[��U��41�s(���Y��n�x���<�:~��� QA���O��>
�c��F�t�D�8#�����:	�8ۗ
�Y��5��7+�RK�%U毄"C
�b�%��8�.eQs�P4ΐ�S;f��E��cvHB��&��M�ť_�/�>�n�|��<�Ja�)F�&ֆ�C�az$���&%m��}eN?�d�v�j��Z�&Α���ԬF+R��p�-, �P9�_&H�	Fë���Ղ�G� ��%"��	��v�ݼO������=�	|��7Cp�.�/��
�`��,9��=�eG0f�=8�v�3�r�PtDݬD���12H/d��V#%A��b��d��in�YUʫ��ӵ�n}����th|0�Q�/��O���3/B	;�]{�\���ȣ��,uloi`^>
�yi���L����^�LC�63X�<�"���sg=��!�O�RG�<�@��q���Ѫ��H�������U�H�e	+W���� q��Q��k.���G�U����Ї�Jr{�C.毣WM��d��ݯp��nh�%4�Z��w����e�ܬ����%���_�z^h�����`[�P�k��UT<��c�����ޭ�����f��9�C��Nz����C��A^/V1�d���1��,��o ��?r4f�.}��HWv�R.is,X�އ4��N�
+�w:n$bYus��|�+��� �b,bV����w}~c	�M:�Bd��ǐ?"�:�km�ʭ�Y]�}��YT�G���F��k�n4�A�MJ��%x����}�؊^+�)�+G�^c�%�%�ަ�d���mNt3��I4�x�-I�M�u�I�]	�Q��"� ���A�9��	�/N��!u���ɦi�[�I��9��R��r�0_�J��LW����J�5�#���_[���Q0�!��h�U�->P�kE�C	�SPP�W,߰�x#u�YueH�
��T��%���D�1ȶZQ��q��S�#�� :n��8�
!����"?�`^�g�J�h{�EJ��&��P|o��=k�ʧ³�w���VP@*�*���\B��s��1�Аc@�cL`�?�:ߟ4m� ��F	��.���DE�����soi ��t�K�!4%g/.�����p�XO�HRj������8�e�>L�̴��/}�]r��6����>�nwߠ���R��Hv�k��*+~���&0�)`y��g�����tp�M���4���V�(����4�^�E��/�����6��
GWl���y���Ae�<�zbpQ�%�I<���1��h4
2y�����J��48dh�)^��Mt
Zdoa�[[�;���aqP�� ;����_`�2�6�B��4M��7iRT�t5�%��Yvr�Xw�j�a�F4���
cQΘ�M"d uc�P����+j$2w:�(]�����?$�Z�.L.1�A9���+Q´q�#�_�-��5�۴��Ij�QQ���5�	;�6�.Ʉm�4��s��*�o�E���
典e�
�/D.�� �AzȪ�HꋋL6|p��ތ��l��\��H��,? �
�̟փ$%�)Ф!����:j�,��������r�t�4�;�Q��}9�j��i�8v[�`�4@�T�URU1(^֭�aM[H]�d���m�c6A����q���>�elŧv����#�Pө���9�g)��$��lp��GW�ۉѣ��Ĩ�WB�=����\m�1���e���.ޔ���Lj�wUrSt��rbj�]�TB���QƵ5�)�@?ȽK�4�D��WY��؊H=�51��s 8���\&s��/3��Ó��4IRV�j�;���+��}�A�2��:��gs��=�����c���0z�4��ć�Uh�0/�.��PN��FmD2�|�� }w:�<�n�����9�k�"���T��w��\OGK�O�a� S��9��T8�e��N�R����&d&*+��5�e��p���)y�V��$�1���#'M$���;S���b��?�ojT��C��n��DI�6�|9�=;_�5i�۝^���?z�\���#��+_Y�!��; O2A`굓�3d�	dc?W��-�H$�p)H�����:z-�:6��.m ųG�^^��g�$�A��>�W��ܚ��%5Z�
�(�Ī4���b៎�J��N[B�@�.� �MT�
}�N���y{�i 9��7�v-h�������������-&�_z�Yw��bE��FlU��c��?�Uy���q����S9���qŝ�g�Ғ#OM���f<�_5�ljn�樇�}���"��sKI���>X_Q9%Lڷ�����W�]���J#ܡY^�V����h"W��]gG)��r�G���2�ݚ+�ȲhDW���;ڣ��2�vv#�UEv��)�[�4 �>^j���*�1�m��~�c��[{�G?����QJ/d��pB\W���o\����f5{/��nڹ�n�.��کc�+�n�h+�Xf�`�L ��t�~���6L�"z�%��;!�����۰E��wH�
88��THځC����p� �c��K�>��`z�$�uG��C�%��R���<xG���H5,�P^`���G";u���L�_������גc��iZ�,�ᠹth� @�4:��J;>#pj�"���O�<*�R��u�gM�ʾeM��r�)'9 �.��)$/��e�KM��P!2v��7�������;���Wu�ŶB,�w�%rP��
B�l����"(.n���*-�4j���S�Bi,��]Q򎼶,�p�Ѿ�m���RG�t���=c�fWZ|/}��qn]��'t��Q��.f�c���2vj��M�;�E�2�k�X���Ǚ�2#�i^�!�鏁W�?:�l�<���8�Et��^#��n���1[��4E]�|s�H!���\��*�y��V:&]������e��f�#�C,`
ǔ�:���i)W��tu�a&-��JM��R5�6�zڙˠ�G��V|M;L9+̳"'����4�cFԵ��<4�Fcp�P�w�W(%��: ��V=ړH{���_��0���DL���2�a�d-���^L�9#z7V�Cf��J��]�
-�_�A��6�7��Ѓܚ+��ch�^�|z��s��N�c��vø���/ѧ��u|og7���8�[���N2BOf�`#�0�ڑ�E��*h�¶�*�/M3��g��h6�U&���ԅ��t���C(A�$yc*�l�����i2 ��tz�YMs��?��;����`/��4�������&��e'K���6���.���ͨ`!����l�
��Ӭi�ơ���r����늯��,�%ں�{��T9�bA���B������fx�<n!��#Ӱ��4��p�z-�,�U�K�Щ�e˙���D�\��<N�b>��A�p-�B���E�io��O�ӅD8c��P�L�B6N��kzе�J;PXʐ�Д���7��e���w���Е4g�z�W;&�ʓ�vZ%c��=�����m|�a�g�4]����q��	!۷����dx�gjs���3os�ɱ���l�T~*Yt��Vts�+����;�M�w���ݱ�U�έ���v��	t�������l��X��a�߻����ߩor1������>��RexڌI%YC�ڃް�)�Lٗ��V0�\!XGvUr&5��_�ﬓ�MC0k:e��?�RDg���.��f�8��� �3FFy�Q:G�~�����f����"�H-�3�8�g�_gTUM�YV��ɩ >ڕ�fn%w8a�t'����0o�3�@M�ځ��{d������c{�H��?:«����
�N���Y�>�fYT�=�n�4##�M�l#��9�z��+s��|����0�]�����i�{�����2��t)t�J�}կ;�7�ۏ�h��n���[p�Ζ����X�%�n�7���w!���٠�OJ����QLGD��!(/��U#c#�Â���h8�@P0�Ɏ�4�G�{���Vކ�O��:��4��c�7���=��է��x�Dl8��q������m�(��2��r���e�}OQ���z������Ka�h}Ѵ�DRpr�g�)���2�;.^��S�&@��Aɂf3�G9�bܤ$x�L�p��c�2���p��/���,��A9�D�VD�c#���p�>&�i��hq��rp��[b,}9�wc�6�R!����So�($e�LrQqɢ�h$v����ٸ��b�� ���[���յ�����"U�KQS�]����sW��+��(>jc���S��SX�����B�<&AѮ5b0�4�
�x1�Y���(	�D�ߵ�2&��O�H/�ܟ=X釵�l��,��v�|�R�&��OW+�I���*,�>q��9-���a��`���^�6V�`4��jz�1�	 4�/�y񵧗ZP���#��Jt}D�]�S:Z�Dئ�"	X
��AW�}�=&J <|�����c$�U*%��ip���
�!�Q����h7��*��Ƭ�.re_��d־��o9���Z�i{n�s��"е��7�Od���z����dx���&qL5�	sA�(�5>�i2��k�p+����m��)�"V�,�]���ef�m����I�3�r�b��q��C�����$~\��l6�,suI[2�*�#`��t��'1'�N#�(��A�
;�0h>m�6�܉?��jծ�4$�ݾ��'�v���YyJ���O�`	��Tf��fr�����s`�u^G�C�4B��z��HU�����t2��]�Y΃p+�T込�@����Mb~����	/�ϟ���eT�� �s�gq�r��WA��v,F戍�����mԖd�'�}�tt.�L�*z*iyW��W&�N^���M��w��tVN�1��XJǚYȨ�{�xȃF��:n����a�w`JNa�)k<o�!5�L�"���.�Y�U����~1~f�|�u�ͱ�(C��Z�v���n�l�٧T<rg��3����L�� 2��h�W�E�f�:�6��P��b2�wn0�OL�B,���ÖW9�`�>����u����;N�i��	�c3o����x�f�
E���̬��)C�)o����Knq<�G�d��&���fQ�k�R:Rc��e!iC%�VAќ�P�F�`�j���/L��{/���3��v��TH(�r+��{��Rmf8�/���&c1@Z-?�v���=#J�
���C�-��j��z�|#Tl�iR���u�Q����9!+�7���N&�m9g�t �ˊ��t�Iu�+�HL����~m��v�gMB�R���f�X�M�M8� dA=s���M�˿~?.�T�k�8k�H�ױ.̇�6���9��`hO�';��I����zAŘ�Ϗ/�0[M�x̀~�O�(9�y[�	�N��x������:�
u������_R.������7�%ـ�f䁆E�Mo�i�������z��ֶ1���e%��z�r��� �"��`n�P���/�J�r\į�o��t�ؾ��n�[��(?TM�,�� ����|�s):߾��P��(������/��x3���5����"�΂���YQK��)!�ǵ�A����}%��s{Q5J���Y��
;�L�r�,ދy��a�5q�7n����'g�_���g9�����9hn^lm&�d��,&t���%O�KN�a��L:�#"�J?�,/��g�>g*���9y���t9���nY�咉2��/���	��7�3뢋# UDSC��Ykos��?����^�&�����s��fξ}Џ�b8X~�È"0�ke��O��臓���
���R��~�#4}FE��n#���L�(�L���&t��Uܶ!ro�
���P�{[(),�:����o������F^Ѻ�`(����.s]ή��vA��<��)�&��U�Cք����Z�	�U��ۀþUW�F���z�"zL� ��J*�`>���˅M�n�!�`�Nv��'��$�푬��7���&��p��u0 ����/p�������(���E}ì���l�L=t2U�9��G�ŒF,.z�JN*sl���玲9� �i��7y�����<Q�:j`��vԝ���f0"������.nS�\Kb2xo���f��ԡ��l�O�:��5jdN%`��Y�M�XA�O��gP������ �'nz��������hs6ĆqtAe8XyI�c��h	�y[�t���ņ�[4��0��j�,w�:~wΘ	:0*�נC��G�# ے��� T�8�_4��ݧv��.��k_r'�p3���Sm��b��"|;3h G{l�W�V�ʿ�|��W �W�L��Ģ��y��G��ve�_.di�l�ױH/��*�.�S�����vd��3�G��~[�Ê���i���h
,	�����x��%�����#����%�ő��ѕW�nl~r�����7�!	�KR��W��d���ǰ���G�y��;�a�?U �Y_\���y�s�
<�r]���	��L�|GV{Mq{Td76����Ww>o���7�a�cq}���O^����45Z =�M��𦸹����Y߅�\�F�/����j�*?����ߌ]��=8��>�7� �Qcfz�*������' ��e����[q�h�����:��(vp���a����ͱ���=��\�N@aa�=��vw,^=�ݠ���0�q�Rǥ�U����CV����+�|����2]Tt�j�O�
����"}�J���v�D@ټ|ie��������!�ck�U����"����^E���7;������������2L��`lh(��dK% �k�]w�f��b �l�%���q��(��<�-�BT��=�Í/���}
ȝ,�K��'n��'��؋o(��U���֋���E�k�4@ N���}�Հ����l���X6��v�K�}�����/��Sӱ�
��E5U�"�>��M�~�K�DpN����� 8V��$r����+��S�f�@ݘ�~�4�qp���&�)�(uz��/���J16��� �t
�������@�;5�˻����dM�kj�"��HV���.�Z.�-��)�i��(g�'^�tπ��6ʋk�2���~]`-������ �en�_�z/1��\���I7��b��%� [k��~P+X)|hӠ��T�ޕ�^}���
:�ˆ��^9d�|J�#�.g)�$�W�u���E{>q2�/����)��N��~e�Fd��iZGDO���ד���T�uMR��Q��No,k����ւ�pE�*&9� $��*� ��F�IH��p�����f:�H!q��sN����!�y��/<��)�4SƧ��Y����6h2#���J�V�hr!�ȋ��#	~�w(�0
\� u������2gġ��CM�!,���_�)n{�O���j!�V��w���A��5S$�m3�ǎ�2��F���K�z^��ҁ��#z�^٧�A!����^���	��"⻨�Lz��N��00TPеw �C�;2�'��R�)�sȈ�Um����<*ȖQ�TM4�iu�F)X<�G�|Qre��l�7Io"��lm�]�i�+Q�����cE�V�^ξE^L�(\Mh�;��3��V��]������g�n�z�O�hGKN$q���$z-(�_�N֣���4��Q��\��4�+R��s�����~���ߥ=���ٔ�
{�?�P�_�l z��Z4#���݌����e�Û�g»$�N^�
�P��!��F� �]���)(Դ�n�˞Q�>M!� ���<��ǆd:)�����g�؆�K[A)�j��:p|�ѕQ�N�_�kJq��}��#�"��ٯ��� c�8�Q����(��[���{��]�ʹRT�8Z�V�D�W[��d�;B�&��g���Q�e`4V�)�ͽo�,C���9L������T��Oc_��k�,�
5�`h�������:�D�M�$���^H�N�1��"GC~���hY8����z��1�%H�Ai�PL�/O5����g�Vj���5t�2Y��`�����8d�4��X��4WX�\LO��{XSJ�ze@�Y��T��Z����;��6ֺ�{0���p	���[/Z�N���ڒ�%[����r��P���(������H<��c�E!T�Hޢ��c��A�8���|y}����/9�5���Rt�̀+J��N�����.	�'�u�(>����T,����t���ӆY�����^��cJK���Q��F�	2_/�U��Cd�K�[�1�
�����M9�1�3�����/x[^A��(���Y� �e��3ބ&*�Y�������1K��L-�ow��`x!_�w~���~(��t���\���F�_�Q-�˪B�Nmz+�K���F�OS���m@la=�}\̲�]���yN��v�q�}
����`��r9�+����I�N����u"'�FGt�\y�̘�q��C�!�T*#�d��ww�9+~�
�%�@,\�
/�cb�M�q_8G&��R���cr���8i ���i`���;�gv{b[�<�������$���2�.���v0��t��Ш+��$i�qiY�� �aΆ�˫�|l��G��a�Y�I		��Y.���Ը���rsY}��$i�ta��t� 0�Agp�����DA#d��ZS*x+:Ͻ��N�eX�QEU���]F~�ٲW�b���>X�9��Maաͱ�-�c'���(�����?�X
�w!��~�LGD�0��Q^���|"��e������q�鵟���_��,å+u�����N�-����LP�(���� gl	�ŜY邈<8��CjuvM�O� ~T�Sv�ݪ��R$&�}��۲gLl�1��%�虽	U�j�>�\�m�Y�t`�)��FX�EZ;w3�Ӄ?�1>AD��Vg~������6#�P��W��_-!�n�1��m߸w
rG��G^d��?0�V|����w�G-�{�߽U�#��Ns{1~��r��B/���2�W��7	F�I��+D����e��-�b����Ȑ���]'Ęޤl'/��2��a'��_�yZ�m:�3�V9TL�����m*}-Mpཫqz3E��W.������M�ELBš- x+q4+�AaM���+�L��>�<�s:�'�A$ Dle7�0�����,[���c��-(�DJ��&R�MZ���G�&�W$�N�J��|P��(qrԗ�)/��f���O|:ȳ�Nz�
^B`1���%��k�rǝGe�b>���������v����c����gb�i�G\�G(/����K�5;����]j8qi̡uTt �41�(���C]5�D��G���>��µ>�6�/�,�p��M�H�7��X���8:�6�w|��w�n�;����f�����FV���_��X�#�[�W�"C="Ba���"9a��fQ'�<�^�/��'ֹPN�OxQ�u$(̙^ޡ|֮����r
��t*� �_1�n�t9�:z����1K�D�T�p�Ť��KcL���M��VPګ�Y4���[���h�,��@ڃp���ALTi��RW�m�#Ek��P��38+34�X����
u��ݵƨ����b��+���]a'v�D��+M�^ �:��ؽ^~��&�X�_P$�%�L}��לH��������7���i�PpB�S��R�'~�$�=sn9fFі�j �v�����OKIcJ��bz�Eo,��]�?�JL�^��>�=����k��c��3�q�+�63�0}(��2�u"�wN�(P)�����d�E<C��M���/̯���c;qTŚ~�7�*u����hC�汀LV�N�ж������n�kڐ����5�5q �G�/j�6�v]���0�����)�Ϲ��˵��ݲ�m�Ny�'�*1�a<�p ��m���(#���#�q�9❠K�́"���#�Ŏ�x�3{i���ۦ��fM��N�+}2���{�ہ-f���x�:�7�-�vt��i���B C~أ����\4��� u��y�MUs_!a�[U���b��i�h��
5vH���S*h�P|�e�]b�Jk��zQG���@���n:�[D�F�'���wZ`���-Ym�9a��+ф���� ��RB۟�Z])u�҂rN/i����C'�BO߉�Jw{-F�ʛx�!�s�!���f��� nҘ�74L����o0��k�;�
 �A�:4���s?b� 4;�`�tq�i۽)i�̛���Ț�*��*�/�	(<�:��N��x���U%�����=��jS�P�_���]�0�髞�B�����ʻ�Q�FN SsG,x��%CWB��H��Y��>��]�l��9ϥ0�vkC�������j��Rc>�Dۋs-U�Vu��"#t4���1��?:�a�9-�.� f��o ��n�o�zD�N����ULE�>��c�9��41Ώ5N�#֡�Z���#(h�ب��S�&\3P3p y`_�������dɹn*;�7R� ����%��@�VT��=4e��y��ho6����Oތ�y7��8�ٓT�ʇ �)��_��u�V�?5��[��j� U�2�T�XG����� ��Y�@�Q��E�b�*�^���sQyn� ���2�	�Qz��]�޸����_d5,[r7O�n�^������
Xh�Ѻ]�{,жN^�|W��ڃW���xkz�|(yI��=���9a��Ze��n��=�3�ϋ�u7����~b�l�ڇz��mC�s��J~~�>u��W��Б�~"9�:
�U1�AHd��{'3��KhƘ�H߹�ş����H/�P,�.F�y�5����Ӵw5rk�9���C�˷g��.M�������O�[5+ڞ�؂�r�������u,�����J]O���A�(���Ƕ��*�ۨQAS�M6�Q1�t(TX�轁� �b�#M�A�!]��V�h����g{�d�E�e�������p�@����oa����G<2F��c��6b�1:�,�΂p��Z�ri���pC�*�E�c�5 �H}�WUv��las}Nꕁ�,��#3� �v.��fQ�px�ӨA�w0a��n���j��W��)$ВQ�ٍz-��k�u@��6$��L��@P8�gj��>{1s@�AVĸ��FVn��޻<Q���b�C��S R�A c��8��V�~�����;�=O�2��y �5�ϑsN%zf�}HhL�*hjW9�ͣ2 �β�h#��*���W��7K-��X���3:t^�Dڰ�y!3y�;I �e�1~�Q�u�ǉ���k�g�؅�RˁxIZ�G�X��Dv���� 	��L�'�=z��h?��y��&7�g�
�y<��tc�4P4� ���	ˎ�"xEtW'ډ_kƠ�7+�N�pZk��jm�T8��	�Za�I��o<��>���T�Zi� L��F���}wb���;�_ʦ�#G��C�_��U�T�Z�r��ØcGSV>����k�|ĭv�����O�7s,,_�����m�$��Z|1"1����A�P�=��%O2���1���~
侗�`3�KyB��6��刈���`��7��A2i�`���ia����i�ى��*��t?5j,�U�����\rg`��6��K�,Ҍ�V�ew���>?#�\�k>y��$P��Zمa�y����3��}�����\$�8����b:�����j�v�)�,��^^��JzQ��1���i7�v��!(�r���b��n�}�|L���'5����KO�w���t��>���j4�H���~��d{��)��>ȃ���&dfY9�Q��.�E�Ұ�ZD*� ��IH��C:����7 삿�����>D�Z'� zݶ_ʀ�s<��/F%o�,�čpm�C�A��Υ����[�)�06x��eGNh����}�Ԑ�_�t��}o#NW�h�|��?Z�Iá{��%�ј��:��M	��N�vX3	![~��󁑔QÑ�_|���Z��
-K�:��@����m9�zN��Bs"P!��iM�4�Ņ�v�2Z�=�}ϫ�p!��EQ
�^3Oՙ��T5"'�⹣�+��*_6"ڑ�h0]"[D�J�+!�в���}=9O�zR�뭀t9�fO'���Ѣ�����xx4#�����BLE`F�X�͏�>������tTY���@Ød��t�M�-n�v*ԏ��W�j.���:'�A΃��nA7G6��h�r�5S����Z�uE�z���}�D�|(�N/Bt9�	zj7{K��J��]�#�0A�������O��H��y�N���k�]$Q�RI��K�K�* ĭ֙g�o����o�J,��a��բ��D}��,m]ƍ��	�����,r�YR4w3~��^�㧔1j\�#N�jP`��DU��.�j�}]ge�l[� �3��p+fCa|�%D�m����y��C���)6f��sG��ǲ�p�Q2��V $|F������oc�>�� }�����d�[�,��Qb��+.*�te���؈�Bh��UWf��<�qE|�Ak���ŗhڦ����f_W%r���ff�7�yo���;����6�f_3c)�zi���3�>BC�p�B���Ըg����w��Q2"E9އ��0$F�y��^
.�ն�Z�;k:C��ޮ�l6'c1� T���{�C���I,1 �|Q1�9���P�1xb����J�닸����N�SOL���𥙸�["�
&�Ҫ9XO��:Q�`$)�̰x'�0�����ph���yW��E`h��uksq:���j[Ba�`G���~6*U���n��
V�+�gyw>.]E���'β]1���}����{0�-�I�=B�: �20�=�WA����`^냗 '�,��eu6�1x�;�Ȩ���U�~C�g
S_��d���U��t�v���%�9>���y��/Fs�pd[E�M�m-���l�/�����,D)c����ձn��L6���D�^�hA�,8��b��c��xN^��e��<���O샩 ��+��?��	(�TL;�xl+����� >�;o;��F�\rmKUR��C���Q���Q�����z�f`�`8A�s`�G��!���I(�?�oXM���?$��T�.}1��D�¥p��D��L)LLe��	��Jc�xj2X��Hg��?�WW�Vq9����>(��de��(��$,rX��)�l7��a�,D��~�B�M�{��~���W��0\������.�E��!��DoK�vT�-�ޛY%�c���&ã5�����?�����^F�S��PC���ڗt%������H��ǰ�S�m�G��5HW!��8Z�O�sXv@Du~�@�_j����'�mv�2m��}��(q;b���5�c��i<�:r��ؙ2EOy.�w�H�u��zHh:������[�2a�ik�h8	K��i�����Snd��F���@,����(*�ou3$4RU�W���K�#�r��({Y�7��_/F��Sl��|���kO���w�������Ժ� E�lU�%[I%j�����(��u�`t.�����~N��ʾ��*�֣�����h�kK�Ԇ�9+u-�r�^ʐ����e�B`������9N��MÑ8�;q@v��!Jm���q[`�_{xf��E4D����鵸,��^�s�ϡ�$�)�V�Ӗʭ�����9Y3�ܣ�:`�ѫ�0�iJ6Z�^��靉���;Q<�(P�W|tK_ԗ�hnD�c���7�!��,FHO�;jq��.�]"��Q��/�-����S(��1�����%�mM¦��)Oz��b;`5�=�N��K����L��|����`�0J��ŝ&a>+���Ț0��`��	����}˄D�pm�qA%rw�h�I����ե3孔��H����.�T_܏��0�t�̼:��U�EL�H�.C���@8-W�劦�{-w�)��!mi5G.�S��E��6⼟_S2,;�J�����ۧch)���)~�ëv�h�6D!�����D��u���� �h}�����p�n�Ҭ-.��4�>��+�������_�I\^��P�(Y���0̫�َ�1�*���� �Gs(>wو�5���n��.M5i����g�WD]�D7@0��SA�iPό�f	^�ݡEL����IX��OH��&ٍW�([$�u�-Fяܳ�#��-.�g��r�y��e�g4UF�-R5yl%��!��l�w�-�a�%ȳ���?v���əL	�#�����ј�K4����t�()d�8@�V��#(�|��S��$|�Ub�lSx�K
{��MF�PP��f�،M�N@k�Rm�����[>@�"��Kϯ��}��ԴK o"H�z����Y�[�^)�~�塋�/��n >��#�����x�C�њ}?�0Eku��v��oP���gxA!�N�Έؐ.a*�^a�c�Z�N�+K�/�d�HV�I�-���RSƋ�(Y&�M����"e���šGs ڗt��A��qsm/ٱ!SSz��t~�^�uP#��XU����{��E���~����`�
���@����6k�"m�P�Du���t�ī����Ҕ��ǖ����8�4���▦ ��La�^�#{	����hP�;�Q�D�K�P����G:��[y+G�C9 �Q���\��Ɲ�ǜ�,� Gn�3ҳހ��T�4��L�N�¥������P�O�y���bv@aȩV
x�݀�����w���pu�u�90���z��$����\a*�!�&��tA-G5Q�Co��/#U#wўʥ~C�I�eV��X���������aK�n�� ?����V���]_�jP&�#ͷD��N���i?�&�o�>�	JP�:�p�Ɨo��������D0��ԫ=�\0?P#G��M`3( �m�*�.��f�T��.���c8���$�܋Z�·r;���._�ҟ=���!�1�&��&�Zt��u��yu7�<I(��Szz��������\�ND�{|߿���A=_���d��pNE�r]�y	�2n��,�ŭ����TDI�T�a�[C��5���(\x�7�(�*�#Km]���	U��k6�&�e�hoV�g��	�5n6�'it?ǩF��C~0H�!B���W�S���$��ȣ0�G-#.n���دs��:���2������R�&�Z?�rq����;B@xz���F�Ma���u��J��!�-hs4�W�DZ,�D�ބ�=k�h!g�>N���v�F:���r�A���is��=G6A�֢������Z\�3��3_��咇�C�D�x0<,� fe����qR���ah7.�2U��vHE��x��#����do��Ҹ;��Q{�R7g�8V/^x���X>�HL����˵HJ��e��m#s'^=x]]�����Vd8!�*oU	��#uB&������u�1�R毺�}�S�"��v�!��T@�-�J��@�l�&4��}E��u�jP�o�
���p ;Z�7��	5v�о�9���<�<ƒ�]1�``֫�Љ�-�8��6�d�/|N��4g�߇��>�pc�����[�	�0#5�c/� pbDՙ����id�词�U��.&w�1�Xb�hX�?�fRaY;I�_@G�/q�z�d��%��;�c���F�>��$�.ҳ2�a�!����`C��d� ��!�̺0�C��YU�P�j!a�*Q�lc�ZJx	ߕa��b�����Hg�_�M�1�^��,k���y������߼"8�S�T��{�h@�����R0��e�\�#����z��O�,��Cm�]���>	��8�$@�u4hBR[�3���f���������O����/*��1)
*�Y��nk�3��HL z��
�ީ���5b����?���� X�C�nY�����b�NL���f]D����]�kr��܀�GMb���r�����F4 �'ު7����G���?���p�5�Nmn��;�%!4�M���G]���8�h6��SP`���ks9�W�C����id-����5v��M$h{x?���PA>�-I���q0fn������I#I<#l˱f?Q+�8f�6�ez�1s$~�X�*ᙟQQ'Y��\��1�:��\q�Va�gL�R9mP�Ͱ��U$��u��CR:	�v%Bb�:w��O`��U'^��j�@VG�;�Ӑn�r��c*!%���<b�o�=C����Бۯ��@dz��u8۽��G���>�Nk��:+&
