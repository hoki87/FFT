��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#���������l��U�~�׏O����j9�PY���`T���x���s����uí������P��"��b%>�1eτy�<�gܰ�N�Y�	� {��I�ɍL�ݫ�G�R�k��Q�!E	�5E��.��:�͂2��y�m�-�.E��i�����YS�
��@�H�ۼ��nD��Y�l"BU�.TԊ�=�-�����q���Ǹ��j��ԋ����tr�a�ٵ�]�b	��%�ɔe�)rYOjX5;V��R�������M\�	D��ҏ����9c=�Vͼu��Ro�P�Jf�tRvsY��c�"n�XO��	3g���Q���^�Bʹ�7gQ+Г���$�-��t�8�����A���<����l-��*�|d"n��% Le�]�z�ˡ��Y $�v����z��Η�{?u9�\CT�J�~}o����ܮ��q�2��V������ Gږ�LK�}_�YF:�}��v�U�]�	?U#$�M�;��GT&n��K����Ń~^�(A�@�p�fy�&��*�Ƕ}9H��k�K�dFd��*��H�i\.+ג߉�Y�(��`���5�㳴R����vQJc�h[�;�B7�����b�:�0�����˛�G����|�;H_4�P�O��Ғy��u��ㅡiR�_^�Š�y�K���JX"�p�j�_kȱi��Y?0���ݍCVӅ�M7��B����<ǉ�p�GPS����L��oQ�d������ ���,|�A_-Ჴ�ԓ@zm��,������ft��
�%^���QG�������� }q����&g�=���5<<�\�^#5:�צ.����u:xͧHW<GC�"�¸��,��3$��oF��k���ly/�yJH�c�6��UT+th/C�#�� �U���9�p1Y�X�t7�\"
�g[��:qxt���̌}�����@�%�g���}J5s.n�N����'2М����5,-��g�t�%�	!�KC|�#�Mn�J�t&roG]�n50���FnQB^�l�t[4��h b�:̣���E�71���gK�݃�.א�
��$]�ɷ0]t�=h�(1��,S�˂��IV|���S���s)���~�*�:���U{s�|�d<���%��Yg9����%5�G%�&�~����x`�;����J�����d&d�9���X4�n�8�I�F 3t�7 6�"����?���z0�N�;���r�f�1�0�&���A�J�=����hZ|�����$؜���;xV���&�a�9���4ɐ�����M �'�Ԁ��Dg�J8�4�x���S;ȉ"���Q+dͬ�����s��K�ݬ��%�9y�=�w3�F�f^�1; �mZ]b8j�c(��5��-�ޒ�/8��2o�w2?�<��Ǒly���%�Ѝ}�Gp]Q�U���`�ǵM��&��h�{�;Ym��hk̚"l��-i��$�����1�+�ͣ�;-�B���#�n9F�c�꯮���DP��'�r�bEʬ}�j[�s���.�v^kp}�h�_Z�PΤ���iЭ�(ܳIɩ;.� �n�I��k�����p�� 'c� TW)Ѣ#4p{��t}�"Օ�B��mI�Q7�MGg+M~�ۋ/��U���{���ݷ]�T��{f&.�}W��͞�ͮ��b�V���sg]��5�����C�S�3,�,�7N>�Z�!ȳi6�הh�_�(M�A��zH������j�$<�_v��ݥ6�s�<��g��Z���.$E���/:�VF�����s���1��3��pT�"ss�iN&#�FMH$2 �Y;B�}�N|RO�����������r�({}	Hn�w&0��Uj�-\#c�.�s�ȑD�#��e�uHv�'���|�ڳ'�JF]�����E�ZS�m��W�%�!�����E��i4��FU�t*\)��m��dK S
���N�o�{��5蝔�<�J����GM��K��l՗#J���z����p|�r���Ub.�f�9�\�G�f̗w�c�Ն'�8RÔ�R���(�gM@-��|̵�-���8�f���RO�M2�Eݯ��=�,���I���[-[��sS���]6�~�U�!�%/�I�!Z=��u�&1�y��R�u�g��Z7����ݠ2;�� �`|�7>�S��LC����$��
x�}�!^��G�g1��g��F!����A4~�z��Cp��pMN�I1��g���`��)`��D'�e	׊�0k�%^B�Z�r*աL�s2�	X���d"� �*���_>�����m[I����[w)��HMnG��D��Օ��t-axtr��B~L�d�n�r~� B5�a�������+е�?����,��7�J|���hJ�
�o���ղ�L\���������r�g�g}M%\�Cm"�J#J��;D�0��������ѿ�aA���z�h�mB�F�b�ʫ�◜R]�5�;���o����W%�{�%蟥�Ox�Ȩ�|�<j3�ދ�뤓�_���ҏN
�pS����P�/�����5�d�㊌	�]������R�fe�n�#;��!�v_`x�����u}ua��"=j��;���5ae��SFv���2�c��G �M9D�֫Ѳ��E4��d$� ��'�Ƚ�S՜F[�+0���v�
��Ѧj���:|��1ie�:`%&a�C��� ��无������������1�g8�d!	���
�N��(�RB�t�l�7X��S��u�U�0�[�\Ӓ]��
�7~���
w����ߊ������4�֖��k~�?k�l�F���y]���b"jI���	��)���X��"�d˓�d�j]�IO�mM5�{���n�	;G�f��Y��Ÿ�I�,Pv�3�����U&�}Ǯp��ba��)�fۈ?��%��Fdv	�[�o�
ӱ^�������w?Ʋg���5x$EBL��]�?����3��Z�7ܿ�zb�=����f��O�T(��n�Ϸo%�nZ�[��[5 0��C���i��'gG2CGw��~d���%c���E\8�d���������Ndt�H!S�b7�H X�F����8���Ɋ<d'���L.��e�.�]A2�D܃�1WY� Gu������frD�/�ҕʽ�'xKl���=ŵM�t��a�߁�ԄÉ%#��p�������̿��P��-s�RӴ�!eg�޺n�lݏ&;�ɇ���z����3�	6e���,��G���H;��$�`�S�-Pl���<Ʉ�� �g�dh_����3�o`�j4�1u"�9P%�@:oMÿK�mΙ��YA�$���bC�����_*�@�o�J'�bu�KN�?�O�!�C<h2��W����7��ޭ�ȕ��~Ӗ�8I�߷tU�=�#�y�F3p�� �a�H
���z�葡0���M{��?�~�6���#ɩ�'E� �������fz Gr�N�����z���(�nSm��#W��/h�/nԪ���͂�p�C/|�9z����.���?��]��=_�>�P �m&�Sd\6nD-q�o�Ϝ�#�0u�g�౮(T��s�k�q��%o|2��ØY��y��B�����t]e�1��s�����;���YGD��T�RrþJ2�J��9������D����p�`����T�D�n
�gs����l����.W������+-��;��9���Y�oT�Ǹs��'��ى�Ty.���
�(�=4G���9�v �H����W�����݁Lv�����A>��'Ȉ��W���|��jZ���l�C�r`�nd)8���y�;��
YZ%�_�i��żf����]����D UT�dē����A�Z����I_�5�|��������U��I��QZ��W��{��sB��w�̌u`}�[����?�J3��k9�'�"
��?Z�*��U��A�,]�%gr�tʘ��ΰ�J}��y����iB�>O�Ɇ�RB K$zt�z���9� ��X��Ĩn|O����e�#W���
pj�\Kb�eo(4���9�QȎ�9�9;#�xc����ধ^��B�`��ň��b����}U�s��� V������
g1���ˇ�=t�d�E����-���d�����JQ{���l���=���  B���/�e���Ƽ��|��;�Nkqe+��fh��w�!���eI�L���b�0�w��slw����S��>�@)���ʈ����l$����3�hI�)~� x�d?�'
q:	�-��.�q��zOHF�H�3U^rlh��Z�G.���Wq�&�ҟd��ɩM��Ģt؁/.���v|����ѥ�ԧ>#NqN.��O��^�uA� DQl�7�0��������)$�����������ä#j���moP(����7��|��<�䭜�]��;8�Q��.���V9������/\Д�x�X���͒L�7��Hb5�=���TG|�W�A�6~�t5P[�ꊦr�*^Z/�E`��:���;P�mG?)�
x�T�b>�o���.B���S6�|[aE�����
���%9���Z�u�V�ۖ�Xe�%�y�n9�62�K�]�$��.B�����'��oQ->���m�ޫ��]�����!�=̢�[��"��?o�ފk:gA8BO�Sb�_tE�^AI�̗Xt�c�P�?�6l�nKs�m�4�4Nc��S_l��/��e���z&Q�L>$�(5gY)i�y�Fz�v-�����d�t,>� b�es�I�6� �MgLY��/.����exkR�1��/:c]}����;ۘ�eξo��v�ND��D��n��;o��%�α%ϑ�?�9!�kf��QW�[�pIƈyl�������I��#���o5u|>�%�fu�5�2���Y�x�N�N��C�?����ݐg���O����aF *��&]��C��ã�
��H"��9q���xކ)���.�/$�$SEE�������9Y+��NnP�t�YA� ŶҠ�Y�Yjz��r��ޘ�.v�Ʀ�n���!nv��[] ���쁲<��-���T���gW�3mt蛮3<�*;K��?-����j�B�g<�6�?*U{t�Q��X��B~f��8�q�e5���3[	��ׁ�����$뼘e!5a;�R-7xQ�sd,�h]��p��8��W46�"�,�K}ꌤ��������i�>�N��tǆ���i��i��}��x�r�d�9��^�m9�/�Պ�Z�{|��ΰ�d����^BI�����/ޙ�A��A��B�+7�W�LV74i�4hF8!��C]s�OWR�/S��y;�Z�b+����� ���+�=B�ks@���[u��|K�e�jÎ���/�(A�����^8T�!��	�,�i�B,�z�
�`" �e�H�{�Żf��������̱,"?AR���yj���o�&���:yC�^Ț=��Y<(�_�q�	kTCo�e���a��Q�{�!4E��)����[Ai�����KO�יP&��-��ި�T�������)'z����|t�͕�r�^�ɸ	�~�����5 E{�4��9��xx�R�3��2d<oJ*0s�%w*�Z-SxJ+3`���rn}�X43��[`�A!���N2>�S���0�;H�Sm�����D�����.��J~m�y8| ��uA��YSXg���zB�"Z^�Dr�<I�,4Z�㺱�f��zA� �1�e���������:}E�Ju�j���4���&��0)�vT��&��l�T���*I��P�H"��@����U����q(�g�8ǬYy-��_�<2����a�_mq&%�A�λ����#��9zc��"�5K`�5�q$A�y����D���'"$&0ͽxK�l^l�!	qq�Ĩ+Ӂn/�'��P�������?��yW~��z-�$�5u-�S�6��d� �]�����v�em/6W���|�tK��KXcO:kþ;���ӳ\�_���6e����{��gn�L_��(r?!	,��&|��j.{�p�!A����skb{�����kI*Gx�A���؇,��u�"*�:�?S�����@�&�*����w���!+�(X���=�=�8p{��P����hYDn��.����Ͳ��?�(3{���Y2�<F�b��Ɓ��Tq\}tV[�76��w��*i�8���%�r��/`��)��ΐ���N����Ҍ�Х7�n��i{��f��F��+��K�r����nevz� p�'5M�uD՛�(��vs�u᥂bM�>˝���I����Ugq��Y�['��!Ƕ���k����P�F���k��l�М=v��Wl��	�Z�O�:U6^|�'0;������E@u�
7�^�\N"�S��8��v�v�Y�Ũ�q�o���q\h��*�j��#F72�RJ�wA��2����%⟮ ��4��qo����0��Ӟ̗��rܕ���)����-�~B�cfpڧV��z�CNM�Y���;u �����Qy7,���9EY�9�E�1(���;`�!��%�R�.��oށ�7�싵���Z-<���w ��ј�Di4��.y�.KIc��uw!=V夾�����^��ACoV���fZc�E�����U�J�;��Q���W:���ⶖ���y͌�hV�ծ������Q��w��Q��`��*�Q��a���Z����y8�n�O��N�Ȝי�=fL��>l��Ly͞$0$�+V�T
�/�T�^��@~�EAI��?�����1j��4〃������|~�}��'���d��*�-L[{���1���X� ����eϼݣފ��'7����)j�/�W�����'�.=&���"{�|�"�@Z�fa"�n�+�s�e<�$W��~i�b���1:J���W��P�$���L���������uN��R/q��f%Pt�*��4�06�?ݽ�]��L�~�V�Q*ςq���\�-�k�1����������gߩ�����vу�En*Nm)�@̜[���+�K�(���$�UZll^�k:���\�?��Ko�Ӂ����k�p����o�^�wz�zM5Sj�~f�n!�,�
f�KD�,
����,o�=N�q!�8`�b=Rճ��,
����np-]3�ԙ����J�-�^$a����֓���]pJ�v= an��2"&�D���Y� B���^#f4�W�)˘��+��]{kv��S!򲬹��I�w�G ���� "3�CS�i�)��x���ǌ�2Ի�,��͊�)�nP���Yc�c5()MHtp�Ԗ��5!p!ȧ�֙[��l�|*@�"��'��r�����X`��p�h�Y^#� "O�gm���g��B� �åa���+n�xn��1��� (ß!I'oL���+\�=m|��ﴔ&[�7h,:��yLo�:�|wƠ M�4�i�W[aT�u���W�8B�#�cE]tf��ǡne���Ó��j��SI=3#�n��?�;�Y�T��LJ����裃�u���:Byj(���_ࣁ�fM�	`�Ly���>u]����h�?�Ny.�O>���Q4���ɴ�YjOze/�����{BNJ��Q���'3k�IN�k1hȥx�ھNek[�?�?_9�i��E�3�<���hD^�яXI}&1Q��d�{v�Kg;bdV�wcw��qL��`1��N�4��T����N��u���Q�f:D�9r��Gx%���
���?4�8�n
��@������2
�O?�����x�G�r���!.��~�[�B;�n#��%fkR��m@���^[�0�����1,h��6�nUq@(;�}m�JB��d��R�������'M���}Y��Eӗ�tB��|̵ᯧ;�y֖9P��q�C�"DP�G���E���y��
����A��]�B�V/�c+��mA�w*?��_�H�ew�v��"�Z^�|N��ĩvo ����]�7/�����G�����̿�]^���=b����F����9Saσ�>���I ��ʟ5�-�s[�W"B8��9����t0U@�
����U�Y��Ƴ�/�	8˕��L�����
�tPW�Y��'��g��nqzk�WI��9c��3:�"�Y�y��LCI!�z'�Fh���'C����t2��t%�%��N�h�b1�f�q���W�n%Ʋ����G�!+\D�XI�����8���a��9V�3�E�;Ӫ�GC6�p%�KZ��aNe�%RDO�~�r����y���H.W��w�ʷ���Ƽ��r�-�����نK9�����@u(C��N=�4෼�$���D�ǹ��8�^gm�}#گ��g���줚��i_�����(F��r��5�h�=(�K��u�h�M���1 ��QTD����/�j�	)MPjW�<<��3����Lۣ���$~^�>�<����2�6�}����|�J�G����x�fw�27�TvWU�HR�Q; ���C1'ql�t_<����`*}E��A �(%S��z�����������[����|��٦jn:@l�BbԘ3Rv�l���ώs���
�^� �<t'������f\6��aRخD�E�Mi�2��#(��|�]��Ϋ��|XE���=��@��i�+�,K�88�;
�w�g��:j2��" ��),�w&����8|�I4�;{����h;:���Ķ#لi��/�k,��:A�'@>>[|�nL��;��$M�6ǟpS���pLu:џ�B�����*��L<�`P�v~̀",9(�nq۟="��){�8n��R=� :X��ON�������>+#�ew��s�"����6��{qJ��Ya�>�ɉ�,�Ѷ��W���$�$l"�w	�$�1��!�f�PG���<�b��윁T���vI��L*7y�C�CR!���Ȅ�(.yl�-g�GH#"�aS'�MڥnM`[��2mK�e�C��k��6L��a0A���=G�l�ΐ���5'z��+��M��eot�(�f���*(���tϒ���QY�p ����tt�^�f�����MJ�#���;�j$�~	�l;vj��V�aD�%��èjY��+ऒĞ�@�A��6�]��?����)��L	j�w��+_�h�_�7N���BCZ敫��!��������@)4?�R[їڦ�Am���3s?�\����L֚z&>9��5f�,`l�9[m=(jN��`�+;��W��A��m��d�r��WM�Z��@n��ё��@
�p�T�p:�F�7�f�)5-�|��Z�({o:�w�@f2j��"�hf�(�uç�;S�>�Ý�c��$�W��Un@���t~�탆P���@Eѱ[�������~)@MI�����h�x#Zk��cfmc�j�D�ܺt
F��x��l��窏}e�;��-w�t����_�-?�vi�v�\��k4�6x �/�-y��޺���o5$������4����G�}��y��|<yIY��a�	KK�h�.(Pbi�6�v� �r�����	�ԙ;��� 5Ը2,��QCB5���`D??1���N���F|<�1]��O�m�2����z�`Ʈ[��Lɕ��
�e��W�yJ̭���ȶ�¬B�)�G�������D��G-n��8Ѣ=���j�q`pXCip�	�AU�xa�7A����۪���}81CU�|b��"���-
���}%t����h�-��iB�N����L��plQ�Х	;�����~�No� &�{���,�����YHX���q�Cй0��	�*Ȋҋ�������e�O=��׮�ӌ�0�_y�l��+z���+PQ�:bW]�r8�C�k��ce�B]$\p�O���#���y������4��`��F!��m�[���X|'�E��+�Ⱥ0`�?�לm''�;)�cL���/�R_[�$X��݉9�}Xk^V&s�ٕe�$�d_3����裲��?�=�P�>SN���^�Z0�|2�!f��D��3�G;w���$-|p\R�֛��1FPŢ��(�kCK���Ǩ���,E�@Xd�k���a���C F���Ly�g\��_�v'�V{U�`�6���iSc�@�P�Ck�G��4u{���;�ʞ��N[a���@#D(��-�7�� W�jo4cY{�+K��8��@(�M͹�+̆
�m0��zS;�V��1��&��<�%��BI�����݁��k�F�1|W�	.�s�#n�_y��5*���v��ڊ$%������*岂P��l֡M� ��,'�v������yPͯ���h�CrL�(�c��"��j;Jk����T����)A�ٕ[���ξX�������+j�:�)��b1�F}r�z�ݞ�ұ�H3 ܡ�r��KC&iEjPQ��BzW-&��`O��!�λ=��q����W��y�}+[�������Ux�]1Yć�"V:v�6Z[����G"h�ݞ���o�[�<7���h�b���s�;��8r/��/���]���5o��d8J�e�	[�E����H������b-�rh1�k�"Q��׎���H��U|Mp�٬ű�sr('0
B�Lt���b�A��W�;c&1��,l%щ1����:�~>.��8H�P��f�A����_+}�$!�s�'�/�dy�=�sX��s)^�'d��o���J��G��;6*_p��b7a�| Y���}����%笿�����[�]u������P�L"�W���>]p���؃K��uk���۩�qa�d����UE� #��ڬ3�[>�;n��=P��H!����ơͥ��m~�Z�Qt�<m�%�E�l���O�1�V�My��O�6�34kR���Y�'j��׷3sY~�\u m�3j�IڢϠ��ZG�:p�_�G�nCJ��I���x�����ڬ�8 �t� �gR=>|�f�Ģ5�C����L�xY�}�#�x~۩ �� ��ws����4"�6�lV��@+̵�ʜ�> ���_�ʸ��V��S9��kX��k�Sc�c��z���"�[���R����_ $��o1���T���=�rk�a-39Ձ�
����լ�`O��Q��+��-�C<����F��rN)�g��I�2��f/L�S]*�z&1�u5��rvo�b?iA�������D�:�m�BA-
 ]�b�ΒZW����J,��|I��i�0��o郮�̃E:L�X. ��ё�q�(�u 	��R�xq���UO���b(�At�g�Œ�(x\۟�~G���fBT�'^g�^0��|*ѩ=BI��G���4�+u��}�6���,�	FS��IoM���I��žzd��=�ݫ���%������Ch�(`I���㪛���<�� u`w� ��A�q� �N2A`d�Dc����UL�-�nI�Y���G�`z��$�6�����&�zf(��W7!�'�_�o��`יl�R��M;Ʈ,�k(��R�b��
��h���$g�6i`09�S>���L����	��ױ�LH��_��U�6�|��t���A&��gx�!�[�C���/
Ψ�����JC4:��)�_��9s��sX�'��<|)�e���jRG�%�s��&Ҵ�+y�&����*��$ٱ��F奆╈o����؀�I�ܩ�w_�6�V�ˏI���3!���L��i�T*_��%�(�zg@#��v�1X^��:���:a�`����S֙�5Q��dԆ�~&%��-�$��6�QC���M7S?i����i��Sv��ӳ�o���'`�O󬄿��?�b9XL��c�	_7F�
[��C�!��
[�u�����B��3�q#]��� '�33Ԁ�#q�Ⴏp��=��+ȃ�aǻ���*6���߶Y}(M�7�N�W�Z7�Ute"���	ִ�t�fZaE ��K������~�b_u4��dS-K`Ҷ�G(�v��_f�=gCq����E�O�Ɵ�TI
--�jz?w7�)g+���Pf��_��IN��������������B�ُ�ީ��U�f)����)d�B�2pl���J�p%�z�h}^t�ci��X�YLLةHi���n�i8�@y�jF�<ݜ��jjٕժ�|kԹ�8��"Ո{ʓ$���z�7�Q�밻��R�}��ٙ�������3t��/�c������Z����-*7E�C�t�|Z�L��/�4a�;[۳n�S��'X���e��}Z�{V����q�r��M�R"D�����0;�&�g�~aT�g;\e�����2,�I��C������{�S�I�%b��wh0��?���7�C5��S#��UtE�t�>�̹�Os�w
�ڔ�Lu7@[��jD�9�9Z�����k7�~t�P��}��%G�u��#�ڇ&����Le�����Y���!O@�ٌ��������Ώw�z����=�N�n���c�ܹC�ߩ<��/H�ߪ���*Tu�j�z�yg95��֓Ѥ���3g�A�K~�*���[�^F����j�w֮��4D	�Zr�yRX��Ffv0�n_�l@2�J�%5� C�Nł��SY��a;�!KWӀN�3�g�� ���x!rr�!��*�kG��E��ʾE�O��QT�h���.��\�G&P�6��gwc#-�;�I�M����`�'���.K���:yT��w��o��6����p�8���_�6^'|�����4��/#��ay6�O'i"���}nmŭ���p[|�K�\��F�����z�m���g��P�6�Xΐ���c �%>C	� ��M�����9�g�g�� �,'*������7�u���a��y�뻖F������c7cG'd��f:�Ƿw���&��ݷ�1�.�����bޫF\kF�PP�$lz!��m��;.��?Rsk�S�t�-�cWQ��Eq>�/���gA�����ն!��k/�@�+L���l��o�'�^��M?%\jb��F�6�%��Vl��8nӡ	�����1�I��æy�qp�AI�, M��T �o��G�|?�oH�p���d�=�D�X���px��ڔFU�xyQ�Z�p��1䬸97�=.�@[��9&���"��������zB8�������նZ�F{��]A��,�ڈ1 �s1} ���ÆW�wb���$z��S�l#վi�9��	\�K�������Ͱ`��+�*������Whw���B��R�%i�7�
�ޏ�N�@(��;H�L���[����-��*6��ͷZ���J����9oƂX
�t8UvԐ��?�J���Kkݙ�ӲYG���Gy]�/�ܲ7��-^OS�^ޔ��"e���Q�
Ϲr��f��݋�B�4��1f'�h����Y�
ߒB��[�T�?B��z^�ĵ���ɴ<�6r�Y2��	:/uue�6ڢ�,U��OAx����S���7��?�+%�L`�BjOD���2X`�?O-0�v����u�!�C�bQ�d�ӗ��V�6���~�N3ro]��e(h��[�`]���XA��Y\�15�=n���G7D�}��B/�a'��b�\37\����*nnu��y��Y�q��i��~+Bf�UZ8TS�}��q�C�K��y���D��
n�%�
k�2���:Tg:����3!
'8>S�.uaV&NS�.��<Z�V4Îè�"�T�E𫅮����w�F��M)������B���r����?�|DS�9�:K�V [j�]���x>��M�����Y�X�b^6�ʥ� ��M�M/���{����?݈{��i�\&��E ĆW�ek���T�������ّ�/�'�}f�����Uy�k�������.�N~�*4�v��)�	��L�"�J�ćJ9>q�ۏ\k0��C�͘���"�JqbA���+�Ȯb7�2f�}zQ���Ѡ`���qU`���#p�=���<�Ȥ��~]�@/�����D�09`	$�\��:c䑪ݫ0Ei��n�n'Ys��C����X�t{5av�1k1*���:ܳ�d�.^������,�;�6�?hA���n1�CPXk(��9�|�W��Cb����^���3ѱ�s�E����JPI�(VKX�A!��|�X���T��?8�!5����)=e��ܛ�Ę{%�'�AMɿ~� 92F��u�mm��ٚ�S���bf�l5]���A0Z=�J~��y����61���X��J.r'�ڇ����;��f��*D�{�����!*�?X"�^]�*���F
�
5�8|�L�~"��B7[���mbޭ���>��Y���p �8�������n�~:����a���R5��aSQ�e|��V|�3C�)��踐��#tQVE��-i�JTH�<���-��h���P��a� þ�b5zlA` �D
7��\�"
���\^��R�Cf�Ϛ��WХ�j\��RA�|����8r�sU��}���%9������C��M�:�28�p@�.0E�ב#/�֋]�O�u��h�tK?@�����=��'�ݓ�	)?-�N�z俪��Qc��S���*�T�M��Y��d�N,s~���5��/�^�9z$��gb�����̮4��m�mn%�Td��ҥ�k ��FG�m?迟ѢXx`aW_�7�~ر���^n�)��u���-��u��-��]�]u��� ����k��;�c- �:-㑥�����kлj5i$-F-C3�v�e���q!�T���
#v�h:�&��2J�\4��'+�ΕUdSˉ��Ǘ-����(�x!a@�R뒼�Q*u��&|0�A���kL.*�"�n
���-:h�m���#B��P�;��>U�h A�ж��޲��*�2��xP1�r<�݈���3g�� �r�UX���l/ST�R�5�7��wh�>�R6�fP��T�/�tS�X�޴X\]�*)�"c���^�_�iU�yl�Nʇ����� ����4�^*-s�����Y~beZͬ�[�ӻK��(/�W�be�[DH�W�*A=22��&K�*�A�>nv��Hƌ��}=����ނ[rĶ�Q��"-��#�����` X�<l[t��� �`N�T��ǵTi��eϗn��V4!z����CtC�m�-#��P*��_���'��y�
�?d,����q�t*◬ʯj	�Y�6�W̥S�����K�E�xi�i�9	"�("�$1*�y˦��e�U՛m_q��ӫ��W~����&o��h�i�cB7O�=w��I���[ ^>E�"�����Xm`�.�seV�ō��S�Xn�{�Ћ^�Q�#�j�LU���*Qψ7Z��rʐ����z�Jj��Q|A=%��0��u�'B��X�Յ�	���@�O���d"2��(�p��?6�@��נ;��l�t��7�U��cl�6c����Tj��a�|�тR+ B����"$�P�B^��y���w�rsT�4Q��)�M���Ecj����Q���e��d�V�[���q&���'~��n�(Iy���!�߃�t�9����!.�ݘ̹�z������dƤ�e:����z�}@p�k��E�ha�Yg�MԞAe�7��T�����	��V�A�?EE�H��o	d���3��w��^�_�2C���U�'���OG���VR�F���҅T�l�Աҝy�R���4H��&S/�p�j,��G�&3�����%�@M����@ �<��T�΅M��޷L|`�A�+�I�fW�$/�F������D���������T=�ϕ��gV�!��K,&���E3�:�������(��c����Śz��ܥ8D�m��D8�iX�Ղ!��Z:�cZu���\�Q�j$f.�	���;�I��&�=y��9�ݒ��������L�M�!�ݼ�<6�BYJ�8*A�w�{J�RH^�þ�Hd��99��t��&p��4��SeͦQ%��N�5nJ����4M;�Z���z4C��~������T9�7+�M#�G��ߚ����U�;_RA�3�y���1Ch-��RF�j�&�;
I/(+귝ā�O�[��V���cs�⮃U�Ii,�+u��{X~�r����-n�&^�k7��g�x,�8�B#_��Ml����h�Z~��X�}F�Lu._Fi��l��E9��M�Fi6�� W������+[&�q>� �����7'�b�������">ƹ��la�kۓebs>���c��^� @�'����ĉ�Y�;�D8>�̝�����_��rAe=�3����Ƚ[�jd�h�ҫ�\�\�@�&c�݇�84�5�=q9���B������NӚ��,[� �� �i��9"ք� ����B�|	�xg�<ux��o�C xB(�*�7���ƶ�q\�Դ9sŎʝ����ׅM5A�����<Dk��>Z\�;\S傹11 0�^ 9B3�OJ��4��-`B6@l��s�^�=�m�֑-܀vv�
g����������B��$���mȌ@��b�^�;�FK5�r�({@Td �6b8������š��]1�{kn��ğ2�r/�_)x�,9�M'i�������������a��`^�5�$ �~��,cx���Y���bLb .��������m���{܂�T��G�&ћ5A-�_nS��v�O.J`���B�:��梠^���G��^��U�q1�S`�Ĝx��r,��^E#l3��Z��i"���+������ר[���p��.)T�9~�����,�e����q3���)�p�h��La���Ň��9�V���$.Vߋ\�[��:f�sm�<�&����FbO�%��BC�V-60|ȷP�[^��١�ձ����J�� L��;��a��h��+6�(��&���^v�%����>W(�h0�v�`T-�(�P��.uvCU?�0����|�G��3I���l�{�����%SIl9l�>���0I��
t��4��S�_Tsc4Qv��[Az��"���G>���K8�/����r���@3�f�}FWJ ��Ya�_�*�����?G���>")e�=w�{�u�MA�
��S�O�VN�UZ"�����g
�.�����1�%c��;!� ��ժ� T�+����}�kN�f�s�L�&�j�Ȝ�@'��Ay��c9��b���Ua��[��~�0����@r;J�Pkl�,����GQ��h��j�ϓj^��i�nB3k��Zl�[��&}m�i��D=�^X:v�n�w���!y���7�č��/%�|zp/~�r�(�Kt'����t:�5f�Ѕ�,�"^�B�0�&,�����D�P���,rg�\u�sdڛk���\����т�#xuU��U����HW^�qP��J��4;K���eU>r���%	ؼN�;�X��]��<��9EDV*BD��X�����,J:X}���pN�>�z)}�4��t����e�U�% O���^�r��?�}�ρ�P宓ޒ$c[��X�L�'�u��"��\��קb] �	<_c�{�Ϸ��=�WwCt��� |0�f�rj.�a2��MR���$\ɷ�+�5���g:ܴ{�I�\3����R�a�}���M�S�cŦ(�9p�Yi�\҅c$d�7�9
F�C8
Nʠy+�'��7��u���e�|N䛧�(8�
���?����;Z��>���� U��cv�v^�VxFÑ0r���J�ڽ��\L�ݗXę�%x��ؠ�A���`"��	B�&��kk�Ȭ6���ܮ�|Y+�f�ج3о�i�������((Yq�
�'eqQ��W�=��⬓��u����}�f�z��*��7P�_;����3����#�,� �|NAU�5집V��%:],�	[����YH
hn ��Wt�~��dy<) V���`�Pg+�8e�QE����?��ŞZ�i��?7�  �S��*��gA��$�������
�0B���⼞��נz�&�E$����c�G��^�ƴ��zI9�^+�Iĸ�DI�϶���
	j�?���N-[[ՑE�ࠕ����p0[�kw6�����~6�$�Wn&��I�j�[K'�?���T@U����X�$
�f��^�i>�D����'����7jn �#Uu����B�B��M����X3�{l_`*�~�V��O�?Jt����:�o�r�ɍ�v�.pm������\������!�N4�����n��C�K�����]�����z�$O�{�"NR�Ʉ�;)��]pJN��)NJ਀�4Hܠ��\��U�.c]�UVp�4Dr<�ݠ�N]����]J�~�qɵA:��8Y3�CIJ���	M��s[�L� Ѳ������h=H��%�%2��~i��\=�]����e	lc?�s�i'��gO����)�E�+�z�Ia��}δ?}V$�w4|��/����0d���X�$�Z��JM��ԶU��p���V�k�������֡�ٚ5��/ڦ��fj���I;|��\[H�͉��l��:���Q�6�!'G5W:p_-���ܦ��W��Ps��ʚ��U�fsEqR`FF�������4{��Ql䪫m�k�����|�3�H#�P��t�:�\?��>�@o[��k�A���A>��^)ߦkrKK�>v�|F�V�3j���5Iz��m𝷦��f����_g����#6�c������f}�)��ePT���%��z���PB�-b��A�OS��ܵkV!�8��p���˲;�ַRm�ΜV@�Ew��X�!��q1���L��Т�X60�s�$*VF��{�t4e�:�ػvA�[�fS��fwtc{��o��ȃ� !q�߶.��"\n?KO_n��Lv���	�*ts&�1vO���l2��]z2D�����GB���]Mo=t�m�d����^�Gq�����S��Y�~�פ�.��Z�6*% &ذ^� �pP{ϔ W�!S��x���+����c`�t9�5����Ԋ�����+�o!
�3A�ް���n�-i��u�l$w|K3΋p�b�Bp:æ:���VZW�e�A���E�\�n�9�0�~��Y�s����L�H�f�x6ޑCccû������O�88/]��L,�
.F"��=f����Y�d��9�1���\�����n*_p̭�I�0�?%�Uj�?x1I��(���l����c��<���%����g��S�\VL!}|[s���42I״��O3���Kc�{Yk��׼@ͭ��1!7cm�DD������)J�dJ�g)��vX�Ø�����,w=vb>��h��]�5�[���E�	jV67���́�a�w�b���i�,��};h7����`8I�����+c�S.�Rrݾr߮�����t�տ�Cջ��m�
6��=�?z(T_��!�X�q����h���,Q0�2���q�u��a�
�,dCA�.��3J�l�ϖ
���H�쳆)�LTm�St�GqZP�~�����8���e��/���\�#�Ȇ5���?����e���,|SB���r��'Id�!���x�Jy�|?<&\���`l6��L֕��u=���c5����.�b�@��3�u���m)lRӬ�&��'G�����p&+�`���`�2 �E�f�`���Æћ90jۋ�B�E<��V�*�2��Eg!��s5�A�s5b���苶ϭr�F1q���OvT\v6V�؃V�0��)�1O��@R.��W��&9��2dtז����'��R���bA�#�;J�5����G��\����*cA�	�o]ehbo���?��G^=�2̛2m���¾��ګK�~
,�=��	��i.P˿���S;R�O[3�VG�b+��}%H��>�<;ܴчM�e���e���XkO��I|���u&�|�zkm�����h�<o�|~�٤`n�8$-P���N"��
M!�V%Mn��e;��g��G�4<Zƣ�|��a������_���~�v�ۧS?���#6��ᾢ>L:OF$�ٔ��M�>�"�n���xB$��R���a����H�a�Q�:a坄��>�hE�$T}�Ԩ�0Ta�d_K���ty��G���l����.��q�"#��5q�R�ZR�s�6z��MQAhdY�����a�f���&:%<��=gU����`Z$�*A�I�3�eX%m��jh��3U̴�RZR���@�<y��C>���,�6������'�GG�@�����+A��if��f���R��S���&�,��0�x^=�r�r�_�/zya .k
� 8�//4jƹ�߽_���vc�R]���������}Y���D�nwe`���);�O�]
:�0��	|₌e<�S���� ��X�v]r^��e���q�5��X���8l0��aj*�?��J�X~��#���,a���H��'�akh�#��c�L?���X<�:O�C�W��~��{JM�7VG��W뿼���x��M#�U:�e���vƃ��M�ô'l[m�p�=tٚOI�Q���"���7J��[9��廊��y�3�����/G���	{�(��t��]�&���?ޜ`�?��*�ָ_�u��ǉαjsr˽H�l���7���/��m8��Le�d�C�.k�� �� 3����C���S�և��d&%���p�0��Q�r[/�\T憎L�{*��O�i�~�4�q�������;L���s۞\��\�Q�C�(W����NݬOh���6* 尘���9�m��a�o;�1$	Q���J)<(b��
<a��"�>6���%kW����䱱�Տ�\~�*+�+ӷ ���6uwo|��7���@�L"E�?�%��������5	�@W{ ��ep��������j�[��5���w��cl�+RN�6��Af���6:�Id���aʀ��9Z�[P��/1�Y*	mb��4k'��x�Cx,�'�]��ݦ�g�\��̭2[N�~���#�����oz�`���(���-�8��"��
u���=������|���h�H`G#¶P���\���Dez���ץ<�����������jv��nM��d�]Bt����p����j�(���ӸP^@UG`�X��4���I�0�y�X�W�a�{L��m.���J$�!�L#X`��غ��!����q̍�>e!�Sx�v�߄7if[\ߟ1��τ�����p8������EtV���iՆ�=�w`��wsՎ��,�֩�(��͹���ڵ�����ՁE/����������T9d��a����W�:��Y%aly ��fB�};���9���r9P�Ї�O�֗�·���h�BD��q�&*������u�Dv߿�f�����'hԀw/�\�)�Z%@�C&H���Hi�ӌW��F�z�ڔ��z�x9�Ӷ'	n���o~`��f�n�#�`�����7�h�qB���6��x�@��JNA<N�8���࿚jf����h:~)&?�}�<��X���4��V��tc6�V��/���;�	�k�����H3Na�1���})d9�^�)őcd��x)��P��X`�i��v�;���b��6T���Z�67��z���-�w�of֞\-��mm�p��^��fh҆MP*@6E1���z���jF>�ܐ=��q�C�0T�%1�1�KG����s=��>���1L�~Ĝ�SV��F��73�8 �E��Ӫc�d�~������&�Ú
]�8�ڌ�����Q�=@�x�韎�3�.m�����y��P�H��|GO!����prX y��|�yV�I�-��.t �4��!b�ܡ>����۲ N�z3��l�wL*�Ys�?�h�1c^HZ%�TC��}�9?mlas<^��A���� ���2�Y��d{���k|��ܘ�T�ff�����DUO�J��Q�:�D&�|�h���ᓫf�2��'>��~�_X� �B͏K�#)UB���7��m<�������p��W�{�/s�|E)S���(ap�|=��H"��U\��w�|(��_�p�����	���z)��$�wlj��:���*W�oD`69pOƐ�Ԅ��Pl���P�OŶ͹ֵ���^I��b9IM����5��e�;P�@�~�NJa�\�8�)��dϼ�:]���\#[8�F���[�m��ۙ�o�:����g�q��}#��"��,� ���d�:���Ld3���G`���3���KDc|�>��$��u���f;:�ڵy7eO^:p�^��f��� ��<*K^(��}�����P~9�0�W���	�c4������d����ۋi�do�e��r�H|���2;�d8��#ew'��D��I��-I����QP-�p.��_t8&���U)�΃��&�a�zQ2yw_uÔ�E��=q�L�po���3l
�u� ��l�x?ت��P]#|��w1���	霦�T���Ρ�I^G��Ԩv_����Z'<��8\���N[�o�{x��鎦[�2�(G�c(�y&��}��)�R҉]]�ӑ!\���]ju[��
w����@�Z{Clw�R� �0?��A}���[��!��){a�[d��jN���ū��]��B����cF�abb�Y�>ߡ�����:�mcZE�_�`z��i���uQ5���a�V�����LڈrG18H�Trh�U�sn�3t'�
W�ӓ��ŏ�~t�[~ݧ�����+�r怾���o(r$�z��+�o�|���)^�R����9�BT�)�q�L!Pv����:{��f�ř�&���E82�H�Ĵ"M��loO�	�����N�����i�H&����э����W�J?�7�l�����4έ�2�@�B��Y5gJO�;���,�>��y���V�c�P?�=К��a����2�w
j�T�UT2���9��L~��/K%�a">f|��ì���`9ǚz%j�G`,�aIo�D�j�����b�d�v��6�.�%�	���	�'%��i���UB�+N��*�]�ݧ�Gg��㒴iD�,���f�g��"���q�� H�,���k9�B���ӌnAS_��U�"d.)�H��g���3.{!r��,� ��n�M��J��E��0�I�!4��Z��%Z��$��z�#�\�`��-�;�.�q�dz�AO���}�����s~��6ט�"��O���3��^l4�Dt���Ec�����]nS�η�ѿ��4��:C���V&�����T�|sM�w������@XK�jz�qUW�����X�Tb�	����k���a�@Y/�&wk�mBC)�^T�#�#ND���g�v��m�̽�#=��ᡩ�qT0n������5~�`����Cm~ܬJ�m����{�e'���@�4��x�k�Ul�̰eJ��P5����������1��.�*c�}s'����D���^��~��3IU��f�V�B5�j��jo"�P.�{�Ď�7E�sIA�Z�f�a4U��>��SHGw�<�n�������J�̯����N/�W�6KIj�Wr����F��>��G;�sl��l�Q~x?��B�i����q��}ʽ,�o��G���햏�Mʹ����Te
wä��N)+#��/.)�&:Q��v�FW���<�K��|֨�ec��J�\לx�mIA��*��p&VnF���œ|�uЉgLj�4���1e���h�2r�j�:!�3���B/$x���� �<*�{��eX'6��U�~�x�l�MD��d^�^30T��y���W�"tN�����̽�V�$AJ��+;b���æ��U������\�J��l��#nl��H���`���4&�h�("&E9V����?�5�vV�� ���D�x�� ���a||t�1a�����[��Al�KV���.UQO�d���h��-����<�F��?��,��}$L��[��/�<)A؝)I!۵�ޑ�RR��X<�@B�VE9�{�L���D����eWV1/����PN[ ��N�6��)/��	����q��\.���l�����,����&\�.��x���7�	BA��S��0}��P�}���gy��L�R���Wp��[.�H�����\����.��~N������EP1<X8�y�����|
Qc�7p��קj*�=X��|Ѽ��e�@�������ו2�,8��|K�4����Y!b�\��a0~��q�E�)ѧSb5��0PUt�KagR����h&��j>�3���;c����;�����Y��/��&����H��F9�dB�F��Q��̓�޽n����s�X�t�]b���4P�u'�zi9��z.b���G�>Q��*��%����r��(�%��@Kg��/�#?�r���	���m��)1���0S���q���L{7�$�%bɚ<Q��?	�Zh�]هa�;,ڬ� )4�i����� ��̴DF��)����Z_F�޸j#�P��E9���s˷@-$Xo8�w!Y�!S��Ql��Fd��b�J�2����7�?�޴�D"�iP�p4p��K�����ݨr�`�KH[h�W�A����v������.H[p�s�)�r�yf�>aA��D�lnO-�C9�1��R9��W9�ǫɧ�p	k3:#��@Ўl�-j���������!����e��DW�rT����=B�1���`'Z�Y6�1�5
�P�%p@aH2�(F<�bAYYn�H~wh�'�5oX逷ô�b���N*��������-���3��zc��v*��N�{;��P�{U-��4� )ED*�������BHu�)n3�ţ�����I.���n��9rp�A�2�W�8�����"@_�f=�7ډ�/��Me�uN,m�L�b�)�(2�Z�m�NkB���~�����C�o��b�Pw`�8\�_V�\hw$v�8?�X�8җ��av��u���j�d\�ܖ��u(�a��>�l�^y,E{L�/���" ��<�f��ȧo9����b/����µ��O��:�����R�~�^���L+�`��p*���9�9�v=ⓤ���i�xo����~���Vm�z�� ��6������d��~���8=�kx�1}!<͡��g��S�#���ȶ8���_8+D�)��k9�����*����kU-9JF�ZZ��*`�v	68�mςy��*�x�8����'���w��G*�ݙ˶���{�v5V��>���3Vv�:5�=}���,Z��|������U��^�Xk��Bv��f�b��w��[AlX�q���L�Xt��U��.�v�i�.�������h��3�o��rñ�z��ؖ0���)����Q_#a��0�����!���8��?���P�'cP\��F:���*渧��A�ؿ���yq҈��y��!����A|q�9��/���/tᓂ4��,�+Y
d˟���!֖�������q	v��2�I�o(��-�}�-2+�0_!�6��dɋ�A][�I�L�,��S��r	h]�����2ǡßi���/�!���̺Q�⚼��M襁����K!(�K��$����ӂd.Z}�ji��ueY����qpq�u?�8�Ѭ��h�J��~aG��ԓB���^eq&�q�y�ZC���r��`�g�d�!��%�@k���*e}�CV��mnEB��F3�'��h��ӑ�B/;E���L����{���Q7��k�-p)�ؾ��L�yŹ_�?��%�l:Z��m�ΐ�i�(Ĭ����I�K����UH�'�9_�5�Ca�9- ��yHb_�2q�M�2�#���S��bwQ�>�䁄��p���'��Z��Ϣh1q(�&f�Kg�w0�/1!�-��k�{�Yc�?E����0v>�xm��ck3d���72g�xLэ
c����"�vc�R��(��s3��?y,������޻�ak˦o���e��H �
��&~U��f�)錽�e[�T��>:H Yb�CmO�v�E�aE���V]�<��t��k�![���+�_T����`y���|v�T���'1O�<��G�We��̌��1�)�j,YO�{M�O��y����9nBr�5!V�O���=펪45���VlXK޿/����獧�B�1u�N��S�O�4+�^y����������/d�ڊ�;+0B	e� <� 숊�����h�J��jik��Ɨ2r�*W��B��=���n��s�0�2�c��/�^ N1<�nA������OR�7k�-���Ss<��b�`�m��9+�GA�0��fh� ��'������s�~)!�X�����&WArŏ���4Q^��6g�7�.��b\��3P++�u���
	w�����YQ�C��Dk���~�z�1'�n�/����."T'��p��(����m��-�u�!��}��\�W�ka"�3�FO6�sȹUF�SYo�%\IC �?7�Yk���A2ԿE�=�G�z�E�d/�E!�I�'M	xQ�|*��7�ϖ󩴸�2A����U�qB��%̏5��zH��ФSh|T/MFv�d��^�0ѳ�j��΋������-�HV5�ו��+����m�xl�?5����т֍�J�0J���,���G)X�+ֵ�Ui�� ��U�sTy�j��p��(L�Y!p6�?fa��,��o���\���tt��q���"ۑ�scgØ��x�R�s��J�l����6��X��2��v�fw��K�K�.i�4ki���@�$D<���
���x�Po6�Z�~ ���ʞ ?{:�7��U�����<z���_���;�lt2�H�[߁�~�Nӣ���Fatj���Øi���q˫ڂ!)�a���H��k	9�Ӑ��M�|�4�>��sr9Ѷ�v�����Ui(Db��ڐL~}���$���;�cSw-�0_8��@sKL�kQ�}4U�=�Ѿ+8�"*J��e@z�Z�Q$oY��W�6v��/j5h/p�k�	�/0J9�,���_3:-�^��E��cՆc�Rk���Q
+����J;�E�sx=��-���v�YK�|tN�ez|�%��D���
t"�'��+�h������s���������,�dX�,&�(PMָH���^C;�S�P��r�Jl2�g�f��YtJԌ/|<�B�-����'[��ݷ���hv�
=z�UEİT�DH�$�bT8�2�[B_����,֝"�8���DT����*7�zҹ�&��
Ɛn��о�,Dc�q�ǘ�jŅ@2�Nܪ����$3����\�qA��\��q+�
�Py+�s��d%�r��_��B6)�CN�7b,b�G��5�R���Tң�\�ii���	G�s�ո�]B<���� �m�{����>O4"�+V����L��Y{+�my�4�>#V�IΜG�:��Ľ<��A��C@K�9�L�)k�̵�Q�� �z�mcb.h�.Z����:x��`(9��o���sNq}`�l8S���g�k� &�G�o�ʞ46}~�ѽy�P<�b���6ƨ.�_�ݩq<����@+��Y�;���F�vտ��G^���9�����4U7�����{ăxp�n�<���KS0[�N'��G%�Wǯ�a��`ۀ�r�7MMȒ?)�#
U����h���qC��6!�i���A���94l��-	���3��l�p!&$q��������9�zWt��J<�d���h�����Mg��q��p��}#n�AG��_n�^z�LM�k����G?Mq��ᾃ���_l���boI� ��`:yf�r���C�3uP�W �K�LJ��o�'|��u}��5L	?�Y����D�>��ss��bX3рg�|跇c�8��Ą"0ݗSk�������V)�i�\�6��ņ�M��d�P#{.e 7A�����H�%�F#^8y
���3$�q���jN?5���=8f|�K{�_6%�>�rլ	
;�I�c0ZO�MZ�;�J���1�d[�W�ĉ�06��&�n5{�i��z鷝K�ö�6]N���m䁖�\��D[F�W�v�!��!�]�h�М�NU�3��՗Ŷ9�fA{��R��`n�0�y��Ma)
 ����?=���;!�\���\ߏ?�:qvOΤ�v	�@�}����Z�f��4:Y�/�Ax�r�/�S"�E�~j��gTpo��&�7;q��|��*�����(�������`�1�.�R�a��h  M_4��e���%C�fV8,�N�A��Bӳd�o_�{G%����p>'�����8ht%�鄶����1��D���_w��,<A� zw{^A/�X/`����k��A�C'Q�t����,@`��Z��9�H4C18 1`!�R�F
��ή#��nJ�QV���3��)��c��?@-���)	��D'�ķ���n���
;F8�*�:"�=�.��pu`�3��/��HA�~�T@M����dБ`>�+��#L���S/�E{�9!<3�	���n�ԃlk�,���S�@t��zkg'�8G�B�9�9�k�O�ʊ^"��3��@U��T�P-#׻[����H�׌����(������'����j|3������,v��:�����ݢ��$�����`�A�s��j����n�h�6�-�c���<��|�����'�s�\����]����nϦ��0�{[���}��/c�q����0���&Ƈ�x"��6�@��})�k����4W���~Fz�>?:��'?;g���=��]�^��d��D%�HB�][�3���e�=�uO���m��b�|m�u�YJ�|\�����i����=1 q��gd�O�Q0��B$N�+�6z�cKk{�b	G:���Ү><�~��ick��	���N��e޸��^������CD��4K��\ _wf4��*ׯ�Q��(��8/�l�֚p D��NGn���0�L�_Z�!���$Ɏ�`+>�e
@�8��֦���U�(��)�Zڠ���a�4䯐���I��EK\�|=>������ӛ�����AyGѵ�b'Z`��]9���UW<U5��'|���U)y�/�+=��U3��8[�i�u5)�e� A��?�a#�ѱn�T�u�a��d7r}��E`�U���M9r�������CB$ؖ;*��z�\��L{,]���A	@�-�r�n�N�RQ���\.�h|ܤ񿂔Q\���?.ijgYPC�%QF[�sAX�[+m���
R��k����1��"�`�HV0ꁟ���UFIHJ�@��` �uv�\��=�����Y��v��<��5�^UkQ��Vt���9ͯ��F=,���K<����������J����c?G4�˸�2C���A|YϪ��g7efJ-U]e�_�9��N����hK��z��"y�+��E�<�����V���,}���ϞuH��x�o]UX~1�4<1�%\@:�վ�V���C��	�:˻�������x��w�'Ƶ�M+!�9�㝘N�����"8X�!Ct�/�N}|ೣ�=��a��B9ۢ6���vy��Y�1o{�����G>`l`RK4#�foo!(�����d�ŶࡶT<Ya�\r�����L�1*�kN}��\�����TJ����%wB����ؘ�o��ţjd���o�h�/+���
`'/�	�DG���`V��Rg�f���M�5�P�J%[�!m�{�� �ӭ�����������g"!&9Viq8��g1��&2"���ӡ��i;;h	��Y�O!`.�~ƣ�X��&Փ5.��ƼF w�w��~�e�*�X��f��j�P��ߑ����j��Ӿ��êL*���F�l���&���0�چ����/0�?r����`�e$�rKOB��24E4M��i�sy��	���RS�6�婤1�1�f�'�/`�W��d�N��w�﯁�~+P�<�O�lZ?3��}�5.%�a_�
��d���_�Ι�oj#L~DGt�/H�� �
A��8��_�=�sɣ�s�<�o9*=n_�/��ݚZ�;���3��ps�����7n<BP�$$Z�����e7�"!���<P	y�ؼ!G�n@���ɝ�QlB<��=�2
��˨�m��V'�*׿���4��e���$��t<�G�a���+�9l ���<��	�Me�ӑ����ƞ�\��� W���V�2�9'�=�j�,z�+p���j?;������ �s5&�)��\�8Jb��R$q��e��� ����ĝ�_U|	��7b�^9Q���]�cI����R��]��L��&�t�48�9|�d@��g'!io������"}E��Nb�DȧR�J�_0���MyB8i�6��j�_x���.��uʸ�ZO�.J�K{�T��a�Miv�n:�K��uиu��s�cC}�珗`�����|+F4�>�h2y����g���
��S��C��b�������,7����mݒ�&m7�ΣG��傯5�2O�������W�!���k����,�-�k> .9�j~sY�фj#��1?D�I�
5�mbO�7\�]��4[z�N-d|
]wăI`-"�Ny_<�!C�tf�~��v�����V2�ӭ����Ƃ����d��/^�׻6Wu��yGNiJt��������; �!@!�^Tg �%7�l�H���Ԥ�v�A)�3���a^�#v狡��*i��T�}<�VW�Uc��1�mES�q�7��j]Ç=����%W�Q=a3������#���l��%6���j[o>���m��=����Z+��ED�BrV�+��BJ4���Lɷ�</�ɩ��G����#���<�c D�
M��D|rJ�i��D����2pCN���>3� �"`�Ǉ|�eA^91vhV���ޣ!AY �d��L}�����#7	ZzN��f�s��(H�	�w�ۜ��UN7�W�)�sZ��0	�>���I�+���<�enTlʹ���d���B�$�������N	1�����EE_�
7��-�H�W%��V��/�I�g�������@�Y� ��*՗���\���j���`]m�J�:���:��D�0��7�Q�J.���k��$Y
`��t�T�� $*3�0rn� ��c�طvL�|�.Ryd��+�A��0C�lL�Wj�FI3���J:�.V+EB��n��T���P*F>�K�Bϊ�m�!��n����  �#���c{�.�-L[. ���b/ٰ�yJ����Tϝ���lLvfU2۫q#�m}��eU���䆪Y�ڨ�с-Tq��*on���ↆ=���[�29hOi�5�3�\z�`��=(21�w�!����宑�o]a)��E�9��#��@�Ǩ
�iQ����+�l:"�yb��R��ێ��D���}�5�Q ��A?G���5r�_��~A�\�#7b�+�p�%����'�����U��%������	qU�!w��o��:*�DI�õ�	މ}�*S��5��~�Tls��v3/��Y�]9���,�LH�E�q�=�W줓��	L���[7|v����?��F{�R��U��d�1s�����Bg S,k��}��Q��p=ύi�Do��*��Q>MͼE�NB�Y���Oɝ�������a �a�=4"˛d]����{��"F�A�GhV �`�nWG�Sc�F8���A9ȺO]����@x�uno$�E-�k{-���y�#wL�hQF: j9�'W2���g=Fhä����x����3X�յxj5Ql��o�b�"��~x˱�{ͳ�I�B�����`2��Sf��>|eU�n��Į���⒝b惴�b�Bx<p��F�a�ٵ+�3��v�/���2=x��G�MHI�`G�n�PдO���/�'۫q��0C�į��>�[�3>��Aճe��@��p�ߔk�d`9BᯛP_I�V�
J6�{A�\ea-)�h��xIRw/ay���k��D�V����#i۔%����g�/��j;����D��% ���M�Bnly���t�Voﾋ����,��^�������I���!�"�v�����tZ�]7��
���2���z��<7�T�
�K-��cV4�Vǉj;��y�jG(^�J��5�*���G��.���*26f�t�txs �t��� 	x�ޕ���{�H��!Q���x��v����ԁ��0����%.7��i�Z���0����9��v<ǂ�I������x�S��!Z�E��Ai�[�q o�0 �g!FQ�Ѿ��9n-,'E��#�H!s�Α���j����fSz�A#ŵ)�V��1�_G�g�b	���9�by�W�*�B�ܤ.��۩'�!z��s8������{,�ӧ;��߬e$	�P�̡�[D�U�3�?U�'$a��8|�̈If$V��=DWxP���\����a|���uf�C���"�	�rgX.o��E�E>�_����:l�5;@=��:2�O��)�K?�:��`�����S5i��t�����e��V���>������KΔT�ma�;��y���}@�2�^���rn�>�F��h	�������0F�_�n����,��Ћ�H �Q��	8g&N`���n	��ztb���jN	ʳ�d�D�*j��ߞD�m�/���L��t�MYt<��6H8�)��5��S�1�����E��w9��w�(#a#	�ܜ�!��S_HR~�Q���:��0޶�@(�b�eam$J���:W{���ʫ/�y\sv
��fq+��d>8*#X�.��]�u�Tv�t-p�,%WV����5�o�1۝��2��R ���?,rm�A���W[7�,֏�F���
�!�d||:�6 ���.�7`J�8�����M�zO�ܧ�@�">C�@V�o����)����\�$P}�3��AڍFҼ�ӭ���UB]�:�%}�hT<q�B��o肼m�CÎ��m8m�  _J�ra������Ls�^��J�)��0@���<ـ�b|%K����h��4��yg��4P/���i�G���y�� �Ģ��߸0c��?Y��3X����!�%��[��r���0 uk嵠�� h \��R���'�t>�}!��ٌq*��HF�q�ȁE�t��3<`+�}Gb �%���be!m
y~x��`8�Xd�����712����s�F���<��D'��\�h�*�\�M�:>Y� u,��d|jj�0�Ė	
n�������[Pu�fzKt9�6�E4��.�y�t8��Yvu?N��2®׎�����J�'��.2R��D+go�JżAT�Y�-�����E8t�p'8R��M=��=\��A����{+���g������=�ݾV��x4�sj�={�� ��i�~�}ڸ����j��K% ���L63N�\��l��9���i�:XU��F|�Jk�{m�RR�莀U��4�R��(z�tx�o��&L ��@��n���"�D�^���D� �兣�v)�����C�>�Huȧ�3�n$�Ӟ!��+Gz!�@�},y�A���.aj�rm��gg��·��	9c��Kю��NV�_�9U v��{"��W�DI��	a\��6.�*,��:��x��V/B�wx�_����P��b���y=����N�GV��28[9�HQ���F���͆���Z��qE�q`F��?���2���$�_A�}U�5/g���%ݹ;���-��I���0�feE�p�(���T�=\�5OCBjD)�1n�JMYvj\+v�)�jȢ4�BE�0��q�
jԟŢ5�,Rv�@4��]§�O&>��f��֫��4�s%<W�ڑ�����{ж����� o嘟��9��ER$��^R�e$.��4�픆��h�dU������J�)��Ϋ�.�jՉ���(Q���\ĩ�Yfã-�����wԙ��<����Lf��U�{ڴi�)<wm5U�T����ULr���9��H��4��':"�2�m�;
f�|il�+ �ݣ[t�A{���m���0咲v2a��"�5$3��'@o���q-�-p�~���K���H�����oYqr$P��]dSqD������jK(��c�<;��y�v:�ԫEK�M(��9T��!�^ ����٠�^����aq;:;9��8���hm�ZkaU5���Ӭ����Qgp��EQBra-�U^2���O��ͅX��I_��=��{QӑlR=G;��zj��%������t�A���\.M��j��iD���^��͡@������[�!���+J�Ԥ�4?�nq桙��R���T򬏁�0C��Š�LX�n�u��h�%�9��^���c4��x��P!y�m��U���ºI>2�|	:4���J�h/�C�8kQ��	D+�%��Y#fv� �	Fe�����jy?k�$��լr/<_\��tU�i�!�E�"Ղ(5%�?{**�?���PD8d�`��BTF]�y�)���ɍ�l���]lz�ڂ�Ց.dYj����/a�JW��F�0�fzX��p+��g��뜔p}��I�f��J_U\vs<�)�(Fk1����h�a����{��Z;�+�����-=Jض�([��SNp�`x�n�E�e�z������9	�� ��Z��V|@#����8ar�����@-9�h�F�>n��l�?RKH����(�G�f����K*���t�^���aW$;U��"1���?�^�'��7��'�l�ܰƞ�2��d �k��5[�1��js$d�'�_�K��_��>�A$�G�]���������F�L�/��{q�����qDq��X�d�.-�����b�މ�������% �1���Y�v�>
5hh�6)�݇h�~��ת���~)�$g����x�#8�˻z��%�yds������w���9)�N���X{U�k���T%���j��@�n둺�Jx�!(��p�����^f!7Ը>�N<��I9=���~ޏ4�^�C��&iH,�~���1VRg�����4��hW�C�S�8ߺ�SЭ��D������G����	ĂK(nݲA	�	��	��Gar��EK��G
��$��f����Ā/;0U�^O��~D)�M�-��^�K��#���Q��c��ֈ$���x��s_X`Y��Ĵ5҄gw2��G=ь�^l>U�N�1k%ȕ�q�#�Ů.�1Z������QT����^;6-|�e�rbB��E �Z�x��T00fLU�̜��
�ώl��J�m������*��ĖE.=�Ux�
�!~�j�`�3vD�F����r�q����1�(�D"Q]�n���	Pͤ��<��n��UYOT��A�o؟�_���.�F�aŰ���M�=�^��%v��ɇ�X���{��L�j\OPJ�G����Z��i�<���`���9�j��B����)OU/�ʾ����_�HsAõf�8vc���Cu�h/�m�^)
�
M(w{U�o�Q�k9-b0+����2��h��*)S��c؞]�NQ�!�q�CI��=��]�����<�:�n߰'��<�T$���#&�P�JƾuaƼ^+˿��Γ���jΎqzb��e����|+�EUzV�+`�9z޴y�f�6+N�0%�����+��zC� ��e��>z��Z쒏"ЍF��@��EʄL�~��8s��s�����w�h��P��憃C-P��2�j��FB�|bL��<?�HB�s�K,�b)Jk
 �DZ����K%�z���T�iF��;��ě5���nu���l���f:���8Ԕb<��;T���T�{������w�y�v�}_�<شxǫwUK�źX�Rg�S���:�Hb������큈L?Ý���g�e�qVIbx<�JE�cXޮ34N���+��[_������o �P�Z�8�]��B��@>�o;�De���%�h�ah�5GN��c�j�Y��R��Z�I��yu���>�����@�7*,-�4M	�iƸ�H�����i'[�Sda�
p��VI��{6����d��T I��۟Yv��ܓ讪���ZN�!��������������A8O��Mn��=3��e~e���C����f�YU�9��e�<O���^W�����y�$�B_�I�t4��/���&Q����:$4k�'u֒� ��\w��	���z>��3?8�L���qM��|] c����ג3�L-sD�]�s�(�>���1���I�r���¿��H)�;f���%�ߜ�sU�"����x�&M�1�^���%d�8rr7�z%��e���+�������q�]���w�գ:��rθ1{�|1@O����l_��;{h����VN2�r���i�c��7��v�����*���Ɋ�<�o�
�1�2c΢�N9��vG�묤�<l9��}���6�o>_a��aoTu�{D'8���21w�Z�W�|9�L�9���MSM�&�5��H�S����C��R���؜SA璞�=�8-mm�d�|Ք�����V�+9���֑qZH��4O-�6�<נ��Q�F_�2#:;,��C��Hb�}������,���ifmO�G��D�V�=�{���L��5��x����O,�3ڋ/e��"TI�Kt�ѵ��(d�hf�,a2դ�z�F�/��Xx�?�����і�B����X)�����<ڕ$�9��Έ� R������<�-m����m6z�����P NU��8C�t�u�|P��&A���k�a��Y�ƫ�7�m%��z���&"MA��� ���zVu󶢅C�ɻ��w\a�����s�
	Z�B(�UT��@=�)�Shsnz.��-����>���3�8��Ox�^��;5�J�ڧ�2� �x�>��jh$�i*�2�4�jeTL��!��8c4��_Q�CI����P�A܁\�V��u)�ŵ��=6�D�9�^�wp����+݆�WDʹ�A�(�1*��Eu��M���v�8����hK
�hW�~�(%��,��*Y�4�����G3+��@�M�?<I<��#MԲn�\7�s��x~y�T�H�XQ���{�u��2A��{6i��o�+��p���������T$��en0T.�-Q&w�w�KJ0G:� �"���ս�|��ar�y6�����PQ"�Pi�Pܺl&l��ږ�u�J�tϓ��<��\�1E�$� 
K/���Kҙ�� �a��<���9?����s�uW����<@#9������J�3�l�öeĚ	G:�B�zפ���ك��c�Qi�^±�W8�:�<��<T@���\:ຌ溘�c���ǔ0W����C���@�C��|D�i���1��;��>f�Ի+�9�-�ƠGN��[�QG݄5��g��;�q=�3��"��LZǪ
�ꚝj�iߒ�yy�&��Yγ�|I��{�c�]��p(=�RA0���֙�rv*l��iw��/g�NH�����3����;L��N�c9jc?0K�(�)+��"��z�{s���
�������˷�o�Љkg{�SHLn��\�� �`_!�征&!�ѓ��m��1��]��Ek��+1\��6���A��M{Yޢ,�=�r�g$���җ#�+D{9�$��r��y��o�:7C3T��]t�1���pϦ7~և~N�ѐ�f�#�-�D
�����N ��nh^|�g�[?1����G�ʢN�	}��p���nVB�2�y�̗�jj�:��������N��b�DF����'�M(�+yڠ�Ǆ�uߓG-�
e|reZ$I�6�KF~x?W�[���>�*"���C?�0@��\O��ad����i��4%�_������}Fx��z_��g�/l�J0e5Q��w��k����d��� ��=�O����45�|:�O��Q���&/N��������/�>�'W�g��Hh�?-PLf���"%��~�C�(�����"_�O7-2L�~}1�(�>�@��)�g��U�95�g�]��($���!K�~�T�du4��sI�-�7|%P�m8�0l&^.)|#��-�%��!x�$ö1��t��Xt�j��Fs��Z'��))�F?�S���k�o���zq)����Tć��5�A�-�E �j�#(�f!5na�]b0#&�	'�_3J+�W�ӂG�kB�S�+JC������'>2eHJ0E��2�k#�R,�Q��M$������p{��N�"qnF�c���\8����^��̏���ǥ5j�)a���/��9ZiT[1��D.��j��]� qҨ;ZĎ�|35�v��5`E!�$Ǐ%�O�0ݺ���>���nu�_5�-��d��i����.��p����GT�y�p�U�`�?P������8�����M����&l٥Mq��|��{�x7�E�2��q1��x-ϣM�Rt�e5
߾�%���'����៲tU���v���z�n�~[G
֩�[-l1��@�s�B��)��&MHQ�q4�Ed��<�غ ������}�ۚ���T���7�H�&�i6O�ŧ��¾��� ��m�J�ڎ>�j��_� 9�oZ����h����V�◡= v4���G��4��k����YV�>�eg;s�A`�}Ic3�h�@D��z��S���d+�;����k�a�gDd��k�^�q}x�T�T�*r'�� |��m��Lߡ���S�Y�~���3�[���y��8e��1�_����~XN���~{�8�F+A�>-5Ֆች����"b3�pa^G
�����m5�Tv���Y�?�Ui8�|@D0ϒŧ@I���u�E�~B~%ΆR�y�m�6�z��$$�����o��m�sQ�5"K�gw?�F.,�YcD�H@S�Ϝ��*ՀY8C��m�T��8}��@��y�ъ=RA�dz%��a&0��_�=���̰�K4�
��,,�B� �7z՞�)~I�w��{?O�.�ec������+��׷i�:��Q�9�~���l�&����y�6h.`$p	�xi-f� Ev�����=� �2�0�Cb�c���A�HG������50� Q[�H�).�8�xVB��u�<��&�&xz��b�G\�S��y�{�]�·w��㎵v�K�7���*p����G�)�2\��/�<�!��z�z³w�Ly�k�3PW��B�ҏ�vE}�~W�v]��=�N	W|C�:�p���D�,���wp�۟t�zS�h�R�6�[�̜�t<� �`��{=h���հ<�<�X���e�i�j1���@g+�[-�����̺4k�a�1:���`��Ԭ�$$�
rf��Au����;�J�&5� ���l��}r�Ӥ�$2�G��z�cr[���(�6۶Qfw4J//�#:<���3�e��ņs���]�-�c��.
�i�:���Upv���\hS��=4��uRn��j���D5��c-��l��Xq�V�@������k��93'�`
@�;8,t2��@uu2�jk)�"H������V1��v 	���uI��b�ñ
��%�VAࢲ�0���4��������w�s��Y:�Q��+�9?��On�X��Ӭ�����8���~����/1���pˑV���͛��-f�&��rgC+�w��B�#� XS2"�"��a;�?�[o(�<^��7����6�=���l\ɹ��z2�At��H*��Y�@ʀ��Y��Ǭ8J:�P�:o�o���d�y�8WP��AF�� ���k�a��=�
��ydr�-�	��vMOXF�Ӫo�.�O:�����B�U�������{x!��ZC�x{�o9=�G����o��Y x�h[�m����L�K�+�����f�8XS�l����X_�@y��$�a�-=�X�Xծ�"�f�����*�	4,)�������r3A�ܒr�K�ٺ����c(����Ц!�)����[R���\�_�	� x����deg,z e�����É%�vܡ�ۧM(��Ul�s��R��ɹ��a��1�r�?���TĔq��u�;�t���W�A�?�ߝ�-RQ,��m�围���N��=�wS\	|m'1��d�g����zL=��x27L�S��@���*��mUx�ѹO�+8mI����=|�j�����i�K���C��T�e���F_��z�ۑ��3U%r�![c����:Uݠ���z	`
˂��%,�i���*���.�Ɉ	�m������v9�E%Zg\%�$Ǻ�I�����yu����/lMdm��L��l����,���U��?��Y�,Wfޙg��$���m'Z؅���,��Ӛ������p�1��a �p|\�K )��p�Ո�FR�)2�d�@�������5vDs�����<�3eb(#pߑ+Cq�.���`�?����+uTfq��L��[09�ٱeg
IPbM��W����I���CO�1,�;��L�μ�ap�:(V��|g�<�Q�b�̼u�%ۑB��E7 ��<����q1o�Dr�J�=�W0��v|����0���4��'��3�l>�$u���r�R��v2�� �}�y�}�;j�p�-�B�c�>���x;�tK��1՘%��e�|A{���`��_Rɬb�/ok?,Rʕ�.+Gq�*�z���Ͱ=Q�M�䭔=��v`<��I9���C5�!ާ����3ې�C����ϢS�ӎ�Jp��H����
8���B	/ۼE�ȍ�����L��9�|k��O��#�H7b� ��U�:�߀��G�h����eCBH�&7�\��Ly�Py�����f����lՌ����g$��VN�ܤ�fUE
%�6ٮ�;Zne�u��qL�ѧYںs��=�PU �ƒw����f��ڋĸB��5k���5'����σ�*EГWV]����SH߈Fr�y���Q�HxF�(�Uw��t�7���!VWo<��"�'�p�χҘ�`[��>�-;ږ��BpL��	������^$I���<�e��Z�[L�����.�Ͱ�ϥ�9�4����>/9�'jwpx>��ٕ����́a@� tCr� �2��1s��Ff��m�V�GKZ���
�F���{�W�Zݪ��y��ey3ύ\mZ��<���\���1v�Kv~Xd���YG�56�g3����휚��S��v�Ӛ�1i*���Bќ�NUM�TZ�����eqUI<�WzQ���BiR/�iY�}7�٬��Ns}�ͭs�ZRO��?Ӭ�R�c��ྞ]Sب�xVhθ߀Kgnߛ�|�b6�������r�� �O��H�R�v�p�j(-8�������`�����bb�֝��H
���B��!�)fy�7X�?Y��?�.��և4i�S�*S킍.����������i�������!����%%0�,��;�'���&R��fk֮_�@�PI�Y��� ������}'{����$& �	�Ϩ���@F��î~���+�d�nb�L)]x�A�r�ꅝ���R��𫄄p��~�eRm<"� ��������r+�>co�`%r��	���ԩ5�DT�cT��w��i���n��Ɋz�w�⋸��D{P����w��w��a����hs��!	:R/A������zA���Q�iЗ��}I�R%4�p��fs aY���Dbю�Y*p���g����O)Q~I�D�S(�R����c�`ELY%�u�S��=h�/_G�k~d����"cSw��
O��.���\�qD4A)Ч��[�蜮��	E�l+�
o1x�nrV(��Aq�km���V��O���d"�m�](*�������<�6-4i�1��t4�l�-��S��3��P�G4��� Jh�{�D��]�&&�N�C w��1+�'������g��R|��r�Efa&x�Q����?_ސ v�mN�_nUs�u�҇X�Ծ�; �v$Y�K;�2�w'1�M~+�x�$��A��w��ݬc&݀�;_�n���C�����>YK��$��4F*B��r�|xaNH,e����$Uv(��Wk�G)-wGX��vG��Qg��q�C��Ux���[��8#����r1ͭ!fpfa�w���I���O��$�d=vl;:S)�YH"�e�j�� R��N���c���+o"細�Ga4a_�v�Dk:N��x^����*Z�!������2�wCߤ~_%��'��s�`��
��I'�ȷ࠸Q���%|K=���܆� �ذ���ܘ\&û��6�d��̌�䣊ϻ�O��j�|o���Z��	���j1���jo�"|����<K5�F�H�F(w��ch���c�@����sl)��������rh���_�ט��m���������p�t���Ŭ�㔡Y�6��g���&���~�H�rd
\�
r,^��Q&uMR��M0�b�A��$1�(�uiJ&�m����W6@���z-AH�4i�Ac���H�RB���t�Y��r&w��a��Q<���'�=I��^�[��Z0}���0��H�]��,<��B��F����bY�!\E���w�d[�#߾�-t^��$0��O4{�CX.�s����z·62��K]'L�7`�0K`�0�B$�҇��h{R{:�і�T���&h��wC	wN�P�� ��'i������5����.7-�k�5�h(��ćԟ�FP���ݣ���X7@�����1z;u��$���N�S4SA�U�WG��8�����wԅ��g�ː��H �o8�~�O��k�x��%����Ws(U�5�4�-uHǮ��44����/�p�}l�X�ˁ��/�x�{���Pý����25�	0�{�ɇ�,���x�W������YH2����^b^|��L�u�"6�V��1�����Z�y�"����P�	D��s@�BWX�?ݶIGBxG�Ӹ�iKD>˦<ɩ������ic�������A�D*�'�+��P%�+���R�np�C��
�/p�M��{6}������m��s�*Ii��vC���і`�׾��Y9�]���zSZ����pBU�+k��H�FZ�a��ZN(��VrV(b�37�@Y�$_�:��bp����D"��١Ċ���/t�o�H���~�4E߬�+g�\��Y�<:�E�q�p���CT�ժ\gG�!A�A�J��or��G|�f~�E����������3O��zc���Ù6�;v�&Y9}'N�e������������q�ޓx��3MLL�+��-��n�d"? k@��<C�1���g���V��Dg�gN7r�/��s�jS/;�����?I�fҏ/�_�=��څϒp��͂	 �*����b\�#*�;��:�o�M�b���lv�A",�L_FE5 ����Lb9c �7�_�j��g�=4���o]6�C_K{���q�F���-ys#An7N�X�M��e�]u��f��|Є�De��^z��S�r�p.n�wu?W�� {���C:Ҙ���ϛu@U �R>�+x.}��@�[)3�S��?�q6Ԍ�c�]�����<� �� ��(�]`
��T&���a�,�N�K�%|9�VϥID�P���L�	��t���""^�ى�9�p��P+I.|�;4��
��|� lh�r� ��/��_���x��_c�y�D9$'����A���ϩ^���܁�N���҈�e�Jx���i�2���Km���پ(u�+�y�="{���ʆK̘/��#T�^(�]�����YL��n���{��V�b��/T]hų`$�M�ୟ.�D���&n ��@���מD���H'$k�Co������&��5\n�L:�b���V�ُB��d�M����'�(��
��× ��Y
�dj̙�l�'�es����=}��UA���W����k�;ƒB�yt�Ā�+������q��z,�t�T 0�@�|��-��:��G���ٿOh�����S��A�O����w5$���˘��eU�:U J/4މeB�%�Y��^��	v�,;8ń�8���r��Gg:�K��%��w_������$!�?ɇ�bi ��#1�G�Q���v���q��Ve��4���=�p��m�5����>��b���;}��&AWOc��b^�5���cI�'�������p8�y(Y��Y_�dv��|�Q{B���M�N��n1n𜙢]��]�
N�%7�b��������V�1z���$�^�
��\h�;�<Xc���Q/���n�'��!c��+M�k2l�~��J>�G�#�c���6KȒeb���TcQ��P���)�s�!0��آ�ҏ��D`-x!O���{��=��CH�W&��j�-2�L�!����q��K�)°
�Hz��FD&�͋�%h�}yEm�����!n��6yE��i��DxS���N�*��@����N~q�TʦY�������	Yv� ����\1�X�)&�^��l�-#JJ��EJ�@F��߻��_�U�s�׼YL�i2'����ɎNw.iÜA��D�3��eX�VϘ^6E"I���t�X������GY����h~x�ؿ!á�1�E'�{fIa�'�}�r|��y_5�[(v�8"̪��;LC6�E�y?�mj���'��]�F�NV�3�£�P�j���T�H�q�\rZ������d��=˕�ڭ<�Y��"��hl��kfU}so�=�j7w5�T���q#K�h�:+�� �Mm���er��.��T$�2��E����[�M�P�Rd�Л��YR�����rڣȅ؜�x�}Թ�Snq6��p��7�C���"���|�I��M�Jz��f�L�!��DC���:�W��_��8����h�q�;��XH识����x \�a�C�i�$L��U�g���_�`0�c'�� c��dJ�n�/d�vB�������c���pۖ���8d�?&U~�M�$�ǘ|������H� '��3aN��k���nw�r��Ѐ��i>��1I�j�c7��yE�hӪ#d�/��9���am�x��c�6"�����G��嶪�>�`n�|�dhrǒ�+Ha��d�N�����XR(�v�=�:�tH���<��G9�i[��9�?���>��̩2#�۽�<�E3�V�g���tpFJ*� ��'�I��>�sw3�6��HC.85@��.%�'$e7�}�]0�|��:ʱ���X=.U�	.�9j��9 &G� �;���ɇwfco�г��ϦVas�9���=����;���/�``��l6��һ�NLf�<��gR�������ʷ@������D,BU��ߕ{zp�ނR9`���v	6�,R�n 3`cqh���,E��'}�[���Z��5w�b��°68���G��������E��'!�< y�7lA�r  �j�����,-��!d�Ck7� �'Ǆ��^�n@����F7,)6]�^Z�<$���j�-��͚ȟB�ÍΊ3��3�CO���TS~49�u��OH�x��X`�}��
�y�Է/r$��p�z[����z�Q��nHh-*,t�$P��RX<$V	eJn�F���2�s�{����9L��9N���ﱦ�xg��(.LN��N\��}c�	:�����28����\N!�j�~��M�=��V�C�%�`��O�`����J��H��XË5�5�����`����d������8.�$�����Ǜ�c)��D�8	�~8�|�p��9�����m�����x�����=@?v@K�*-��j�sX��G�#ap6\�YI�=O�6�1�H ��>��f:�4p�P[�r8s�Nv��J4G?��SK�{ BS���(�e��y[��rM<񖱂�{����z����,k�t5�R-�fg�������mC�����KC��s��Í�� DΖ��֐��@0$�߁-S|6S�#�qj��|�;W;�}\?�j����_��}��x�k㶸Ӈ\�Y�a�)��fǭ��<�G�B��#f�w�:%v(���� .f'+
L� u�>3|�O'p�;X�M�+��0�^ִ!�z,#�� 
�"3\�����vl[ݥT]�l8��~�L6���E�ыl��o%tE?,���J���)C�ħVoBT���%��!e}F���/����IsK����h�j}c�7�����R�'�u��B�$��p�)����;�0�����bG��υR/�cn�!��$���Z��iJ�KM:�Lb���p�z]�,j�������L������g+�!5a��5�6.^����H5~Ιqݘ���K ��?�G�e�����@�G�y1�0|: -T�:��k�~8U�*����&p��$�/]�v:v��3�p��x��5���F�#L & �{�e�EQ���,Ry|��3B��M�ӻ>���-����+�i�������?�� �<�7.]�j�Sxf����YC���Pk>���xL�|��H�����L�ōY�Io���qo��q����	o/{����6�?2��N~�5mR�*S��[��*����¢X�X }�tTL�\��U['�@���#���̮��[��~���W����D�dU� ��<�MBサ@	UX��I�G?�(q���J�7��	�k�
���1}4��8u��2�<	�e�8�egH��|���a�a�C�)�`%7��x��3�ժ�jOW�$�by�T~=���0�	�<KcBاM�̲N4�)�v�M��<�:���5u��p�[���J��?b+�.�b�a���!F�� �g�cN��1�e�_75�E�>�.��GuXC�Q9Q��v�g*�.j$����S��R����mi��M��Xb���^�:���l�B���0-�KB��e.[}���Z����%�VC�INH��q\��^�L�t�հ,m�����f�.w�쿏�V��)ѥ�����=�h�܆P(ĉzs@j3�עٸ��Z0�
;(�3�.�6�hP�&�iC�hR����V�dL���Z�01�_��!�%+Je(�p"V�LI%z�_.^�w�H�׀댉D��vu��Sb�4�����7��(�x2��\r�Y�f[�gEPl�6�d3ؑU
SF�@�K��k4Ģjew5$��oM���Yn]�R|�
\a��,Pn�k���<q���1��a��m�̜���3P�̾q�Y�ry��f��'$p/��5t�H��V!�n���ܩ�*8J�j��K����
���-��"��X^1�y�3�'���=��B�;��S�G��{z���5I[ &���b��x��\�MsBX;���h4q]�ۍ�Ox��B�l>��K*gb��y|�C�Y�j�h��=�*Au��]�݈�`���t\�'fy��7V�^e�a���b�W,��
��P����/�
r��4�p��}pз����tf&B�	�Qr�8��rjI=�N�+��)��o
�k<c\�����}�g/<\����`+t�O7��4Ab;�_%}�O���Y�h٪q��� /ݹ[+�r'���C��t쇽�b���X=�Q�H���l��˾g!�����G�m1�4E��a��^P�J��oY��`�7�%l���hx	��	c���BR3[��V���䲦���7f��[���&�e9�����3MrƘ�J���=6a�?��������Y�.ת������Y�>įj,�/��?��z�����|8�dIos�~�<?���}?QCۭϩ]�=��@�:ùV����9.���jM��RI��)�uX�9Zh�e�0��Z)=Q��P��i��I3-�=K �)K���o��<de΁�ѧDT���r�p\��@\r��z����l�D�>DǑ�#� v01��4G���cU�����We�BUrJ�g���j�~F����z]I�N�ЯӲ)yԫD�
�̢w��Tߑ�w��BI��)F�kWH��S����>m��b;X��Q{7�����[�-����@�]�kwȲ�~�wX2x`�G�'�Z#mCK�$���
��/���1�@�x�g$�n/��� �jm%7�����9�!�NoR���YhϿ�o���_��u�~��gV�n/hH�<���
P1QWOc�b>	a��S����?�R{�����[l��/�P	��ܲ��V�U�w	k��ʹWX��%vSM���*rf?
�WZ�q����{c���=G���7�i��s��i*[|h���O-
����P��..��:�d��g���R�תQ��O�c���9�_@O�J	j+Z$!�z~��c��zG��}�hi=9uĞ���Q���7���C�$:�ɮ�D�f� �J�u���el���;X�9<��t�@�����(�e������I��F��R-��|.�g�1^׃@_" 8(ʊΡ���g�Do�F�& ��(����~a�*z�����Ի]�m�m}jV��o�|�б��|�+�k�-:�(��8��6}B�� �%H
T#�����DQH�@}w�Q���E�l/QO�'�,�l<x��X��RK�.�xJ�����DH!g�ՕJ����xPǔ�L��o��z�Q!�*S�_���nj�B�'g7���Q(���aA��&�Z�.DF���>�/���s���y��Smp�h=�N��0����ә<R�<�^�>�51w�����~�f���{�{�+'��cУ�����9�4ߑu!Z��vS�m�� �W�$D����ގ2�Hs	���,c��Nl�l�@���u��K�hW�L�U�a�H��4"E�x��	��(E*�����b�ŉ�����5^4<!Pz�1n'�Q��ϐ�6�T�ؼ��S�g\��( )��[��0.�@��J�����.u��*[��1b���Y��UWܷM(e츮q�D��WwZ�E%�j�׌6��F���e}-��k����w��S�
�+w ��\c``����P*�V򼛳�`��Z��jxT��i��bhrd!f�21�d�GX
���5�B�aX��ܱwa7�ʞ��Z_��3�����
"��-j:G��U�o8Nc+���VH:�,1�co'<$ �Ar���d��m�Tӎ�$�E���d�F|{}&.?c�T��<R�t�C�I��=7��׬:ۨ5
�(ȫ.�}��LqP�G�����.���?Fؕ_.�(�JH��&�9���ͽ�>� �r�Эܾ��f�=Sy��(��y���d�!}�u�4~�*9]�ʜ��	-
��7Y�򷳑DNgt�{R⼑���E>�{�)��ؗF��]��}� år��	�<ќ���j��m-��䒯�|�!0�-���Ar�4�rB�}�0��lC��'�9#U���Fν�Sn��I�o!!-�Q@�����۟��&W����VX��:��	m�U
|���M!�ƺ���"�����wQ�00�}��0b)�k�t :!�J򣛃)10ME��k��9�%��=e�K�w��9��n�h֊��]z�d*Z�K9`H*}��-�(��e����>��ז�LzI·�K����=PT!I�Ԝ���*�c�u��O�0�:Zf�v����,C�0�L5�L6D0�茗"�dM��$8������8���ȳ�FѓkIJ'����F��;?���o���:vKF����Ad�����P�h��#~�Y�q8z�.wE��YN�I���P�C4[�` ��_�1��d�/�	�v�@V�؝��P���F^���⏹g	H)[�^�H�S��z�e,oY.#;��F,��|rK)���p��R ��S�Cp2�M���� V���a(;w����=�`����z�Hj��A ���:�|��y��[��C�w&Ơr�Ҟ�
�8[�D�㯄k�� ;z2�?0�F�\����|S"<�X�J.l����R+�W����®vp{F������u��`�%��]��ld&z�̒J��Ӫ(
#;ϫv�%�G��^��r��
�L�6�ų��X� o�6����@3�X�����?�+�O�y[����KH)Ɲ+�����	�i|<���YClC��\�D�����Z[��%\ѸqS.}|~�&��ռE��P���W��-^z�(f1/�׺���k��y)�ҍ����^��6(��@��~�qq��>�1`q+��v���A�?<ơ�L@�Nn���a�����*�O��w(��$���sS�⪶jto����`�τ���ǒ�4�i��\��_���V��j��'k����M���cát�McLB�6!?y	r�э��#�|�
��>h(�:���ym�CKi��~��o5��������2}3�^Z����#a8�I^��6�<�� n�7���Ͻ���]�m�:C��DӾ�oБ��#�&-�[��̼�8�|�߶SHR��m�F�����S�����G{�6t� ���E�R�{n�ߍv;�< d��,E�y��!<&|����Qd�1���3�6���+��2�n�z՛�I�;�����o�;j����|4��cv�<�&g��n�0�G��Ɯ^�!
��A��`c-�\�G���[��&��vs,��Wyd!�4���,$��u������^R=pB�L��7�=�"��mJ����p�V��}�:X�3�:.5��i���]�\�~;��<=�XЕ�6(�1O���I햗>�p�$��[���o�-�+.�*���J��FK��o~��l�J������͛��؂ƯĻ;^��qÈ�#OB}l����]b+R�p����J%���Mm8c��'T�v�:��2BEl}w)z� �:~<���Y,���2Mx��$��Nh@!��9�M4��lDd�l5�������bz�W[�Z-P�1��0v ���b8��#��C�x�����#^��a*��d��������3}E��2/O��C3��xkAž1��#����v��Y�:�F�xr���32o�P�/���hU�$�k�3�u\�[�:Q�/ꚕ���^vnký�}����Σ���Su�`�;/�'6ţ+��,=�L��+�\fdIA���H�ww+��)�$e%vrr��=aV����`(d�6�=�x���Ks�
�nZL*�m���������!F�T�K@G�����!�r�����)l*��t�����@� 䘿F2/K"'O������q��}�v�e�7d���(	=Cġj�m5�:�"�}�In�sg��&S_R)6EṔ\a�-��%n��C�Ɓݱ������/�$�7�73�\�g�4�Ijed 0�ɳ�Wy;�U*d_�_��fJ�
t�Gۉ �J:-���U��"��e쭦��|(�)��s䛿r8!HpIB�CN��N�t&F��`�����1�w��,�P�s�d��~ަ�b]}���$�Gh�%E��>`�b�J�Cd"�w�w&�Mbx��0i�w�<�Pkm��}�"H	]��������^@������.���	�nY��p��Ǻ>�z`���:o͞ef��z�`��%�z�p,NT����_���}W�P�P�#��1:4)��f�����~0*���eh�9h-����?YX���F9���e�i,`�ψY�}��$F}�ڷ��\UE��DS����uQ\P�z����-�ZaS��O�zغ�����N�Nf��\�P�<z��s���F[�ZA:(��%0�n��axe��"'a�5�,����J��+�As�V���\V�H��f\�/E�� c�1���A!�PtҖ>���h�}�(݌0�qt ��WQi��"r�G���ő��M1����.�`�a>ܻד�Ӗ\��<P���)M�Vd��	a�o~�M���a��l-'�i�_,�{�R�kZ�q)�}Q�4�ڞ��?��;�{�GJYU#�-���V�[S�1���,���^+�X��^�{� K������c_n{C+q��K������$�
�>��A3ߐy����_�|@�!��c�ð��be�ndt���.y�އ����f�e�����=�ϐ�5@~t�/��?b�l���0����(	�dI�����}NK�4>�r^i��#��wCF���z�2>n2k3�e�]Q����(�2�}���<+yv��s-G����|U}���-��������L�7��k}S��Vt�"��V��ڢP٠ԬH/g�Z����r�M�m�M��Oz��4%�S���U��۳o2�/�����&?���iP��E9�YH��;�X���9T��ð[����"ŭQ��b�۽����C.8����MI���'��S�֪{���J����i���~C��U���u��rC����� �F��7�+�j�~�������_�JF��a��މc�����Z�y*E���u'�l�R?��jS�I��F���X.D��tj(�<Q��MR�����dPQ�`C�h~[��T��Έ��`�8'<�ŧ��> ����0t/�~<�~��Q���@y��Us��E��q*�l���&}�ď�@ J#>8�M8+�;����?�UX��j�-�����x��`\� T��iן7��٢����k��Kr;��1ZVFp'��{���EdzT�툝@_{��q� N��ɭ�-؜5'V1�yʌ@Z$r�@O��_�s���1W��09§���Yz���q����/�Ug��t���w�w�x��<�cfH^ԓ��ANYj^�PE����g �f#�r��_���lc�%5�%��c�X^B����f;ږ�ԤvO�>1�w�'F��/����"imqtU��l�Q�e�#/Y�j��鸾(@U���`�H�24,�!U3X��� j�o�>yS]~�. �n�j �;�M�*+i�.󮭋1U�I��B2�w�H�������!���TO��ީ����o�5�X���޼��u���_g���=M�7����>���׿[��M��;�㢛������R��r�qA�7�	�P�\c8�  K����,Ͱ�aT�W7�CfId`(�^z o�-��0/��k+�V&��	r˄�X3�|�n��#c�.��1�|�����NW�'�
��Y��6��U�@�����%��{�g]����NM�3������D�8OV����.U�'�F�M�g�tR��/\U�|zcm˷��R�Nm��f�Y,�Y23	���L��-l��%��x����A5
��\�^(c4p&�)�>޽
�B��!6 ��Ϸ��A�]
��p����*��e��Ǒ�i�U��3��� t�!m��l�+2���#ȏ� r:�|��/�m�,�:�ڋ�:vV,*h3-��OK�΀|�l1��d=�����[�$�Fl�5k�����Ԏ�����K�����9�,ת/���51v�7Q���������ӽ~��i��[IC�����B�Ԅ�2���F�X�8��e�v3~R�(�����MJ̈́�n���G�y�w�_
�h�_�ia��:�w�����Ļƌ���Yl;����ne����5�%���4:|��I�!¢�,�hi�߿Xb$c`�t{��R�<��<�/�]���f�Tυ=���/9P,^{���"s��[�y��#�b_t�����n4��""�U���C
��A@�cM����9�ysN�5�'�IS��G�|���?�7>Ǽ��aBzc	��Z`Z=�}�H��S�����w��<���J@B|/�؅�:���Ә���>=5筺�$*hw�����P�F�ڱZEE|"��
>�����AC�z<G[��Elɇ?Ww�A�_ŴVlߔx@�����[�`��gԝ-6AW3Ƨ,�,#c��h;��^���������kx��fo��i�FoV!MZ.�/z����O�� ��YDQ
���צ1��V~}��{0�A�����+J��^�g��N�����+��<�6�S�W�@��(f�͢A���B�l��%L��m5��JJ�:���4�O��ׁh�m��Teʛ�R���M	�ߠ�I<6�(\o&��J�o{���<�gGW1A���س���a���?W>��s��z�ZV��0�U����.uJ��u���U����5�w^̰.DX��{,a��˄D��H��r(�h���Q����0ܖ�0tygJ/�g�M%m|���<�����a6j��n^BGK9���M�F���yG���Ub)��R���Z���X8�F')P}�N�
f�X���&�G��^�[�������x!��{�N�fXctr;�9�?mFg����<P��+��9�̇[��Լ'dTO�3� �ר�?&H�`yuc:o죰?O��x��vb�>�\�݄��X�^�F��58鵅���"U�n'�'�|��{�,Q!���4���b�[x���7��κQpQ�v��1
�&SD�h�z�������Qư7�D�rPf�&�{X5�K���w��l�m�F#�����<`0�j��I��Q$��`��f̚~� ]"(��FQ���T�v�?&����z�5���h�M�T�΋g`��Y3�e�$H�M�1��Y�o)�<m>r\+����3`PJzx,4�йVZG�ep ����"�8r�o�`����M��zhL'���H���	�q� "��{��X�+HY^�iK�"Li���JWL3w�!2Bi)ș��������ӴQ����iR�� �9�b&�&��l�<�|���GR5���wj��d��*������:�층�R_��dEږ��ϝs�w'r��dV�c�˼,^}b)r����9��2�L7���a�8Є�<���[��-��󭄥��*�̮�_�UAY�f��.<N�x-�,�R�ռ��VY��D~.�^Uṽj.�ˣ~�͹��w���OB2)�{dh�y���QU�t������;��8?�0!.|g>	iJ"�u}�L��մ{���NS�d2�v/���$Yw*Yj�_��,��Д^�E-�*D�6�b�2[I�7 d)�]�"\O[�T��iO�����	�
;�tƓ��t��z뤀�����\�u1t���DL��/���O�8�q�k��#�+���a��l�q�v�7��Wy�Tj�q�}�D2�hH�r}Hmej~=�6�q/�u.TAw�B��Ǎ���Q��p����,c}�x�fZ���L�iȭv�e�ۨ�/د1%��h������ylk����A�Eo�fVL�BY�J3R�ʆG{=A-w�,W�-���3j�y<������c�g�Nx������h
�Ԭ��y8�z��r�$������N��`[0Ţ����M02^uY�+�]P]�*�� �E]z�j�w���/df��:Gt�agZΝj�Em�?��uj�G�45��Nze׵��Hn��۟ʁ��Z�Nr_��84[	R���N�4U�G+�H����!}=�_O�r���(:� 
&�*&��H"������ǡ"����/���4+D��=�����
����w��T(�r:f�y\{Œ-������~	~�)#-�B
:����m��#���!)��+H���!�S�JN�&��f�|��3A"�I��߉$��O�_ph����>�p�w�:bS�Ј�.�� ��F�`m��m�rn�kܚ͕� �����[;�{�"d���{��5n�C�KhW�H}V5��KdH�e�Z+�Df;2���H����m�����eF:nt���i֎�
]TɁ:�S��e���7q����\�����e����5�	�㛥����Y(�ؠ
��xP����@��S/��h�0��_]��ي�=����b�\A�����&e=]����9�����Ƭg����+Ύ�?o:�]��Tt�gV{�;�/����g��*	��i�h!����>�s���E�(�S����B��;��g[��P��۱�4�7,�u`q������Z`�v�ӫ˛����f�z����iY.O���<|ʙ��ǆ#KDv�%�ʜ|�  �|��_�a�\G%R�y�'��ק(9��Lӽ�V����\�h%na�����
�,lk��l`d�/�p�.�w��g!����ߣ�mY�G㚏<$���!8��?	a0�M}��d�cϋl�b�[i�����
(+M��uf��!X�D���n'��VLop
�˧��v��v��}q��x�o<1F������״gӆn����4�Dw��v�x��-^�r��1L��ʢ)�3z�w(��$?��ј�QgeNm������N���>�H�Z-ζ��+Td�x=+۾�����yz5��a�wW������O~��Z�%�}O�
���f���r>�
\��0���\QV�8$f�th�W*��Օ��m���TZ�A�6Gg�:��L��S��<��i���(=���^$S�W���� ��C>�h1�PTͷ~��
X/�ܹ�8X��YK��fQ���.����)Ai�EQ�[I�.F˴<�D�#/���3DF�+�	��u��J�cFP�/ZD���X�����D^�V�H+ߓ��.��a��vʼ[��ܸAŭDN2�=e=r�X}-Õ���;Tq�3D��'odͮ�wPa� >���'B3�����(&��e��~e�gu��ΨZU��� ��s�'x>�o:��C���h��)�\TC�����,v�=�#�"���g��70\W.�l_%Og�����F���EK.}�\O�d�U��&W٠��[GO� �i{��D��>��p|�C�p��Q	x ���)x��a�3���b��R�
ڲ~Б� S��$;e!������Y	���}C�>����HQH��) Q������"[#Ϊ��$2z����Mw������x���O�Oi�m��
�ëR� T\:�	���H�`.��H�-ŀH(�6/â0�Z��-�6(={j�.~"����u �;���x����&�4�h����降�ȭ3w��;��Ni2D0FU�	
�F� �t�F��7f�3hʞ�| N�\�ӎ-{�����*s?�L{~����Kt�Ͱ5<H�}�����;0�{�Ω1e	�y��w7;f�Z��=zt�~�ad$P
B�ܕ~ j�93�Ѩi����64L��kJ����(*8 Z�	{�b�:�]u�@0z���7����*M����F�L�h�!��_ϝ���"�#[H���z��[�W?<�q*63@hr�ki�z1��
���j`��0=[�4���B�LP� �F���]66�=�~i��z;��Bñ������u�聒+P؂�r&�:�����qd'�iM�_z�-)�F�;���}�Ҕ�����*tP�A~�8e�]H+����h�^T�����X��x�}�ʢ;zA/�Bg�C7���ϺL����r�=_JM[XH{��V�j4����	# �A��b�[��t���u��;�oMn!�
�3��WX2-��H5�Il���	_�M�!��<�!7��~�ڒb{�e'���a���kM"g�L[%j��/彤��	dª^řoX�]��XOs�K���S���1VY�@{Xh>01xXVG��B�:��>,����_di\>M�0�`n>@6�f�a�4��E0�DRk&M���p��ȡ������R�u܌*e�Y"��2e�8��c3�fd/��Kt����fEdpR�SI.�$*Px����h죶���ϩ><��a��J�.2p���30�Lv)&G(�=!	�	2j>B��L�w�1j�T%�Y"�:p�A~��Ӊ�����-�n'�fUA߭U��td~�b���)(C�Y3V2��)$ɍ���T0���i关k1��>ʢ��_�$4}�g.����cx�4�mW��L�����7�������κ ��4��z#g�v�.���|�D���,�.zK'���c΋IB���)��.��XP��=�+�h�zҞ�m��pϏ�"�䣭�Ɽ�>�ln�_,�D3��^�F薲�_�@�ŝ�h�uN􎅇P�]ԳD��%зdx!��b�!p�暖��~����Rx�WlE���C��l�J=�լ���0[��2LJ����DA)K��������.W7G�qlS�YMk/$"����#I���tH���)�;���l���5'�����n�K� L�d[N�k1d� /�(c κ�Jc����9S�>j>.�ng�����������Y
Q[�-������
ߦC9�O��(u�tJP=�4d�,��:�TD�WZG�&}�	2��m����ԗ;��8���`�A��~HP����+�ӕ�n�P7pi���q��[~Q/�R�b[��<A���$8������HiQ���,8V��(6���`34vHLP5���`�@�^H��@QA�7���w��8�0\��O���|^=����*qMs�p�MzثE��V��D�X�u~�\b�+�Ub�Ѧ����д��K��������~/��"
���!��Y���������e`��+�3��p�I������	�S��|	)�KW�oA����m��}gtO��.A9f�Z�E����F��^n��\��Ms��ƛ���x�ϼ������̟*��қR^vN�nR��=K#Yө�
Ht�QE��K�i�ˮ�Q���Dy�y��
�N�N ��g(�#73Y��Wإbc}��s��G���ϸR�sࣘ�o3^��!�B��8��$��c?4���2:��#h�\�9����J����$�s���c0"��T�~���1j�	�[|�X�����%˅�� )��2ڰ�7��0����c���K��l���b�c����++�g��Q�V��s_��Q��F����J�;V�=�W<��y9��[r������E~�v~$�,�6&�_�|sLƭ�LXh����\�Lw:R��H�@V�8\�QR_���h�$�{�ٶE��O�:��LE�Z����3Z���rk)���	��SQD��ݮ�^N#�-ϸ�$�ޓS@����3�0V%O��غE~���$q���>�	��*wi<�Gt�aX��V�dS��V�o��6 ���Tmg��U�QQ
1I�K�d�9P,#��5�n _|ۡ�KBI �Pgo�1�l�VS�r��t->
ϗJ�i����L�B�n3%���u8�lD��R�;-���8_��	[�&4���H�)7g P�-)w�Lф�8L۽�j.nRO��6]�i̷����B<��9��ESIZ�;x��׍��OdcWC��M�$�͖M/E1ʣ#s�"�`v��[���?ְ� �2#V�b�����~��y����4���<����_HS�'�MC4�C����P�v��4��s���4�җnx;�0��.��@�-L�,����Q�ҷ�2d��)/�w��[Q����@����]��:m���}NM\�,n���y�L6��	,�(����i�A
�]M���H�#4B�����&�K�'�N���hV���R�n��m�4�����j�~��نn��kQQN�q;$��
�1����>7�ӯ+�����7����Y��3Th���]9�y��d�7���� جc3y����C�xX�s�L9r~���}�k�Z>Y@�+��`�X��F����b#h�i�1�R�vIO ��)RT�<m3�e�h-�6^�'���剽��3\;z�n��o����Դ���+��]��x�m�G���L\-�������� �x��� �禪F�j׶��LY5.D�K\����m��*��&슠/f���w���,2����O��cb���cs�c�ܶy�ɱ�n�� �TZM��ү�����h���`Ҽ�W���q3{M%�1�l�\OQA2+_���6��1�=�n�&@�_��zc� �~�i�~���p�˞;a�X�p�	�$F��,�S0��ʎ���jy�Y�ìܞ�(�}�Ò�ȩг���G֔�r|��U#n���V��(��Pl����zU@G�p��Of��u�Ջ����bЮ�"�Y������ҵ_*�T���(­L�Jw�C����sq��ϫ��q��DVP+��Ę���e�����<Q9a0ՈT�,�PQvs[��S\YEp:I�R��(�O�t)|g��|T���	�����9��2/�����P���@�̳ٞ�����[Y�J�����ء�~+b�-୹�7 <�)��H�IŲ������6�,X��EV�z<�5|/�Z�I2���A��<���J�k�eT��������=c	�x�sD��I7Q'��-�{��|
�6��J����<N�%�����n����������l	V�������$�h�Sǜ��qB6�@S��G�+��Q|�Wgd��7)�k��f,���X�l�H���� ځ��c��c�"�#{��;t&�tX���/׈+s��r^~P������#���8�BFe��EW�/=����Z�k�)�{���UAA�G|�W��q����VS6�����0�j廚xH.��,���H�I؏��Ʌ����/΀�nQ���di_�u�شˉ����]��Ti@P��� �(u�����T�5�R$<q�h��W~Z�6o&Wl�r#�>��%��`:80�C3&������iN�%�,���C�ڈ��T���	jgۜ�,R������G*\6�z��02*sJ���TH�f��(-��&�: :����������nÒ�)@�$�(�����ݩ��=Z��a6�k�% _���}�0��Hd��ԅ=`ҪA����� i�4��M#�R@r^:}�/�ƥdp|r�,�-c�����c�W��3� rx��q�w����~+�2�; ��>��gX"B;4� ,���3o������b{�)md� kB�����J~C�S�Ԡ|'� Ru���2�E�ܴ�6��/��0��°���1zKG�� %��U�ǝ]�A_P������殸r���5 ƨ�>M��[⸰#*���B%��<��Ⱦ�_D/��6j�P�L��].1^�Yv��7&�3��Y�'{�n� E��n�R�#��j������<9Yс����t�@�byA
b������Y�~�?��ko��t����}*�{zu����C�۷/�&����KWu��":B�[H�L,/x���S�5��zZ_J�p�Au�خ"]VP.�n�֐��&���)RO�e(Ds ���~��Mxw�r�G�F~ݞ�̥]%��d���o�Cw}����!�!��(��H+M^����н�q�����2S!݃�%8�-�F�?�U��!�1��g-�r��92En�V\���=���O���G�Ј�1N�������|_y������`�;�UZc����]}@H��#f̕�O�tF�%1E�ذ�,�g���l��J"��!G�^No��	�v$�LD�}/]!�Ip����m�'rT�$!���#gV���]ͧ���Ѫ�I���{����ʍMY�L� �W�c
O�V;0��<E�����WOF�d�)uN*\ٞČ(>�%眜
��E���ł�J�'�U� ����qx��th\�g��ь'd
ܝ�Q������Q���	&{�RQ�O�Qz��ټ�b����\�3�n�Y�'Jǳ�*2��^�UV�Z��]�C�GiX��D7�BҾL&��Ow��\D켶|��*�bn(�X�;�n�>�AtJ�Ogڭ�*c�C���['`gz����z#�j�ގlY�AN���7Ȱ�%@՛zoy3��W��@�Sϕ��u4�iJ�e߻�j�>揵��6��!���~�-��B�*�R�`��9����ȗ����|��[�)=�o��}�������(?��7W� v}�Qq�_��������Uɨ�o�W�&���K�g����(x��X��R��vB�s������0'�d�#���F��)Mh�QE5I��y�/�;��Q��� :�+~�������D�O�<����z�C�R�����,]�Ϸac9	��d��^{��+��u���3<���+�ǥ,0�04������+q�tFR��K	��5Z�0��jo<W̸7�/����ʕƢ�P[��
�o�iuCu�k{K���q
:x�S����F���oS��x%H��}�K�8�P��nX�t���n(�Ĉ�D���]"gij�\��,E=W�Ԛ�e��+D�x��M؟�~�q�� �w��m�Mv':T=�;%?C �[�2lh��Z���`d��|�qq|�Q	.��j��i�l�#w+^A�]�5x�]?$MM�M��&��g!�O����ީ>��w2��"�2g_(GoAw���b�WQ�q�u(�.��%��M� f�fc�8˴����.�ǿJ8�3�΅��=T����Et%�=e� xmT����B֓�`%�* �lA�QNo��ב���1�7���<L���c��V�}���P��	��󚅌��#��x�p&��!ѐ謂hꎯi� ��\�L �* ���<.�vmY$�Z��j X+d`����1|��ڈ������p�u�b��72������]ӥ�	���
i�����f���w�o�}�!5W��k���M�tX��d�3�t3pU������h���w�I��[hA���+?P����+��v	��_��o�>La�O�����"��i�u0�#ۊ<�H06�|4} �sMʳ9J,Xt6 !4&Z��rb t�r�����{�Ѯ=c��o��J+=P->>9��Q��4N�(�׽�4���>_�>���V�{���e�؍�7�fP���Tʮ{ N�Y���>�Y�#��4����wi���d��ƍ<�S�rfxEe�t�[�����a���PY.�6p""AW�HM� �~qG�#�,!�t���Ғ�[�(ӺqW!t
&�п�/���}�a4g�ir'�������U��NI�(�ɲ֩aj��gI����/pl�<*����S��g�:�Ν:T&M�H�"H��<B�G{J#��.��o��uDЪ��T|�!sU-xWj���7��L����{���Ӷ� �OnЌ�>�У�WPϥ|D!5���%oK	D[�~��Գ�f-�ֻma��kֈT�}�ֵUFz��d��20^�z
�,3��vϥ=�rG{�g��kB��$�����l���"�ڽuKD��뼂�oJH�G�فW�j{�OarRb~ ��>� ���\�?�������է������<l1dbږ�D�]AW�}���Fg�
z ��� 	n$ ��؎ʣU��j1K��ޖ�o
!�齚S��ܭ�P����]��b�|0�)�n X��Ϥo+"(y&|��B������2j_�Cn�}0�L9��a� &%�zaN�_ۛ?�S�!���9�+% �&����=i4	�]~�آ� %?��4j� �g�������MΖ�q�������)`2�􂠦��	�4ќ�1����r���G����W9��+#����4��o�I��]KWw�t�@�Rᖓ�@>�uBJ�$�&!�P�7H)s@�-�'-�;qïFn��,�+��e� �u�tUA��}�y��/�'ַ|���l:��:,�_�O�� ,˛R|[)��)Bm+�wi�/�@��F�W�e��aYrV��cٸB��8T!�!k�r���E��9�Х�W[����P�H8����o_����E+��M��-��:�ܜ���XS��}���,ޚ�۷@T,��#�|oI3g>�$��A��9 V~���Fq}���f���y��ʛ)@d�x�(�i?�N�g��)�Ę;L��H��b�{�4"?���o_��;y��U%����+�S�|u��GTlol9��/r<2��hU�A�nb�y��x��=*Y�$��U�� m�[s[��O�&���T���L�iR��/q�E<�^�}�H���JD��/.`� 0)XT�8�	���eB��F�<�'*R#��2�����e��[�׮�Z�?ꌇq�"]Du܈���Dr�-X*�xݎ�/Z��5_�S�7:��:�~�dK;Ѷ�1N���K�������$Ԍm.r��[uao�b_��*Y�R���\��C�<l��:/�z���Ѽ��2���֊����5P�۪��?*��cѲ���0�fW�<TMt����n˯A�b�W���$�&�x�u���l�fa��ݼr���zЏ�V��_��}�tT��  9`t��1þ��d��=����q���:G_ks���L�&#<��H�?i&�$�����<���?��rJ�o��Kg�_��Jte]Y��쮍t��&Ԩ����T����G�1I�D:d�w�y*��� ��QJ�#M��4O�|�h0�#�5����'`D�r�Zj��M;�Oa?"2;�F�~� *�s��wE,������$H!�N7;��������J�v/�N�m�GQ������{O=�xy"C]��o�#���\���j6���SMc����Zl��xǳt�!R��M�2-=���m�B3iAwDS�W.R���������#�����w��؜�J�*���̒
]�c6�]l�X�'��}��n�G�$#�<1%ZEB"Bǵ
�"uʎ�X�XT$��E&�ڽ��'G:���N��m�L+�z����7��n�����*�t=��)�Ōv�lIX�!)�;YiD^��xb�k�^19e���c�;O�_�ؼ��ؓ���+ل�������������?��5���誇�=�mYr`֤yW�8]�J�D���Zq
]���T�I{V���î!���q�̸���ս�[�u�|q�^̀)ԒN^�s�q��P�U����L� O�����`���S�hUSd��T>�nSuǎV�8z�6
ǬO;��0ft����%�Y�u\ͽ鄅Bi�&3�������,��,�z*_��i��ޜQ��ꀤ�ތ���j$��*���F���򈽝ى��Rd\Ǒ�'Xw溭YK�.k��Gke#�7�ID��2�R!j���V��@$0h���]�6�i�v�Z�L�t5Iֲ�ۑPF!NB��*����}�!�1�V_��x�!X�������Uv<y��ˌ4x�̦�t&����uM�V�"�<RJA2ai_L+�a}x@_J]�XYV��"A0 V��`b��7�b/��Sh�吲� g��b�zbH'��.ώ{e�0�`Eȩ�d�2CC�	!�e!�]���	�B�l��L%��4RO����57�o�Me�65hB�.fLk�hl��.��|WǾ�s��5N�d}�]Qk�Q�K>|J@��q��zmu@Uf���҇e����AW�M�M��`����6��I��k�]�/hh����J���[~p�["�bE��9i�8�M�����p�{b�(o�C�m�#lCYs6r�8���B˝Ae��/���hM�3k+_Nre�h<w@�����T8�鮫t�[z$�b?��6R&���VI�QX˺Ʀ'�S�j���c�j�դV��� �kn���@t�<6�h^+L��g�m�#U-��l��	DD*�Gl$���>�Vںiu�}I3}��AI�x�cD�6!�A�^�HzFx��d�Gj�aw�V�Z;/C�Q>�m]����0|<�cc�#������م��">{c"��8?մ�~A#blM$:nmZ�^�;�K*ɋ�w�*C-�>r��
�t"��h���!E���@ܴ��k7�֔�G��x����a��j@I���.t�UK^`N�T�~+ͧ=���Z�z�C�����k��71��I=P:�Ȣ�vU�_X��_���v��'J�N�,�xE��} ��#*}C��NoR�W"�4t�Y �:����O�Ğ'u���k�~��͟GR
�|�G8�\b��Z d��b9���9:T��(�&��<�$3] DݻJ�8mdn��evP0�GY�ٝ��+An9%&�+�Y�>��I���[��UJ=vfO��i�͌����E�mbcM�qx�d�����w�v�"$�����$z�FBڿ�x�T+_���%MD�i'�#�BCJ��4�g��#�y�H��7Z�ѳ5�C4d}��};y�8������zF�F��V�z}�j��$�h5�MJ:��_�J˜�q;���#��ކ�JhP��Y��jW���C��E�_J���<`ق�1�b!��.~m��<�Q���86iP��0�a����X2����(�N����*4�$s�ƭ��{����V�8\�qj�fPA��|U��ct	ux����$���-���-�3�qv�[��tD|_���!i_�"͋�;��n3�0OI�$Ez�N�^�,���nFm.�O3��]y��鴉��5�`��~b%���h~"�_JD��,�XH#M
��Ͱ�v��<V��6�B[iT�4�YM��+ҭ<��p�,�5w����́g��U<���ܾ��U��8�����AO�\�y:�=���y] q�!���I̎=L�>�1�?�����ѩ��W.�WX��c�����7��#�� � r$$+�׏��zCk�FX�5��׏= W�q�H��?�k֜o�a�x~�n1�vWf����t�iԸK��\�������- &�'�A�9����Sӆ��:�t{�����Ů�GB�&���qh)u����:"��:��ˡ���v��9�����=�-*�&|#}���r��o���rT�N\���E@g����Sz=@��7��ߍ|����Gx$o�P.��EoeX��5�S�n	���̨T��k$��"b���LDG����[=y
rV[`
��T�r���M4uD[�7��5Y��^�ˬa ���^��<�D�y��@���A^衂��&�0�:P")ìQf�i�~��@آb�Qr����~d��U��x{�ay �PΈ$���hW�u���"���4�����S��l�e�k�`+�.��}�G�AFW5�V�(mR��6}�/���y;j̓r�
����ۍ&���	���ʹ{Q���R�')d�� M��h�A�H��4F�	H���L�`��� 
�-����MQ���S�jZ˲���#$�@{D��	��aI)�8��{M�NP'�,U�i�-`���n�7]��gq�=�2W�
,UK'rl���O����(�Ɛ����+�v��.u��v�W�zB�S�.��U&��@˶V�`��޾����}n��G�E�9%����a���xw��T0�H���מZ�o���S��>L.�Z��Z��(r���K��5�2JSnL:wx�������&�r��U��(�xI(V��+)�i#�"����r��¶��+��b?&bEU���bu�M�_�������TV晀���5*E�>4^������)�g 0S�8�j���!8E||�tqq$'#Md��Y�3/����bL|��_�W�l�)ʦ0:j�\ȶ����y`�}�m���b�"����V��[����ׅ��I�=��}���#i�c"�>B��n>�vx"�����m�g��|j~�OһtX��R��2e�@�d�C����uw��4!�rcI2ޣ$rl�HQ�� 6�����Z�hO6*]���+Zˉ�}H���B�� �#��V����"d�K�����)o&�[��fy�7m���?s�CT�(l�����Ra	HZ0����"fJbGl<��0�G��݊x-ά��£0 �A�4�QI�����5I>M$xm��pv�����dµy��=uf�V��s�[%vV�z��^ҁ�$H`�;q�$Z���'m����J��b�0Ls{��~l<��cTK�	u
��?Fں^6�W%�+Lx �gK�9e{�y������@�Ι@C!?�sm��4�)8���~3c��$���s���.UUM�̓���9��D,��;$2�q*�F��m��SQ9�;�S"�[�
��Nt�ZK@���o�{���`��O
ֲ�����y���˔��0_�1�3�d�����g��2%/�6SU''��|�&<��]\*�=��Ѳa�(&�:��F׵��V����`�b�[݅\�V���0�'��ug��ណ�Fv��lxBA�7�"�ݼ�Z45�B2qfF¾�,f^@!���<lv�������;�$�Y�'�AJ��o���7�t��� �"Qs)�k�m�?��sN�g�o�a:�%
�0�T��&zއ�:�I:�وs����6o?7_p�(hg%6)����u���Q/�[�����ׯ�Go�;C\d�!M-
�6f�ˉ@X��DDs�3���N!SM��Eގ��6v�]V���8��y:�В�t���K�bQ�sbd���-M�}7��堁��u�֡���w|lk�넕����
9��Ijl�}z��1X�f3 �,R�#���q�5�0���o�Ҟ,���X�ܗe��DM�;;ܗ!�#c�4KD���3s�Zl��T��������9$�(Gmɑ��a,�
�K���q�,i�3P9�Ы�G�><s�u�B��l���@��[�(�|L
Yyb�J�)H�fr ��BS����cӦ�k�M�7֯}���&Nʟ��%�]��bX��`\
*�/�zYA:Z�hwۑ[�ͤdLw�ǧ<£�%�?���3$(����Y�ԡcn�����TĤCAq���\�Oފ�v!��_�]w�9Φ�Z&%�2	\v`�$1+�+M;ly�y:�
z�M0�2��9�)If���4��Mr�q����W����n)�m��l_v�!a#.���W�R,�rA�{ؑH�*�Yj�*�HS;5�)����w۷y��I�F�K-1�mj�rp<��m��\��Nj��C���sZ�ҫ#���n��+����@�t�2whK68��4��E�2���aR��s|0�� ��ˬdX����*�]hs�����T�ط�g�ץ�q.e�|L��̇�s2.���e��T�1����óc�A�9��w~ZƬW�^{�3�8��+|�����:���G��ʣo���M�Z��X��%�W9�4-͘��~Q<����ix���(�Ήi�?�T2b�Q�k������'�m��m��ZL�����W�V��N�`�1�v,YME���ftW�;C����u���@/=��B��o'M�f�rœ	�o�b[۶�#�9���s�E��J��S� Pʴ�ħ���-y����1�����-$^Io7�	m��]��.&i��B��L���n��Y��L1c��ie�j��UZ��G�Ԧ�O��S�c*�;Eq6��t�\����w{6:��*5�|����?^ͥ�F�J�Y�����X8�����@	,i5(J-�4R�e��7�dt��`X���N�^�$����J�v���!7��K
u(��?����y-�ߵ����bP|�ɵ�^���FxiR2��Z�Z�X��I��]飜��|kG��!��MpU=ǥ�ě<G��2�B��QG;	=LKqnFq8���vw��U��t�51 �$S���u�"��d�.U"�z�~�(�F�ܭ
�&L�3��ŧ�9��OӅ%L��ҹ���,كq�_��g<������{�U"G/�△�҅��9�f|A��ޢdQv���b8i&9۲'�xr��Mэ����9ӥ�xn���ن��W;���k}'\���d��(�ӆ�����Bo�(����8���>�&�*���70��f�O�(NosA��܇���Zc�y^����Dd�[I? ��r�#��# rv�\����p�AR�;�Jzr͐'��<Qd:a�s���q&=&i�x��q�l��������׶%�93� +����`��#d�����v�9$tz�M�4���<◑�t��"�K�DH;[��hPORy,㓓!Q�{����C��vDmy��oK��8C!m����(/��.v�[�C֋�����i�C6}�g\hަ��;T����wY��S���F��h�̡���i��R��R��c������u#�h��$܈J2#�E�;�w(dA2.�ئT[1��~��_qrYsy� 3+�Ni�T�v��0��G2�t8 Zt��)H��r�AdE
 ^{rYFʔ�&k�S��'�P��'�a;���\Djv}��٦���f�ڸ��܌8���y�xmDG�r���G�V�C¸��R��dM��NA¹��kb�~�`�O�� B�DR�������Z��J�0`���yOj8�y�l���D�M�𒏪��4�[Z�U)��y�-�8���+����������E�L��)���|C��4#�D�Q��5|�n�s?n<*Ek�eh��m��� <J�8�7�a�>�k����ݫ�H`��pk������y���p�� W��[�� ��~f�
Jת])V�3��t[�Il�TdG>ve�U�����A����4`Q"�������~�"$��[A���q�b�Mҏ������'�AUb���H��+.�������>u(����?Di+~v4�]$��F���b���>�%2;x���v�,�ii�oF�i
WM�5���Wv=E���)Y3K:�\�s��!%��X�I/��l2T�|\�o�����)/��E��9��J�l(©Ar�<vA,�l�IL�.��� ,�' ;�
����Il��&Qfk���_��W��5�}��H}���.������� '�]�[Q$.���KOǀ���b���=��e�|�r��K�Y�)ki��x���Ve��m�dG�֧�4/cw�����dw�*6<S���:��V�F��Y)�8K��㻞d��ҋ�*�օ/�)�o��V�&+�j��ڂ��u���3����I}��\Z�|��t��?�M�3g�ؔ�G@�T\�R(�X�aӮ����8 ��b�����s�w(ͤAP���t+בg����}����ڔO�(-$=�צ� �<��T[���z/j.��w��X��t�O�N��	�ϐIM��d��3wmHA�v������!�:	eb|���0�0h�������^ �`��g�ҍ��7�Z��L��ȳ줷�t�����F��%�ސJz-�@6���$}\`�jE�V���7���]$Sķ�JS�����ǅ�6����G8�6XcY�olA�_��	J5.�b�Bq���G��|�ɖH$C�s'���dټ��V�q0&���~���*���>z���A�N|��F��j�Ζ�%��U�X��7'�Q���V�n��N���t��ˏ�pXIp�֛ߐ?קa/�-���J�'�p�@��iJ���\XH�����H�G�<��ޒ8�8s�0���
|>�O{��HL(��/ M�e$�uN`���1ȋW�b��K׃���cA��ˣ섘is�>�$�EuB�8pX¥�q{�ե@�.��R1߁�]�����D��˗�v�fl6}��`�/>$���jbY[���',x!-�3�a���鵠�29�
��F	ٟs@��@\XY��0i\cd%��َv8CA�O��*�+���/?%!�&4��|m:!7Y9&�3̠� h�B�U������!J��j��HJh$� ��ⳳ�^�^%��Q/;��Ũ	���?�_D�*���y$�%�j��������8�8[���Q�Z�HO	������;��	�Mg}mD����@�]nUf��3���͜o�N@�{�fi��x����m�����_Ǒ�f��*������JB�MSg\��>y�����N>�C�B���w�q�����"� ��(J��:B�D&O-��`��B�IY{�-��VLֆOH��$Settx�Eʡ���s�ǣ������Fϫ�/�X�'S� �+�>`OU����Y�[3�zt �7��U�����W��C���F"���(<�EO7���S5j���1���KO�׳~�C��w>�����#��}u���,��bƫ�2ҫh�p>���|H�h�;J@��Uu��4ZZD�t/�ź�s��3��H�*Y���U�z ,R���D��t5��6}��iLʞ]��G�:�%)�%�"P	k�b�2Q��]����ÑE����q%^z� �C����v��V7/��n�d�r{����(��V9�dk��B��~u��O���6��t�[�"�h���J���i�ϧ�n��3�S�	���`�o�E�ꝡb��VA�c��)���Q�dz@>%)0��~T^���vk�/�tD�d��ù��Y��X�n��8�����.�Y��*�Ҕ�9kIKR�s�S���`d߽��? �tyQ9J�z�U���je�I}�8ҝN,�x-�'S�b%`�!Q�Z�:�Q����Np�~���Ł*�{a�+ۻ��6g9�h90
����jlN� 6s"#��I[�掳�1-�Y�f�m�^7���,Q�6�|O��N��x	M�*	L���O���MlJ�K����ܯ��5�/1�R	�x�ю|!��'+s��R�8�K�nT��F$�0�t����(�a^��t��Oz�R���8�u����#U�~�oA����'�4��MC�bV�8��o.M �h!���*
D���V>o �eyP��O��}��!��>�q��(�'��ТLj+A_��2��I��J�n\��1/�:���cւ�D�eP��$�r�az:�4����S:ԧ�����6x�xB2;!_���D��&r�o�= }��pw?���Tpb#����!��jl◥m�J�d释�-�'�Z/�
��)o`�̭�`+�ŏz�z����`!�וC��7��]<�~�`ODx�\��� �m�W�O"��2��M ��鐃),ۍ�|���hE_�k�UE4�"�����/�G'�m�kQ�-sN��`���I3�7Cd>��4�:U,½��?������沘eD�����.<��_��K;٧���[)�\��������D�,q��r����٘&��ض/)f;�
�mA�l�SRB,��o��
\�j�f������A.���ZH8bܮ?Z�e}�W���f�c$A@ܬ̶0��,ڦ>z���K#�[ރ�08��Z�īsgqyf@t>];��PU�O��y� ��g8���V�4��fY��&+��v�^b��e��H�o��֬2�s@��8���"�C����l�82�6Xح ��cmvl�xź��2g"gp���GS"�Lw�;��Q��d��C�����!�@���p7��Ͱ�\0"f{.O��"@[���� �$?�,bT��g����lo�S��0��"f{��r��p4߃nyȊ&�O���<$��1���]��mC�h؃Ŵ�v@pi>Ñ���}7_����RLV����UMy-2Q�\y9/A������h��-�`D��f [��,JV��qC�@Yv� ���ViE����3=:��{u6�q;���|����у?tI?���:K�2�%����۾Z��h��etV�,�ZRJ*^���Y�2��1�w���@�Ǆ	(�����5Euq�/S���s�n/4y���F�~g:������D]�Sa3��[�+�Q2*��E�|�m�ۜ@�۳%	�;L�_�W|��#O��:�Y�5{�g���	cK�i'+GYp�t<�h*�tx��b�j��e$��4$��"u�%�3�5����%R��]�r_,g�6��f\):���c�bR��`̓�d������}��*�l�5ʽSK%�6��j�!��S�Kq"���[��X��s�F^��5��6ێS�?����g��-䭧�W�����l�Ko�3�;7="!���4�1lD�[�¤�K������)�N��2��k���j}�]�4��O�a&gؐч~�aW�����L���ܔ��l�e��#lR�g�A�Fx��蹉N��4K�����Z4͊�!��!*�v�y~tL�"m]��^v�tC�����{�n^�f(@eL>�n�	N������T�z���J��e��M�Y�|k�뮥��w�[JN��KZ��'�C��5���x�`�
��_+R�:6�*P��Lc�����s�!�
�66�l���;5�W�@ؽ�4��VH���SbLD��5��;�ۃ�_:��*�$,�ɫ$)�O��@-;�Rz�k�mI�7&�#�Y��>���:�Ds�J��W
��-��.���ns�~ۗ����P����?��xᬽ //��IiX�~�}>b���@�HI��$!CN W�.bt�A��8�ĩ�>H�y�!�jY�<��%�G�/�G�Xwd#����+ �" �\5�kg\�3����R|��,���e�#Y��kDK�B�}����'Z������� ���Ey��]���F1�����3�n ��[G`XƅhWr�(�ݫ�	��M�YQU��e��>��|Q��L2jơR���J�I�J��q6���5� ��l�㻺z}� E5���F��=�� �39��^f{�L��[��QS�C�7	���n�����0��y4h��X	�P�P�PŐZN������� �MZ�g��K�~�s�u$0ͷ�%��-�ʝ�;�<cg\���/���l��k�[���4�*W�|Y�iZʩ���`X�7���O�I��3��k0��Ժ�m�(�˺p�S_Acg���dk�[��SƊ��n�H��w�2^�9
E�W�X�=$�G?��Pa��n8)?O��� 3��"<-t%8�Í`���b�Qu��B�t�4L��ϔ��0�:�zq������W��ט5gȅd��Y۱&�o��Ȼ���4u�lIW:�D �a�_5�;Kډ�)�Q���@AiB�*,�M�x�ʵ�%��g�iʝŶ���MCݡN"�9i�$4r;�Ӽ���}z<C�oPy�r��e��	�͐d������A1Mew�V���XRi�;]+V8U�SX�H�+�6{�:B�2�l�  �{s;]��*�e˛��i��N�@����PG>��5����<'�
� ���jK��P�o��#}��L�^+ �9������
�k��?����3�U��L��� �ԝ&�n!�\���3����ȃ|���8���)��'�e����TW!.��]�����tK��['�Rc��r���3o�|r\��-?����H|��R��&���wn�]٦�S�Aȟ��.�;6�KxD�	�A��q�����_�{*�^O����<MY�DE���)��[ҥ)n"J�p��F������^���(I��L c�5������,�@�6��J3�ӜN�
(�Set�Z9��Jc@7��໣݃�wqê� ��)��{ޤo�7/zx�{��	dd�ϐ�ꃅ-s�1����	Ba����׈Pܳ�-3�j*y�֫�d�=���7ZY=�<�#��	�MB�>}��4��R:���_O�Ɔ^۱��{��bJ�d1�!p{%O`=��8�;/��5����VW�j!I�1�;�������P�%���sU_Z�'�v������e�IKO����i5`>�v:Xce�N����\m��9\�?��z�/|��`=�9͙��D)Uk&�?w�|��׭&޶���Xh��nT��t��o'��X����^4������e��o?|�F[a�U�P� B�uN����7�36 >���o7��`*@�>U�j�ڨ	wv9O �����p��Uʊ�K�bWK.}ɠ�
�?��F������E3 ㉽1,��W!���4�ƾ5�1g���$&���BS��ʛ�uv�ʞ�B�� ^��#	��%2�ɻ�D���$*��3�� Y_�,� pd�������!���A_��X�gY����:
��!�~~\G�����Qt�-VY�L�i��.�;r�d�������k�ڥ.z�0�H��{�,4�*�K���4�|��x���ߙ����_� S�K�_T<�&�-��� tQ�\�&�xE4��3osMV<�E�*H*n�6ƛ�ۣ��0Ⱦ�ߧ7�#XF�ӣ�����`nc/��e��Ҙ�8c߸
'
�s�I\�@���V|[�^r|�߳GpL�RSK�`'���i����5����:8x��Cy[��D3e*�Gh6T�E�S�\}_�U�8�i��d�k����\�bF�!DG8�5��h��j�:�?lo�06l�KH���ȣ-�à
O-"��?}P��K�7�_7^�`L�D�����	1�Q�3�Uqn٨�&S1+_���2��D��?<x�}s�'�F�.O��6���6ߛ��U����� �2�b���4R��T�%�'�,�\���/Ք�Uh/
�qҜ��nF$��z=c3N�S�/��Rc��Wc��`�UT��-y����}Em�%��|)�,@����V0����+ߓ����Y�=%�����x"�9�l� ��b��i�Z={���p��`�X�M��!戢e�t�5[T���2��n��$��������kka`]=��:#	,�Ё���̰�mX:�v�Z;6~�����q�_ڎ�m��ӵ���3ŭ(�\)�N��%W4#&�̘E�آ��+=��r(��;��
�qyHK���|�T���ږ	���R�2��"�����x�BqY��}��9˪�X���HfD�B����Uz�������9~���<yE�3?=f�>Щ�68yd/�;���0����iv�������Z�)�(�~����-=���B�eӵ���R���f/��	q2�*V�&�࿃Q�
��������}��fH�zU�vl8Bk��j�^����	孫�xOx�x[�Xs��7S�P�d�i�v5k�U˭�������h�'t�W�Mkǚ���Τ&��2B�Y��"m�>
�q~�
H	}/��o���v�R���B�t�n�!�4GI��A�E��IN:^L�8d+��۫d�.;$R������1w�8�e�qP�x�O��� |�G�p�@�+��J]�	fRq~]���ӻ{�ɮ)��`�$?�r\%6����F���/�v廟��W+�l�ƈ�r�t�P�$6��iῄ�(�Ÿ$rs�j���0�F�*x2$�ù��?n�G(���k�:4�QN��	�pE��&�|hE 57^i�Mϗ�Y/����8����B�IX��^6�"�w���r�(Y�ܩ��	.��XN}�l�����} ʠ�����%�c���n�:�]���ՆF�r骶2lXe��$j����e���t&=Xۂ	J7�A}�J��#����ȉ�}I��H�QѱAy������M	'|j��;"�Gy�F&��ƛ+Ήu��B'�?�����~!��{�'��3Uf�̞���cp�Ra�7�v��-TAn�E�F�G�V��inn��M��� �̭��f?�z��K^��,�(I�n�S�OA�#Z>4�%+@�ӽ�g0�?E.��8�T覤T;��V���\�|X������<mp�Gx��]��O�o��\� k8�J����i8���B_�zϩ#Y���i�=��/��{�2��� R����_��?�MF�q���D�W�l_��v`��a���-2�=A��(�ڋ_!�P>4�z�"ˈFN��&������^�E��	�}TUε��Gu][0��4��E���{sD
?P1U�����9�+�WjL�	R�գO�iyH�)�R�����m~0Y�R�qe|�@:"S��D��,틵�)��OSi;7�D�'Md�(��/�K�N{6!c�Z�$��i�h��6Mj�ܘ%b&R�(5�|i/H�}�7���~�P^�,�^�J#��(�S����T�{�����ä��F�@"i��H�2l�����.ʨ�Kĵ������'�UJ[�)@HH��f�|R��K�N"C��%z��'C�L۹\��z� ��oC��m#-ϰ:�tG��,B�;�9�~��#��=Y �)0������ݚ�p�G�o�j=���+���l��@_���.�9вx�����4���13����VS(U��B�D��T)����s��6W������HT k�{�C�	��f�M�.V�Z�H �;�grԚPm�/���OOV�T��#�4�K	��m{/8H��tD2���w�.p>}�d�:]).��S��$o�ByQ��m��s�.0�X���ᢾ���5L�sE��^m���#����ҡ]��]�N�b�<+��m�]aPr���x6HL���.)1�T@+�ܞ�T���Z�"Bc$���E��T���O�~ b���d1j���� ���n����~x�����+�{{��83�W�I1�v���Y����r�?�'���l�|��� )�LZ�y�4G��l���^I�x���A3�V��a�"�I��~EQ9���
}M��ޑd��X��nh�����G>�:�?C�XQ.t@L^}�f�'%6�������}J���F(��`N��M�ZR2�����lӌ=a&�s }�$�P�����d��i����ԊS�Y�e���h@���q�Uu�����w��NS��|�ޯ`�Y�6y�AC���	�U��+��ԫCĠ>�-Fq�H�P���|[	jޚδކ�O�)Ht� ۺ2E8��A9U�W[z��O[9I;�,���~|��FV���p�-�U_�䅴�)�Z����m��G+K=�����dpsU��ق�Z!��;1Ū�/�L&4����m�o�ި���9�7�@�ʝC���Δ?��y&���G�z�	a9�&*OEC�jn!hWkv�EC_�j��m��8)�������7K�Yh&�9b_���?��;k%Ī����e���
ۜ*EK��S�*�>YT�q��[rY��p ��6F���Q��k����F▣��mn�=����.�$d��B��Nf��w��D�#߮���E6t��Y/��غ�4�i��W����#��MG�٭;��)5�N��7cdC5����5��`�����b�Pa�+��QJP�<P�+"�Z��	K���0v���>P�/ C�j�g��6j"���s�Ry�ʾ����!��A��*����gs��df٬hR= Ě0��(XM�E���t��f\a�[�|��ι�Z��F���E�m�e�B���n�;�tz��S��3��̉$����{�9ˢ�tUl��Ա~]̙�/� "y����Nq���������X�/i[��֖�r���>�Xյ�?��&����w��%�-1'��c��\$òA�f�t�r����4�w/��g`74�؋�
���2(��zV(TH�ܤhp� �v���n!�Ϩ��2bX�p��+���-�_��~�`E,�L�
��Ra�ɋ��|�6�5
��E~�U���U��!v�9O�$գ�w4v��L�@ńM,��g����T��?��cF�1UZq����ãL{��4ׅI0��,}�X�u1�X ��1V�a^�x�t#P� ^s8��)��4�M3D��*�F���+<8�����rl[�u���M=s���@c^S�O�&�NJ��rE�ٺB3�����I��x� �Tl���%����'W]G��w�����9�F Ҟ���4m30�0#�־�Z������}��	R˳7�]�y_w��`�|�Bݜ�]��e�F1O,7Э�H���j�n.��n�W�=����$:�+�2����Q�Wu١�'?:�i�e"����z���#F�#����ХŊ�ޑ/���w�Ǵv��2�Jې�`���栳µ�A��\ʴ8�Fe��%�C��=)�d񝯡I�Gz�:s���To#�X� F�킸Kʧ;7�[)��1�9��S7�	�϶eH��&so{���F������C���C�%"|C�0�$�V��qi�`ȅoL�-�8N��Ip��Xk����`s95m�q�n�foNm,8���
��ѰC�	𫗢���J��,J���a������>�x��(Vk�J
���]f��ᚴ�*Y��J���O��������`���yP[��N1J�q��A��s��1o�t�Cx�h!� ���ε9����.��1Y5��ꏬ���a�'�����������T�k�af��S�gO*���B�1����]ec�F�*2Afˋb/ړ�	�!�)�K)1i���uu�����Ir����μ�s�K���"o��eb��g�ؚR����{_�ئ���еGҐ-�	�7A�����u��X�1��C<�N4K�C��x�����1O�;RL���UM��Zp�X�5�rNR��6��\�*�,]:��ZA�������t�Ͷto�X�?]kq�(6�p�����Ł�r���`�X-�Ab����ۅl5@L<��跅����)�p%�'�=��` ��5�h�fVn��*�y=%w8�]�t�+����D�NT��5,^�ݞ��"§yI��Cd��b6-,L��4bBɏcԘSW�%gl��0]4�>A[��3?K�C���F��/��<�=2_q��-�_�&ep�[�Ȕ`7~m�כ�z?!�E�9+�;�;:}�C�D�~��UЯ%J��K߸`���{TLS�i�~�gW��1���ZY	��ا�ځ�9ٰ&v��/�������������h%�M�=/�@ݓw4ShR����
�� RJ0wlG��,l��J7٣q8Mt�o�y���c�e���k���J� � �^�v��v9E�_1(��v�>+�fY<U�Y��EP���� ��r!+��v�"En�@��(O�8��G1�r��;8�8��!��ɣ��}Yܴa.�8��l^��n���v~��!��í㾠"�5�:_����P�wG�;��o��z�В�Rb���Yw����w5E�g^(�a����U�O����
�5j֍"��Wq!�z`	_����QH|�]Oz�,u�,E��H̴\N��H~�C�_Xʀ�����V�j!�y���Ԓ-�取�����ѕ��t���K�Hs���d�_�UE��s�@c1?�!�OJ��o6�@'�����R0.$�������P��-Aդ�͑~?z2M��U|q8��k�]9����ƈ�Xx�8�
Ӟ���|��R'M>����Ø��%cA��W�g����&�|���i�n��|u�~MHR~��WW4f9�VZ�O�ÜX3�k��e��}�0?GM����^���n�v�Ĺ.]!%Fq�a*f�D�7W��1���!"r\���ヮ�.>w����ۃ��rYa����b��݋�L8�'W����B�C�!F�h]R���Fi⛟��̖f^%Ą���6��j�q������7L��!�Ȋ���x�3я:0c���U������4�45*�]��_f8��2�՝�vշ��mVD�;�MX�1��T!����q��H�h����`ӳv|��X��;�G�Ƙv���������4���r@,��`6*����οb2	4wsb�o�K]��]�(�䣵cv)���/
յ�֒"���T+�]!]8#}U�����W�R;�7"��I�I�Q�S{��:z�_�l.�e[�OL������<�����HZ.-�c�{a���m�%�Ģ�L3��]j��d,S�A�Ζh�z��y�<
������ĬYȮ�)�-�:��eD^%����g�o8�=�l�7:�9K,1T;J�����jO������:�2�,�%�F_�M�r��L�(��տ�>y��keVl���+ļ�iym#]�g�X��Tð�ld�}�����_�(��&҃/��C���B����j>�B�z>�F� ���������B�S�]��T;��8���{~�b<��1s��V����ݘ��� -P�cu�a���z�г<'����\O��J�CD�/"�M���;VV93��Ff� f��I�t1v*�֖F�U6���QwN�(�V ɇ*oB9�[�g�;�f�%+ rV���1��<��hwFQ�{��Z_�M�B�[���g2�C.����w�1+ި����J9�M�Јsm.16-�1;h[b d�v��rF+q��>�iQ@�w25^�:�4E"Ts�L�e!�Al�_1O��������	��EŃ3V��!|g�9�qiz����(7�J��b[d X��a�1��$�Qmɝ� ��Cz���x3��&[��QA��oP
נ��O��|:���^�;d�S�&�҈4��ش �.ơ��:�M�����'�:=����PW��)yD8nG^�&/k��.��\�kD���&���2�w�-��I֐b1 �{����n�6��̍
�0cH���f2r�; ��Sn2�u*Rf��D�4�C)�ܯ��W�.2%Q����}��)�$!B CB9��T~����������Φ����^�
F�p׏�5�K��ǬL�qt����Zߌ�"2�QN��5�T�&��]�I��r:�.��0�@��F\�t�l��y2`����s�|b��m� �/AW�g��S�a �	"~�x�t��׍T��&T��@����\��?�5�@��Tw��;�	���nX]�&�U��⃄&?2f+�`��j�]�g��c��w�V��x�Hfݭ�4��{�.�	{��y��a�p��?WgG-����i���L��ջ��C���K ����$
�D��N���knۧk��a�o��^����n� [�Rz�'ܕ��v7;��"�4C�"�����0A�R�1�(n��O�ɡX_��J�Q҉6��8���K��[�������N�]�V�F8ݜ:��n�i���?$��(M��qK���]��a�G�yݴ�iw�.����z�22P�p����,���&AL����lĂ���Ȅ�(!�:��F\��5Y��6n"�dG?���ۯr���J�d��7.�e���D����o��:�p�BQ\ܢ�m�jn`����O��%�� �^Y�v��<�bXe���x^�D�:�,, &�C������W�̠/��>;ވ0�a?��[�!���s'
�lVs�*�7'�Mڡ
g��=��2c����P�q9�O��n_�	�*X?Ot�9)����7ȟ�YǱ�Dҁ�"І���Ƙ�͐>K�(;�D>x�:�{7>GA�er[����s�6C����,���^�������%U���Qtl[�ɂ�f![�-�$]�o^�Z;s�+�}B�䦒5%��n!k'�K���J?��)h�R�a�ִFh1���=�u��� ^(%O����K��&�pQ�_\�Ȑ��ė��Fum�Ej3S���O�d�l�T�ߺ-=��u`�ݸG��7=N�qemND��JE��˨fq%��N�(0%�0!'��>,�1�TP�r����U���Y���ȼJ��T��)$׉��ۂg�!�"�O��z�Y��n�%I�EWp;vE�AS��S���7������qi4ȋa�� ���g	L�7�Ř22�mM�Ѓo�z��gj����R���]Ew�*��Iq��G��y�$6�-��$"��Hd�#�["��<@5�F��wH��zx4	]�fɳ���jq:�z#P����p�/�Bʘ�'~[u9q�:�7�!��-�-'+j�O��O�4�$��z��Rm����������Һ���ut�b�i[�́o���?�f��az��C�Y�v��ے�<�0'?�s�}٣�_u#d����/Q_�R��~�5vĪs�-?
C��3��w*d���^��3��q�ڹ^�����N���J����P�\��l��Q�
<\�G�;u�~.;6]�2�����S�v�#��`�����4fu���0V�8������>��R��n��e4�ڸo˕�����ɤt��)HM_]�g����Z�������|QƬ�ZQh�ׂ.ό͕��=����h�$�<3L/D��G�;��j�U�:��ߓ��{n;�0�H<R�[-7�ע�6��B�t�8�!郈M��Ht����y&���XĻ��(��*��?��f%x��:hBe��%s�.iкq3	WW�=����(x,����I��&���c4����t�`d��U�����f��D�ߜ1����;�`� �Q���6��C���G�-�F��T�Zֶ"��+@��C�fN���|�\r����l2y�zx1��Eݮx�n�F	��0�
���7�����or�AԞ�=t�9'�����F.���(N�o�5O`21Hb��b����п�I��aѡ��K����rwQ^��FcL����v�(t�`�~�Yh��ݚ����Y���l��6ѝ���N���#R���z���=�x[����)�C"����i�b�)��6��f���R]��B�\����8���+�ƹ�k������wpp���\�p���yw����_���-���.��5V��2~�"<#i�kJ#�w۞��\7��J�_�6n��(����W�3a��K��s,�^,,����ll#I�d���@M���d�a��ިMVhz#L�+oL�{�xjvA ���"aU�<b��&h��JK@�]�� n�y��"�Ru���K%6����f����{Y�䵷�S�ifN�c@j�(�*�:ȉ��Ϛө�*\;�&t�e���N%B��,s*|�?���r566O0x{	
\���b���w��o`>l#��$�\C�5fP�ɊW�u�n��'�T/C�{��S�q�W���%����o߼��Ж�n��v�Մ/�gs���W���"d���.g\��P��뀋nt�1o~b�|1�P�А�O�n��u[�)";���]Ĵp���ml]S
<���3��g��]���7���ʗx�~��I5$�p�����Wzg���f���3�l%�i@���a&����Z#���ݽ[͜�O0s�)X�'�u��h����u�b���$B�OhK�|���]�6)S~j�C�b�ph�k����Wn*�D|{�-.�8\�"�E⸍���Gz�\ג���}�P�w,��t�W���2.� K'�
^*E��߫�i�N�rv �`Z�����M(�n�:?�@���!�:�C��Q�k�|kG����&õO�5a��ײ�
K?Y�}]v$�D�B�����)E#���Yj�ƊJ�����L����_v���<������]*� d�,����ڐ����Ao�E���D�]��GXV�=�OZ~9[|���h9��H�P
mIHob��z�s�ZMn�I�{�P�DX�)��<���^p,�_,D]p�J��k��iڎ#u�1�sNl����������_,��<t)!$ھ%���Դ���=��~7����XRک-ΰ��C�?m�9��S����=��|H��)����>U��/�R��7!M&R�����I��b�នI�2އ3���^��n9��Rڡ�lB̏��ݲ�H4D7m��uV�$�#A<W���U�0[u~��^#�������Hk!�!���=e���׈b��""a�4�ب#..���+d��Fר���h{�f8����i�t��H럇�E����9�����a��Y~Kpk���t;�>�P���V"FQe�ӽ(�f��)�e�7 ����
�|��X�Bi��`']����ꑶ�aiR��v	��Y MZ����jΝ,��m�z�c���ݲV�h���r�*Ƚ�r�(!�_E�l�{ V��E��ȷ����������O~���9���#�v��A40-�Fys�O-�W^������q�ʹ��đ��s;C��d���
re҆=�Fg#��ӏb��X�%�T��[qUa���R3��b���4`MΔ�b-Cb �Pw����"��،��D"O2/Η/F�M({��w[d;��O=:��l��&Ay�XE;���Z�,?Z���٦}ӫ��OICB��4�&��l�I ��P���|�������-8C� ��S�V�aΦ�P���x���:e!�������Z@�o�����%��0vwi8�ʨ.��Ţ͑�*>{��|U�j=I��6{�i�'�=�M�-�r<ʡJ�O��v2@6�oNfݎq��J(��ۨ�IB�|8����tWW�t���V�t� �U8��RЎ�8C��c1B�=�*��`�2)t����:��j�X������P2Q��/kU$��N���ɷM��r�-'��u���M'��+Z٩C�����E*+6�x�M(��޹�8<$�S�P&�W?y����H���^��;�M�3��]����d��MلKUl�ٟ��;[��Ԑ{Y�v�gc���zl�^"����aI�y���B���T�r�8�����paŊ�O������[$��"��5�7FD�Q��X�e�et0�s�<Quۅ���Ő�#@ ���1�C���:�m��X�\�i� Ȣ}�3u͞�o�ʘ��D��6��Y��evs?�2g���҄'����3�\��)6��y��X���8g�/�h��Fw��sX�n��2�7?��'k��� *7)n�����A��l�E�&u7ʅ'W	�&�{�r�8Z�D~I�<n41-,��s̖+J地�8=̊ʟ-j%qv�L1űm�Ղ�Q�&�^߉��-�S�����bbw$�[u{�k`�隚1]+��U�����?4x���]-���v!��j���cF�-U�`�(b�Dw\5^�|���z*MęcUF/�"НՇ�^�$��Ӆf9AGx0����?��y�'BH��' 7�!��.�v�����g�f1������[��vj�s��T�4�O�|8�<xj8�X�i���2(�2ѝx'@*�3�yw����!���w-��Lg�_}b���8��M'C�ˎL�9������O��NVi����5�&��F��(�)��:��=^��L�`e(f�a�d����N���Ӎ>�y�k��$�Şc9�Je��O��Q:�ߣ��I�n���қ���P�1G�]˥[��R"&�Z>կ�҆|jR\z�9����]ir����!��ak@!��B��ߟ��[P���/����&j�Fb���TR�%q�U�ta�`ܬ�u���@�4�ǜ�!�1����<�w[ckq^YJ6�>"����e�Үs��+��n��^`���� ��~��F4	�mv��tû��J��@�>�����%��+�_�u��ޱeS��7A�g�s::ԑ���"�BKo���n0 hV����Gk1�N���x���j����a�^8�g��و�[����g�b�����T�ٱ�H��r��t/�C�S�#_oZK��e������zt��6�Oon�͔��ߓ� 6�����(��:'���F� s�{�!����ت9����«-�=>Q>����D�5Q��O��d���fݤ!KBTT�ZS/]����Q��F�+`�Q��������W�A8�޳��y-ʦf��Иtu	7���S�y� n�%J��=ʖy�"���C�^�LF���V�t���1#\��=����y:N5m��һ�b"�J%j�������@�i[?�2?������`]]Z�-���
�dJ�J@ o�tr�L��+�]�	#�Ӄ%�,�U z�H�ͣ�7��/{+�3>&��'z\`  ��bpA���R(�����,	dZ �٪]LHN�l�?�z�	�Ѣ �yq����w4� ��a��P2_-#�����A(ʷvh��u�4G=Om�>;�#Q��˲V4��X�7�cXdlR�oi������f�1oѰ*�ʪ>���������iNN�H��P9f��&k��gI3}&��j!�^��!ٺ�X7�T:-���bK���E+\�3�GW����'h?��\�Cm`�`}IB'E2�Q�o�vk0�%O�3 W�=�hަ/rϜ�ݚX��y�E�}�����ʜk�'>@`��{���3�\` �kYc�Z�L�#ٮ
�T:�lЏ�xe��G> X�`m��_Ck�%�~[��=�Z����x�q�r��J��_�T?�A`�^�q2����JΟ˼J�c�Y�l��4}���o�hR��-��	��
k�W����gZ9��E_JIi��E}[�> 0��í�Lm�F�'f蛫�7�s�t�R�%$�^��m׳���_9���/�95�����QZ}�A3ub@Ny� P���6>fc8����UG_��T4�灬�����"m2���dρL�8�V�\{��_xnAI��WBж����\�듄���'��D�?�xo�7�P1��Z�z����ܴ�=w��ҨR候��e%4��r�@��*@/r�Î��ջ��2�.��.�I�c^�?�p;�}�L�0V�O  � �Ĺ�Ԡ!�_L�+������;�{����9�Q.�<m����$���#� eL	�ݷj���_d�3��S�k�цL�7����Ѫ��)|�����^/�v Ǔ�����(� �˰aF��B �ԛ@g�o��t-�������
����s9�=&=��v��͕L�V��)�X�����P��㌩�V󒺧�Ǆ��o�]G�{G�m2�s��=g�n���,߉ϊ"��X�վ���uvs���)Cg�tL��jP[
f���!���+�=���%���J��f��EG�.jr����ˤQ�@U�;���؃��oĸt�+~�
yO	����>�n���	��i��ɇLn�>?j4]�nbm�4F�OmP�5]o�����\���8>��u�S����Ul�|�/��|���O�<��Za�Кٵ'R~%2)�Û�|��χ��a'x�$*��f���W������u,hX�R� ��{����4W�d�̾��Q�q ���0z�3l����N���	����!pv�tK���:xCf-wwk�}��`Z�r���$j�A���j���oNVW�de��F�謁V8���ك��y�C��<����n�ws�l�ͱ�� �|���-R#ǧ��@\z��^&`�!�3h�f����d���p�3Z�����\L7����}�d��6JX�YQ��@�7S�߮O�%}���i�"��� ���.kH��Z��I�&����}̩�.��}���0���6�meI�nʒ���09$O����]j�V�EI��_��6
�d��}��E~Q&Δ��fS�'S�qV_V�gﰦ�8��P�0��,Q�p�7g�f��"�w�F��t2�_Бƨ"��TSrM�	YzI�G�>�L@�s��2TȜo"�yq4Ըz�ZcB�p���ԥw��RU���i&����T@ysG"9&Ȏ��j����Y�~�C��hH�ězt��s������R�D����a$Za�C�Q	��%ª@i�/HǱA�N�f��9H6�َ�� Z�X�������?�n�=9,��jO����u���Z���&佤ry�J��dZ����u�\����#���!":&W��a}���`�����߹l���3�z���J`�5{^'���"�}�X"H��rHTU`vnD�w[6�Dugl�}����K@E��@���I�-I��
��7��LO��G�����=����X_��8ɋ�����"��7S�{���������
������ߌT��E��|�#٠ƿ�]o��������u���F6T\ɸ�)eK��C;+����#��2���9p�����3���B_���o�"�����Y�@$��u==�'�~ъRdBxȾQ��/�>A>���$}e=�n7yu��w��Vd���]�
�@r���$�F�t��1�.y�����^��Y���$�H3�d��Г�&���X!>+�3zG���&!��"��C)@x����у��X����U�ԑ5,�)dϕӫ�PR����V��yfȂ#�QS���@Y�)8m�����CJ�7��
��X�,�A��������\�
�*s΍
>v!b ӡ��8������+�)�x8"�����LX~ۤ?�%!����V2;7q Ѫ����d�jB]�.}VJ@�d�V�>��b�,��� �Y���^�@'�J*Ǹm�|HM�`)��䔂��"L/O�����DuLpy��M�!وM-d�*�hVW~��lƼ�j�Y{�8l��w\���2��#����v��x��\�����;$��%�o���r��ص��ـ�ٯ�~Ե���N�����U5я��'�~fۼ 1c������ш1��̔�'��y��4�L@:"Ӣ
��YP`X0�qZ���[-�x�.�t(��hu�b�Nt%m�|�qKn^r;<����'�t��"���dɑ�gP��4+�F���#ʔC����]M=����b�n�����}��AS_��A��3�b9�ay��)�&� �	 9�]�4�J��@��k[���,���T5O�>Wd��{Q��q9�US���ϫ�іJq���z�E�ɱ#a�d�~���$~���*�LA �)W*}���j3�s�R���,C���3._W�s��.�O%5�q��^t�Q쳝l�^���ĉ�}�>�TNK�_��ϴ��߯¹E@�����x�W�|�T����56e���`�4zS��%��&9��w�eÚׯ��5-t��I��;�=0J�0T�k�Da�H`˿�f����Z��"��m�~���[��I�ޭ����c�*JӒ����Y8FN��J[k
�n c�	5=�����nO#W�L���]�46��'x}����ȄP�8�ԭ���qm(�m���9�k�J�ߘcWU"���\m{��U�x@��v�~��aM�;C�g��o�nKJ�&���?c�Z:F����7fcZ�����M]���^�p��������M���]<&M+������ރ#��^���ѐ%&�Uk��&�5�K`��z�b���P�l�]A��p�#G�Un�;_#�׷�A����'���ګ;���i��ڂ%�FW�;�D,������p���S���A�Y'�xSU2��/�=!�FZ6���	�!��ȕ�6��J�;�c����lv�Qpu]����)QD��4�%�vBKŹ��!�*�{��]ҧ�Mo�j�$\>x�\�����mi(��.�a-[�Y���>_&�0���؅�'L��~��S���L�G�߄�CD�N�qg�Α�E���? _��h�2xl�`f�����X�ی�'��v�"p�$�V�S�#��_��S�3~��Q���s�?ǫŋ#p�����40���>�e�|44��D�L�&�歫@�M�Ģ���-����;�5��r��gsP����/	��tv��q�����;�p�m����{�+Vd1f>c��S�9������#�F��S�x�%��n�0�wȿF�O[ck�}���>[X?<�2�j+����X��
�TҢ1vȪ���e�m[vi8.���jq,�l��f9:8�]�!�����$���'���M��j6���>�	����Cqz�[�$n�u�Seէ���TG��l�����-�)�i��z"A%�y:;��W�([��P�<VMG_�)�,Bo����)�}�4�WC���e���}΅�ҝP~�-!N���>��.Yx���v"p�P�a����=�E����K`�"WL
�6zV�r����-ݮd"���]~����&0ʋp�:#�zfm��`���<���1�������g���~|��R���y�2Hss�G�)��s�$D�+�쭨K��JS�ј�k�{��EP[�� ��ȟRP�L-v����t�S��Gg:F��fJt�FKh�j�D�(2�J��^��KsS���&�_FM ��;��&�֩����$��N�������'�ŧ�V�%M�'���0��X��<q�_ �U�\�,iHp�r_v�t�!>��Q%��o!T}¯e	�ʫrΌ1�/ٖv�kp�q�|?x+%%��=0�a�&殭��&������;N/�^�-D%	��D
��&�k���OIm��WS�����~*��'��f�U��Y�$7;��ҡyA�M[r�+C%4��{O���ۢ� ���iΛM� ��>I9pe�_�p�o) Ƥi�r5(�q���$��#��g�ՐD��Fi�ׂF}� ���m�r3��},8������>���ίi��/����i\7����|E
���bD ����#R y�� r5�]�b�k$�!��G�쩿�_b�0�����ͣU�p���Y�N\x��~<��c���yZNJ���C_�l@h��(Ι��9)��X,�j�P�Ns1�7����5���_�i�{o.�ǯ�RO��i�C����f�k�r���"�T$ThG�!�.�w�Z3W���}�ɣ����ۖ�.x��k�G��C%腽9v��N��"����M��Ƀ�@��-�)}?{R���8���f��9@�M��*2�l����~��Y��n�e��K�["w��s�8��Ր���J]9�e7�K�!صO�O����ʻ���:,⿻��'J�]M{���Ou��n�Ć75K�^���� �?�Bb��ձF��4BC�A�+#y7OM){0���2��y�)VsZ}��=�/�P�(�1�`�U�rl��;z!��#x;�&��!��gOum�Zy�0^�,T
��p:��^�f B����v;������;�c����=��<��`�"E�T#d{�R�쩰O�D������q�F�t$��.O%\~�=|bMF7�Wy/ ^�%1�~�S��X��o3��!����S�0A���q�k����=Y�݉%�\udl9>��W����V�gGm݈Ǻ'G��T�It�du�K��� ���XӶ��y(}DFd���Ғs�\f���j�#ǓX�����_$/�]!��\�Z���JLAfx�."�n_j�ɼC�jan?o��6K��{��8�����8��%�rs�<����L�A����8v�ú�|t��u!a�M��p�3�9��i�7P~�f����˿B�X����Y��w�!�[�U�w��q$M��/��0�Z>��VB�Z�p�2˴�ɻ�p;6���xGA1������	O�;����=彌~��EG�z�����~�^K1xY��H^�~ < /�0-?7R7I�=��rMt���֌�e�@��e���	ا��Y:PĢ��h>���IT��?J8����U(�65���
2rF�k�J�0�h�F�ߢMe	ݩ�3k]�R7��9��S�-���/���.B,��TJތ?;4XP<dh�����ʿ���a~G���\�3��u[|s����˰�Y4����B~�	s�(�m!;ο�(l�Qy�:�gi9�Sq��`��p0^�sl�ߙ��6���m�C3��k�^U��UK��B(�5:�����B���73��hit�}�@�?^6ǘ� �[�����~��Kl�Z�wz�20	 �Wi_!ytWr���q�Y��!���G\8 ߼[�W�w����xP��1D������2o(�#��~1�QQ�*:h��U���oD������(���ɿq�BP~JD�oώe�ǭ�y.{��Q�ڑ$�Rz�"Ϣ��`�>��Q�̌:'��5�H�L��tOʹ�D�
�B'��"�B4:�]ai>?�*�;^�Of�Et�����2z$ۍ��S�o��&2:&��=��%������&;��%5*P�>< =	�]ɹ�x�5S������ĉ��ۭVG1&���ښ� �,z~Vv[�@�G<Q��ٚ:����|�C�,�����Q(*n��{�y��*	b74����7*��	��Ե���{�ά�Y}8&HbGk���Aa)AzD��g� ��ǐ����T��B���l����Z ��޷���'�ذŢ��+/��CR�Э�k��l��ZͿ��@�G�|�>���}���~�U�I�N��&j�V��R�+�T�[=n��ާ���{t,�ޘ�xqF�!�"�~��L�b�T?���BDP]֑N��@��nG<�&�i8������18��Ff���$a�ǡ�fB�L�5g�� B�hT��Ld��rX	��s9'}@���[Qi�O��I�O��u�3�K.H���\�P�×�V�ĸ��O�u����V �U'�3��6�°RZ����Q�7CλT�Ҝ���LE�K�B��xO���D��dE�f����O��=��3�P�l����3�&�=	�3(�O�avE��g��!o�������[\l�/���q�lJ�t��K�\�;�X�CK��A�HoTV�/zS	���9����vN����b�~^d��9��Y͚�t���(ApY~��8Y��*G��p�bu^KouX����H�F����	�P�)��/���[Iu�?���f�<���5��d>X��~�˾�`s
[�1��7N�L}�׶Z��(�t� �9m��/����فG|���g�>֒�7^j�@5�Mx��hNK���d�"_��ڪ�x�V�����a|�<�B.��$���G:����l��I����ʼM�j*"�U��/J_��m[��\�Uw#���)frR����?x��s�pi�q�s7lp(#���?d��9����T�	4��BDK�ڳ�c��E����M��(��v��J4�֍��%lYKZ*/�w,C�0�@���6"��w�n�J�Y5��Ԝ��)gh��/{�����)5Ƴ�iX������yʶܡr�7L�N�;j�=�H�S%Nm�w˲�&5�o��_�b�U�M�fEc����`����iG�ĳA��	��.�SA0M[%ήmP�F�.OyLޛ����_0�� g,UB��n{I���v~_�_�k��莉�wr�J�4�/[��Xm����+��*�I�JfTz;���W�nu:F�z1�S�$�ߋ:f�b��;���/�į�nU)�%�} �k��nk�J�Q�;���"�W�s�-�w�E�3fS�0�q4�6��g��y�֏�x,$��Y���Ѭ]d;����<�	+�+�Ϊ�G%K���b�G�eHpH��D���;"����[ަ�0(��p�0ʼ�QEk��*��P�q��m������ ��:�9z)J-��T/$#�#d8��v�m�o�.t��٫�`\j��|5�M��1អi�;����80�d,^�r6��-�?)i{�kfO� [��khJ�[��R�VZb}�}��]���и2.9H����<�����rS���� �"�ȧS��¬X�`Iu֯�)����i�R�޹|HwT�Ir�<���~O���?���?NK7��:���KS��]�2���5K�����+���ɷAE��W��8쿢>��k�)+I35_/?�"�#�|�/�����U�3O�e�Z+��&��1��3t�T�Ⱦ�
�L(N�.oyV}{!lx�>/�d�7Ll� �D��ʙ*����V��f�<��)�׵��}V-Iː�3��F��^k���ڱ>�a�~��˳;�w�ׅ��=�"�'f�TOkޘk�y^.vn�f�/D9�f���Y�j����+��P������PG�ù����pü�+�����F�=�M�DN@���RȦ�ފ��T	�VN(Y�;G�kQ��<Buq�^��խ@P�SAw~\�:B�g�u�p�hY���4=������D�$�\P��b��u�n4�0��H��Q�-)�(�����IE�q1=v>CQ�P��3V�TpOo5��sEn�e�sK��
�T�p���v�׏Z��,�l#���#���źg�ǐff�ԫ�s���,4N�֕���Z�>����l#Z	�Ҥ>�_��3����tNV�����o	)S��Y� t�ɡ8����\��b7�Fe���>����VL�~d4���ε?K�sD���A1��F��R[V3}����F��M���:��t�J=�9��Ǜv��ː�Lp��؉���H%�s�TEׂ����h��-V_Fb�_������4#���m^��o����X����� $ƮT��o}��p}�e�sN��;�K��U�h���1*����c���a��#u�]�'ΣE%���xln��kؕ�j�x8��w�"�\kq]��fq��_�� E�#�������)�kإ�u�p��;���h`#����-��p�˽�<��w�-H|	�B\p����<S��:����D�������/��ŉ�BY�|Y��$�o�WB�)-�Zv��H��U+}������>Z(��'Z���@y����HLUK����>����?~<�X*X���?/�g)t4�vϼ�(��ઑܡ��֋�8e�4Wk��2h�f�X�~=������+�d�Z~��TB�6�o9�di��%AP���,�.+
���@8���ܽ-[��ʳ0퀧Hl8��M�����F$Wl$؈���g��E��;���dY���A���㡌?�a�~/i�ې,2�u�(L�?�ȓA_8���a>N��+5�f�3H!mB��*�TQe�ɵ%v� f�)���-��](�\ӃR_�;B?%���t t�Uт�&:��P�w}6=���SL���o"��
��\�=y���;���%<�vw��ԡêuC~YD�  �F�'���<���+/,���O�.`����@���Z+0HM���ݐ�&m̈���Po(|����򗉋�+АJ8��Cε�����|οh��#��b��^:����{�܆�[a3�)#�"~]�9k��q�u0���ΈX���li��ćCMvp�?�ӗn(��� N�$���4~�����Uc�g��~H�I�4)2,8Kr�'������Az(�-��GU���S<�����]��y�(��������t��D��G�P[��d�d�Dg0���Y�!��n1�CmND.�l���͛�.�p��H�t H�#@b�aQV����G�$�d3i/[jณ7h�<,lP������9]A�e��M�mǨGr0���E�`4!�'�c15|�
��WJ�L%x�P�v�B\h��,�~Å�q���Z��?7��� H��x��A�����O�����+����\�����s��ڀ�ݡ��98�v������hb�g���OY�� 7��P��ҏ�/[0�]�������Jt� �C~U�P��"&���,��2�f���j��Ҡ�����L͎:��EUq͢����N[�NVWE'���/_�����:�@S��y���pe�����nd�(-{ �9e"�����#5�/��s��4i�$<L��c�������_u�he1���%v���q�05�VQ�F#��ml�W�6Cu���Γ�-|04ĂըwTI��&��%���ّd��H�,����յ�������b@���F�Q�7n�G=��L�=�'�����oF�<��܌����q%��k�}�%�z�/Ӈ��|�B4B[�Z��tE�b�A|Tb_����dʾF�T'�᧭(InC �3���U�s�@E��Xʦ�U)�����@~�`G�5E��3�.�����Q���e�+�ir1\2����z��K���xYb>�K�"f�[JExfw��JT
�W��N�����H�D��7�#�ՇD/�*�Z��Q�l" �(^%+u�jA�M�wI�f%�Lߌ��P�Q�9���-l���eu��}�5���EeS��W��k�R+�OH�C9E
a���p�B>�17� D`��u�D���#�rwx��$�@aQ���E���U�t#sik��@Zcn����!_Ti��K�aZ���#�D���9����f�k����U�����Aܵ�4K�Q�Κ�Z�����ܣrB��zmvw�)��0�{�ϞN��,fA�ƲT�P'�7��媴�`.��T�XY׳e�݋�`5����\H�h(�?/@-�VYQ����J���u(d�Yj)��E�AӣtѸ���rE�q�ԺJg� g������/��.D�M1p�}	5yND�?���AxU����>Q���Ϫp9�;�bn���r��h]HPw�5����A�͞�q�����D�c�`X���tU~KM���=�k��lN�eﾋC:���C�����rm�L��Ȯ�:�oӋ�fΙ7Q�\#�|� �-o�,�9+��x��	�w���}?�]W����9E7�ʰ�E6�U�$���/����/������#�F�ʥ�#��:1N��5@��ڼ~+����5�$�f�T�/"��(��%�P���i�)}.�A�!E1X��&}k�HO�#s��.�)51+�{�n�����
'��d6l嘌p�Ԅ���Z �0$�U.�w��r���گ"#���N���̧����@9����H�H�L4p�~��
�Y�#?ca� 0å7SENd^���t��|�A�$1S��Z	�3�N6(ie��P��fm� v����9_���Ո��ݮN�������پ|r?D{ŵ��U��Xk��m(����ng��|v��!�_^(~S��''ɣw2��N  ���|�o�3念/4z�3?�QJ#�AD�����Qw_���kS([M�MC��7�{��JW��}��K�S�)+@.��V�+��a���������
\�D��.��s��(=�Wo k��A����-���\���������S��,�(#,���g�n!��@;ܲe��5�)��6J�DP���"�s��OU0�E�i�EDi&�R���u�k�f:+�	�3���V��\��"�t�	օ�+����܉�?7d�����D�a��ۺ� ��H��$d"L�4;�����Bt���:�ў0�@�����G#y�ِ��WD����Hb~VP���.�(�[��?}W���E7d�1��Կ����6$¨��mllځ�ߺ��"�^�P싞N�|k�=�l9�&�J��Kq�Z3O
����<KT۔h����� z�K�C��B!�*�V���b���%�)Q_�g@g�V��N��c{�\��|i��<�`�U<1��$�O3��k*H�DkD\F�|�)�v�	�}����z��.=�Y�b�*�8��Ј�:w�����3u�^�Ʊ\,<���}�6�K�C�kRS��.J��]~�Dƒ�)��T������U���9^Ժ��̺v�pH��cwǤ��\�Ev̌z"|��;�U8�&���+"��o��tZ�jH�t�S��/��Mb�����e����e����u����LB�=���x6��KD]��	��i`���Av�Mظ�ܻ����2���ϸ�D�/6�	�$Or��~|�Z�����k��$	 C5�N���0!-�,��X�})G{ί?v�(���B!t�\A���M�㛠�Ae�e�͒%�ͦ%�956a���7��H�}��*m�	2aC����x�G6��~ű�+�����&W/���\2e�V�<�)}y{[�OO��h���tL�MH���c�d���r#�f3�e�5�t�I$=!ּ8���S�#9d
|�VH���wh��9�ҷ�n����?6A&_���k�ǱY��l46=�����^?s��MQA��{���� �&y���m�������]�lA4e���+���8��J������ ΐ|���(�|)�n߭��;+�;�l>��	7A�N� aܡ!ɼU���7M�#�j58�+J�(�l)�S�u���TJ�襽_�-���-C|D��읏*�x��B�r�X���TSv;�ݞ�t.V��H���uP�l��(s��]��<g�*�OPߦ����2��#�X�T.�@Ǡ_�1�IV�~u��
�+8Y��H�NtF�6�f� $`���E��C)nmt	v�5��_ߓ�Z�H��0��`}����'r�2Q&����@�vJ�ݟ���pJ��\�ڢ6(F�LC��\6;yG��c(�4��"���f���;�}j�8ܭl9���SYg����¢�|�D�E
�����V���5���R|F��+���!�<`�����&�lnŊ�����*&jQ�yõ���8���EC��;��0%H*������V�Y��c�*�:΀�LTë�˓wc<��������Ǒb����4J��즚��a�O�I�vO�o��a�c�Fk��,KF�#�񈞇i+g�3rG�a�n9�d�?��}(jNm� W���N�t��>wfan��U.7��Q���\����/���\]�A2`m�N�0�]w$y� ��j���.�[˼���"x�L���i�'Z`y�	[7F*�-5bn��)b(�!pz���}���K`e��	�ދ���i��A@�b�� ��d�K�7(4�B#mV���M�<��<v[,�i<�T��� �k ���Lxd���b�RM10;ly�2)괥i��L[*Ab�:˒hŀ�-�hu�^����J-<L��޶�EY�b$�(��O	l#3�hOPR	р��-\�z^��T��*�'�=tr,���s����|�V�I�[��AP�9��TU}x3��g��hb��ԾcK�[W��?�λ���|R�ş�b*��?�+=mM����f8�NV���蝋�����p �|P
�V�kn�N��5�NPV�U�!�]�0yW����#{�v�KG��M�t�N����!��X�ؑ�����MY�Va.��F �����G��x�y�Ne�.?}+�-�R`��a�t)��+�}ҺX�J8���3�[\�f�VU�����[T-��	g N������VQ%� �6���a��%��e�U��T��_��O������y�p&+������F��q�����m�ꝵ�N!�����$�N'���g7j7B��0�9�.�W�rz��{���"�ӟ1���'+m�}rК'	�J��?:�����X�X���gʻ���v��~E�:���>��80�i�&�cސh��VдCP" �#qZW�P���"���\��Y	5�0���C,Y���T���_xH����!z<�9(a꽃�lX�Q����1XQ�w'�>'&�F+���`J�7�{O�0��˄k*l ���*�Ő$��],�>o���R�|2�vܞP�6���E+�W"�Ӱ<m#w�!�����#C�5�aUyE��f�)�	C��f�@�O}��G�� ���j�
?��{������^:� �"�}:����u���S��G
|���5�Et@�5d�n�=ޑWj�7�Q��i��� ��:��LR���mvzI�Z?�	���p/����*�P;U���( �m��`30^�:|�q�a$����ay��*�~�����zl�{�u���u[�YV��Xb&��7z��B�����OK|j
o�S�la�v��M؅ݵ����l�EL-��7_�\L�0<����>&{�j�
/��KúF.��K�3����T�91rb����z�2�Ƃ��<��-��^���5ز��pj}9}��?b9 ��
��^�GG�5��M)EZ���-'���nu�bDp����pӒbR������C�+1e�)�Dެ�����D'�E	��VA�b*f�T|D��\#�C��J���+�����d,�H1ԵA[���y��5��m��˄s{�&��#��p���n!�]
(��ndX�N

-��BˌB��K�b!���d�������gSS���)�K6{:�V�p��K���6�g�����s���@taW����� 
������s���y�^J��.?n$Q��C��a����2�~A/��L�+��[j#���Pɳ���OߝVS3]{�����B�W�>Q6G��Qo�g��$��Q�<l���8�y�.�1�k(��c>�7�(��%"كs�LPs8�h���� ax�&�W�9CǇ�~Y����:����>��`ot+=�(�O�Yg����o^�q;E)��B��p,o;X
ç�־ݎ���I��P��*l��~�wQ��Vᑥ���}�Ć�G#a��e�E���,�^�$���RP�pjۋ��z���鷨�'��"'':�	��W䢃��7Q yǵ�I�mX��;�! �%����?��yf����j� :�vh5	T�h�dt.:�� �??�Y�ި�Ƚ�1��h����	�B�!z���H�@?��IEMbv̳�x�E�N���i��\��\��a�!Z��xx���q����ݬ��>�S�u�D>���#-+����D	I���cy$��#�P
�Ω�{�j����A6�T�{@� �eX�J_�nNO�	ejC��5@
]�tՙ]-.��!��U��h�(I���g�d{�������ʾ�^�����r/��qLo��A"��͏?�Cy*D6�vs����.�ղ��Ьq�O�h�ڀ4���^��l�lp�P�� SW��y��V��P�-��2�s��q��0��eaH�"��8J�s&$W�̩]4 _laqT��>kˎi�Q oo��z~y6� ���N4��,���"��xW�j�;��ai>������s_ӂ�nР��*� P?=�Y5e����F��
J��hC.��0��4M���[���ԻGCU�.��d)p�i��?������8�G��!%�s�8��R�~� 0�)����]d��)�K"b=���B��K���P~<�`��9���W/��{zF��K����ba��=�
>�v�#�JfA��]��0;V ��/�)��	��;�x�f7�	" =I0�/�\�l��p��SCRҺ��:)ټ֘Vh��']��&�	���ʏ�W�S�&�L����.��ԓ�[2-�ɵl���$G����U��1,T��?<d��l\X�m	��$v6��������b8�&����v��V�F�&R:��o��^�%�����"��Rfdz<q�:����s�l�-�t�M� �7�W�e���ՊL���t� ���èF�{W�gHЖK��p�G�<0I�LS�^������+;$�p��!`S��;����2��j\��j^=�Vך��`���$uV�쏴7#����\���H�-$����q�N��{�^R����&$p�l�
G3� ��w�R]��*�-s���T=!93��ӆ��X���:�h�'ɏ_��F4Sr}�m;<tYbN?$TP����g#��H��a�[����y[9f$�T��[D��a���^mNGt�Xl&�H��\�a��F`xC���wgp�CN�͈���'�<Z� ��-��Y|�q�?:���5�_��k)���9g��/����wU&y*Y�2�GZ��m��Z��h���*��E�h�Xi���ߏ�h��[�/���|r�����N@X����!����-R��Ѯ#��F����,]�i�4����$�x�M?!S����e��n���^���n��V�Y��++�I@K�J��,�G�-�_�@a�#���7�	���\\	ϲ���O<	Xܤ�[���!ˍV�}d�X���"ס@�O��0�X��/�7]��` �EN�n�=r���ܗ����t�{�(Vkػ��=U��PK��^��~�j�
D��JE�'k�Sr�x���l�x���y�x�A�Xc��;0ƚVc�6��	7��nTX�8�L���[�1j1wTL�`V�6�y��gT}��[>-'@W�:��D>ї�8zg��F��O����� b��<�j-��@�D86n߱x�#��}��:���P�a@OmL�A&|����������Ш���q��`C���>��C���-�.�gžA�Pc��;p���ߪ�ھ�|�5ʌC*ʯ5H`_��l��Z;E,��!ar�<?yYp���s�Q�U�O��s������_r���9�	�?"`�	?��]4���)���ե�%� �<��I��./;qa�5��ɦܯ��i���֭�tCk�6E6�N5_tgQ4p\z�{��C�����i�u"4���4��Eb�L�%��c�z��Rhz�=SQ��s^(��4TnXś�p���&�x����˲�!�H�6���|��s6�r�_֌�g�n�/tâ�G������y?�|z��)G�g��N�$��N8���ԛ噵-��Ƅ�I1�u/���W�N��GR/�몕n#N��#P��@\��;�)�g�';	h��G�����V��s��-�.
Z�Uϟ�����w-T��;B�����RA`�e����uW�V�.��JT��]�=#�(ԟV�Qp�z� O�h&��O<i��%w����_���w��u��?,Bq�2�`�������ֻ̍�W�Cu��yD$P�>ȸzAcOJM�xԍVY~Vh@�W�_��ծB��ʽdOA����5����XI��x�3�Ծ�%Y�e�QF�Z�g���b"���/��:J֬��Xe�I�z���9`?i�@
�Č�mʑ�ɊPS
;�^񑋏V��T� b�k���޳�����kЇ�k$b����1Ӓ�.G!\#5��7��W��q�$������C4�-ʷ>zjBz�+�XOϑ�)�l)�m�e��L��
u�Զ���/�,���D�d��}]M�+�����)"Y�d%�`�6�l4'�訌��Q�/�c�TUQ�Ce�yԼ=�(?~��K\% ����p>э,���4t�&��u\��xy�9dl`���
���|�Q�'���Q<�6p���wz���,��W��\�>�x%q2D�́�Z(��h!C��9o&X�WKW����@-D8B?���[E3�T����@Ǩ~>�>�j��ؽe�pt��1G��/K�tHtV �pXq���u\�9��s<�75�Th�d��B�ؓ���n��*<���u<�f�\�P��B�'e�|�h�L�:(#:���i�]sG��6g���Gq�6���@@�x�fkE:�Џc�T����8T�E��KDX�����K��|���b���i՜y0_ī5� ��c	��`�!Dp6���8u'��j�}'��XԗY}�V&���A<���N1껺�*��{+�<t��r}"��z�؎��9�YWԔD|�nଅ[I.dU��(v(�W}�09�s$T/X)@a�� R�&�K��`�_���K$tU�̡l/��<��lV� ���c]�@i�v�f����>+�E���3��n�ȮӢ��ml��qWu�ԩ�X�m��g���0[�_}`�K⩒0�>˄�-s���JGMR G�nh�����T��,�I����2�F�A2Gb(1�Յ5��^3h�е�W�N�Ies]���h�p_'�Ҹ�X
E&�� ���Ŋ��q��..�/�����(/�(�p]�Mu�T�6���9�,���Ͽ|Օ�9
@�z��ͳ�7'�?�1��O\Ev�+�1c����'�P��;qT^�Mr[�ӫ�#��mPg�!^�p
�^׎�C�B	��y�����yD�V0� ̊�46�_�����?���b�(w��1w��Z<�)J]9_��No�qb(I�#��ѽ���Ӻ;It=h�G�C�|�l���+ ��TƲ�t��wp#�����A7qƻ0�l�t�E�O�#���RTif�"��tןĳ����}9)��ҹ������f#iGa��e�P�L\{�cS��2�a�E3�c�$��I�������x�4���z+��9d��q�[�}����r̀QE=J� �=�XJL�����X����:M���zr�M}߳�&:� ��g�9�!3��YC\���i�M����}��`�noƻ��U~��hͰ���_`^�	�Ȳ�YaB״o-@�'O-���s|���2ŬR��d�{q �(+��N�p�ql ��)Ϥ���%>_;�28��.�/T�q��<����;������b}Q�99�C�v#+��WLF��x�q	�$�K�FJ�(ËpF�㋱�x$�&�3��&y(���`1G�
2��d%����&��{s/=|Z_�������Q�CAƒ�{��V`����8��KX=����$�uZdq)���K%{��1q�i�[]ˋ{�E�SZVV5�~7�hb�z��I
�����)�5\� ��p������%�N��:h���dn�w�pH�TMt_^M���c���I'��8,�W�n��7O*�뽪E��?�հ3묱�"�A�eO�~hqa�.������d�h�h��d�ώM[�j�1�xS}����?
� f��rDz6ukSP� w*�R&SΖ��U��p�W�j��y� ��[�����L�3�<��(;3!2�� ��_�� }�w;�
י)�]��`{)
7���;�T�'�E�b�q���+oX|��^<��[s^. �����=lY��
�q ��	��h���e����<�?o�>3�O��"Y"@uy�d� �
ץ����X^Ҧ��G��T�v-�� ��S
���k����rH�9���G��;l?ʴ��pP��8��"�g�4���ק��H��X��˄�}���3�h��1�.����@�L�E(p�JjO��8���d���FG����-��N�N�������6[)��<s�dU�ka����F�U�S��y��"`�����pҖM�g��C�e2�1�I�?
��Xn�U���pA���a�DyO2�Z<��0�Ggj�
�ǢM����N&��8��G�xB�?[��~��0fu>�
;u�Ef�D�<���az���-����X�'meW�K�/pDG�a�+�X�9�h �ٷ�� �s�ua�濹m���NNK!�Į�Ǘ,-
_-$�: �݀��{`���K���j������k��@���wd����1����7H��"H,�ݲ]Hk�r�j�"�֥N`3����,�n��؄[���f�/JN޳��i�@p�L؞�V�1d���^�f�ս]/�Cc{���ѿ6dg]��
)�Q����l�cl�_ɽai����O���F�x�s܊bn��ɔ�.[���YƏ�4��X��s���n�CMe�Y"����p�����n��a8������Zb/�4��?d�7<��@�N���\d ��#�CT)ҏ(��9ys�	_	#�^��,*�,8(M9�l�3�L�w��9��N�~ꈬ#������~��s��K嶶�^0WV�96�u�o�	�����Fw����d�{�hf�'t��}\� �?Kz@�~�C%t�F6��� (� �S��#z�L���m��ow��Z�Ŗj+��D��*b�y�8/'��Է�Q�q�Q�pR�/o��o��N�ƪ���	�5�~�����	��Hx�щ�Ĥ5|m�bm��3�g!φ!�R	�d�N9����.�EEta�g�3�l���L�`�^����z����Ϣ��'��
��V;x�v+q%gZ�x5��J:̤�{�]ݨ�\GhᏜ]#�R��F�o�*������6
��I�Pc��'�]EE��
2 I7O��Z�������	��
o�߷��t����������s�m�b��������:n�Uzмc��^�VWo�aa^v�ORuF�*= �������_bf�:.�E� ���MQIŰ�HW��DMy?�#�#o�d���k7���u�
���A��3�b���9f
 ���\�4��Ĵ�������nm\����[<��j��\�	���v/��	J�Mzl���C���T��(��X�L^�mB���R�/z&��ۙ��gnv#��4z�A��C����oW��mA��Ӏ������K8�o�_��U�Tw��
��>v���'_��NzJV�1��3-�{���4�oa�N(�!�x�u��:��zȈ�Flⷰb�)���cj������m�*�H�b��JU��}��g�^䝟�����?N}p�,BE��@jRR��J�&bA�/�����Pgh����6�<�0�ǳ�QT�����r{7�������~J䨯#5���p!k5J�d���Y&Z��+�D:�?�ri ��?�ڊ��"�pz�n��nM�Xڤ�
�z�z�]�^A:��@_?�tϭ����c-���/7J�@�]��R��խE��p� ^�EI�{h���-:)�bڅ�#��@g�U�5%6.��*�ќy�0��͜����z�(�h��h�/�D}��W�f���\-�Z:��lF�"�	�����Q����9!˷2�"�ݍ��P=+���E�;�	ܽR���ց�;�����g������T����gޜ�4��.��2r��+z*��׫q��c�26��I#GD2K<�k�S�܌"�O��@�3:r�Q������A0u(�:��iùv4~��[���z���Q��X��Vx���:Q��g��L���I���]mF�p�Bwu���`('�_���g�&�G��RょD���1l�d}�կz���{�;�/�~�Bh�RJ�O^v,��hr���1A�s���*od����u���*���G�3q
Γ��@���bI�1��X�aSa%j��mg���d����y�~�s��n^)�R�U6Lܸ��;�6��.qE\�#l�w��֦��lÑ�K�ҋ>�|�OY��f�0�:s�M�%���|�`�C����gsva��[p��׫��]�$F`\<𳼲f�k_��r)�w��@�~��λЃ��e<���A�y4E�.Pv�����œ_�#��˰#���H��jrX��������,��1kw�/���3td���6-`&[[�q?�o{V�Q��_�X��W/�o�`� �����3Wc�ٛ� ��b�=��3��n��蟁u8��5B9���_J^(���)Ea�vr[�C�.�I�.�y%l����ľ��_�]�B��!AU���I��JR�>��F����$)���ź��B-;�����"&�``��3o�v�w���6�-�O.���Q���FS{1u. '�rK��9��}H
b��0��%5�TF�	J��#;���U6��(�馯��5�Ʊ�JSO���D�7�(aQ�E3�8���眷=�q�����j�����Nǌ�_�o4��%P��*�� G�F^�E"O�����%�u���?j�װ	��>`&Z��Y�����B����(&��I9�FjO,�p3?n6Jhh| ������-_1��$�����I=�t�d�����<`/�7����L(�\�@�h��& y�?�B�ߊ��/�'2��~��^3��weU<����^aTw�f�֏h�Zy�`IS����ω>m�]l|�>�	�/Z���d����&�*��P830g�z38�g��Z�؅*�p���:K���p]�Ex�~�?�r�7�ѬA
�}	���yb/
'�+��<Ĳ����P����R��9�*�y���Pw5�����d�ed)h�c{�l���^�F�0��jxFE2�!�s���O��X-^��>��*����ֽ5�D&1	��g�u9I�^���Mn(m��%�j�+�9ڍ�)�7�F:��Pg��Kn�����'Zf|�⯂�qd"�W-�%<�E�h�,�3���~ĩ�."!<b�Q��|+�}� �C�IX�;�հr�����xj<���#�U~�˛�ʋ�T9��ӓ?'�X�w����!k�De.���q������	��}�h��j�R���E�N��w@|E=���}��,c��gQ�l���.3|��	g�mlc�@�$��(M�J�����;�cM�/����c�=VCV���	�h��zopNS*���[<�I��m�gE!���|ӎ�CO���R� �	�Ŏ�@𠟒�e<}{Z�"�DZ�L[�Sw
#�R��5�Xv'�3�R�M�i�Y�]<����U/0�>ߵ��#�?m��ȶ<A���8��?���)��0���;�����k�����O%s>j����T�ϡζ�/FS��,^ta�!:\R��:� �r�o�<���	+By�0�EĔ�T��W#nr��)�,��[��
�NPV�(ή)�`�e�Vo�{zا^�Oc�Ӝ^�台�d
��%�m�h3����LV7����;�ޮGkSO��uCp�鄅�'��f�!ƇMF���� e��X.��t'��`;�s0�\~.S�z8�P�DTW9t4�f<�O��"(�J���;Z �\y���p�u-'>`L�U:�`h�5Q���	��D����n��8��l��/�����v��;jp�>8y��l���Hp�7N��}"�w'PҰ�q��v諁��b�Y���aG<�r��1�D��(�-�=���e�M�T�(v��bm��T(n��_�N�Q��ٺ}�MX}̟�^��޷��^��-F��c(�B�_��~�d��Y3�&$�;����	���1ۇg�� �TM��b�;d�]�ɐ]��X�q�%��vB��d9p']�p/�ps�v._�֧X=��9�ea}<��F�����~ں�cX\R)�݉&PpcG�$���7#�
qs=��1{��AT�z���Lr�O%Q?����sUv��/�>��W����o�wn��~B�I��6 �O���o>;��H�3�u��z2�6i�7�����в��n����چ��X��K��~{O�VZ�$�m*�y���=��Xn��(#`����t h���k"������]�fd���y^ól1�+�/��E��B�?b6(<�P�.���'�D�p�:���X���7v��N����ޢH3���HB\�Xk1�M���p���ٲnF�?0�\��	��u��h����ޛ���%�� �g[��|%`W#l����q��vR�%��H�-`�1�f�+Mv����� 5|.���sJy���U ��Z@#4耆r���3ҷ�FY*�%a�"���h�I�)bZ�Mt=�
6�D8GC3���l\��J=��.�/BU{3��闧j����� ih�H�3G(��i�8ʡI=��Q��c7n���6ɷ)����P&b��y�4S=��.�z�h�������Ƴ��!��+,s6�	$�����&�q�}A=M�g��^�*���������e�[�JF4�~��?^�ΙB3�?�=Vw��>FZ���YqJ|�������@�P��7-���R[M�ŀu�FL+���_����RZ+X��� �����ه^3�� ���DS^R��r�������g-����0��"��WEf�7]3��,��"�����;�1�_�A��U�/��v�҃Q)A�D�;[ts�BҀ�r��R�bC\���b�=�܃T�Gek�%�C芥�m���ۤ���2����l]�Fs�V��uam��f��<�V�+��6�/B
#�8i� kj��x��q��㉑U�_H١_��V�u4���e�rg�ck��,3r2�є9�>Ab��|����I!��J#�pD0��οҚ)Ɗv�bTa�cx٩�m���/����\4fhnZ@�J~�9=.芽	9�dO�}�BQ�wu��n~���Y@�P���[�x�Ab-�r7<w���TU��BY|G�!�U��G�"�Iy��S����نa�p7d�-��çj��x1���].��w���pgj�LQVoSПNي�Ib"��Y�D� F�6N�������e���4>��m�����p¿���i��1�"��6�g�W���1�����&�hV�qY)j�G:���V/U�� �j�3`�0�wJ�V����y���Ed�M��38b*�ɢ��5�X�=a��6�A@�0ű6�V9-�^d�/�3��F���ޫA���i�����|�H�5�b~y����+�w�(��g,�3	����9�|Y�5Ν9Z3�����MK\/#����ݲF�)�H��$�Gs佾7��D��܈�
 ��wj��<%֐���T��6`l�@�� lH��!6^�����~.�	�\$N�����zX��H�L�Ғ������H6��)_p�d���F[x�Њrq�����hY7���V�UU��v�:��V�Tش��Pa�DRY�e#8H�+�"�5|�Y�U�A��@}+�Y?xk`1��Z2>	!���W�C���;�0	r�������g�[t��<_{-nQe�� �� #�Okw��!!׋#֠V�Yf'`g	{�e�^b��JpX�ɘq��������*�!`v:�{�h;\~EF��+,f�b��{_y�}�Qd��{�����P�-�kP|��[��-���UI�i�ɈլѪ�j�K�6f'G����2�,Gl��ʮ{����/-6����3�A�7�-�+<�L�r+��q�׃�39�#b@:u���GKV\H1�e�pR���0u�.B�2ʱ.s&ZhI0����M��늦��vt5*�ْ�)4ּf���p��~l%i��X�9q1w�D�k�����/���G�6ukT�#B��^�.�ieؙ_��0ϭƕ297���>9j9=\���8�[\H�$:�)uf��,2qx���4��/�hח�e�[Wb�_���H52�S��QX.�� ��H�ЖӖ���Ӥ..��3OGc<���a�',�W�rl8��u�hl\!�[�`W�Θ��,�9���_W����"]稯���$ˬ��;�U,ʥs�S�@tf�9�����'Z)@2|���{��8��؋YȲ{�ы�FV]��ò�q�4���a�F
���W�G�ՀVZ����Mo�op3��c)=�Ȓ��;�PЅ�*Xe�پ���>�}j������t׎ 2�O�04\�gh~Q&�L#?��q;%5K��8����5��0Y��nʕ��5itq6���8��N��E��A@��^^�.O�(X�}�<Ƃ�OK����{�����l�j1�x�ҳ@�oɍ�,_�{_�G�>%�w�D��TQ�d��`�	���_���jP��:X���7��A`ٷ�Iz~��.ٗm`ڀUm�@�;/	�fب��o�z-���Z(�1�H�� X�>JĆd��b�T8�z�Ke��m��;`Y~K�^�����DX���dM�^��{v;k��SC�������!�b��>L^;mO�[�5�Z�?8��=}��	+'@&B(������I�*�+	O(p�C�K����H��uXP�I0&QbӴ9��Y������$�!'��!?$LOyԃ?���f]��!(��1�]�H�c�Vq�on�h��;�қ��0X�Q
��{�
��� oa�O���'��������N;�D�b!G+��9i '�KRn@�H�����,����FH�șxx�%^)E�!�j��Xی<JQ?���{�Q�N�G��&K�
���k�oW�r���'!�a�[��$���p,VvJ޴I�y��SL?̈́ehuA>�:�X�U:VH��3h�xm�x�M��N�kR�U(N�s��Bx�KAQ[�>�xC+�dqL�AwGv8��D����ޥ��#���D�h�JM}��:�}�R��N4�El��M�a7
r*�O��j+U��Dؒ��v.8���A(�� \R.�|e<W	'