��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�/Fw��x��b ayk��]���
t����jw-V��k�d<a�f��xx�Zs��t=ߪk���M��N��J]Hd3؀ADw�`��搥�q��mb����/��7��b���]A�=�!VhtJ���`���2�Pf��i�3�b�Gs��̰�O�%^���rH�+:$���U����88s�ډ��R��g�:}��~b�������z:��F�b�YmV���N���u�Q�Զ��o8��y�nL�D>rv��%OC��O*;}�xe5m[�D�+-��j�a��_���`Q��F���F�L��n��Hŀ���(������{ܸ�*�!x��v�Gqc��^�؛t`�|}fV��'8p�!�B�kHd�
�±��x�UU���e�nqB2q�ЙЍ��a������ψ�=U�ٚ�¶�*4l�6��u���Q'�̏ts&:�����l�-��U�5\�Vg�<��0�3aT�h�a��X������±Q\)�cl�e�� �^�a�<ި���9^-|]�	d�$}�¤���#��h3��D��'U��K��r�j Sמ�PM��J+�qz�E�c
��R̈́J��v,U.B�x�{5��-
-���N��bO�������~6�e��M�7f*#�)�,�"lA��PP=�yZ�R)Ѥ�n'=Ur��P	?/�������7�"�IJB��=ib缹v�+���rk���sI���6&��E�A)�_��N��b�x�h�\�ʐ���� G6��#E s��DyT���	��ַ-�Wf��\������8����r��^�`-����y�=6��t�*�Z��?-�~�S�򣑓lA$�%{	/�k6��ՃN��0E=�H��y�Ӆ�O������ۮ���pH)�Ov��W�:�y�؏���۽G��R�"��mva ��_��B��T�C�3VYcG8(���X0;+w�_5��!�%Q:��v��U���أ��Ј�!��5���A�WC�vj�t���|ЇȽ�BD�bGvM\[��1���e-��a�f�Zʙ�B=��F58 �]XgT��k	n{�3Qm�l��]�4!4і0��F���i��:����n>D��!*��U�^���b�W��g�Ay�I����N䆻��&:Y�o��cDq����q?�dIc�v%Ȅ@|4-=j����I։#&���8�Xv���@���>�>/�yd�u�>_3��]����;ɇ��#�|������3:����.T,J�wB{·�����5���ᾖR�e3���N��׬W�B��G���$س�1�Y�B��5a�`02��%�U���Cأ��w	[��8D	��*_�|���	�l+�L&Pa��e L��j���ǘ��!�3�qPn�_��Ӑ+"��wm��<q]��`VX�&曮�ʸu��',}a�,KEh٩�x
4/�C��u{�N����Q�i����"�[!`P�!#�z�!�n% Q�=�6%�$��t9�Ss��ͮ������#��w�fzn���x�=���������C.�g�d]�F(��1Y:�� �ٚ]��l���CEc�r��xi��`��/A0<΍.�r�긏2.�!x�g�A�� צ'��5wh���·BX��
;(=��_Q��c�V��W?��,͔�k�Ǝ���y�K�Q���h1v�=z�Z�������qI��?i�,�VN�s���PI2y��ώ�㪕���N�{���}�f�4aC�Gv�'r�=��,�A��C�,1y�X���鄇��NWFYu�;"hO�����= 	i��K��+�5����o��jV�w]��}��څ��'�t�D'��bi���e3pR�*���gc��Y ��<�}1����W���n�y��Wђd�dop�X+r�p=�̨$˫����D�F��ob#y#�f�~�7t��{d�V�+.���Z�����a�)�x�zƒ�E���C��ػ=��قQh�P �_
���	+]��
���VI�S��7:���۱�{���tZ��=���zt�;��WU���ٶ�)a�`чN�D
�����ǳ&K���m�� ��L�5�V�^�[���/���c�嚄�f�/���ՒwoeV��?]��W�2�л�K�A%�k8qN+Rϟ�k��e����LV�T��l,��D m��Q���\O��;���)�5iq�
�ŗ��I2�z5y8��#�9Σ�1���>s����o龜=i��Yǭ�'�!C��V*~��?TC�;ba����,�E��$<�~��Ы��h���W6[3@�S�晤��� v�̀I��qH�%�qi�����?(E�:�V��_�b�m+�"��=��3bE����\����:]�'�+�,ȥ냽�G�$3����/��g���T<���R�|�xΘj�/����$7i�*'đ��&GV��b�â�{������͍�B�q�inH�BJt[:vI'�a�&]
��7�X���6��A<Y·�j�Yp�~gi�fй�!��)X��H��r<VX�PHןu�E	'6D�6�IV�2��Ú�zD�5��� oO�wV�t���Ԗ�p�f�E3�U�z#��$xB�$Cn�nr�˿R����;LM�▟|p�����3d�7�e3�t����+aYv`�g�W_�~<Y'��tT�7Q&g���ʥ�M*��n�8�7��������I<R�t���5�&y�c������H�%Ѝ�)�ߊ��]��
g�