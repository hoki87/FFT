��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�#&��#�<��������T�]NA��M �\���(�	Bu� �k�A�=���:����V5p�N�=J��s�U#(�W�Iޖ�2�0���d��&����V�3@�&�E ݊O�J�O:0l)W��:@�]*}-�i��P0�3�׀�����8�7:�����= ����6Dg� �K��� ��;K����띫r��3�\]�?}�C $��\�tt�d��8�\>Q������v���3��ڳY�M�=g5%�ħ\��'!�t|S����O��!ɂ5&�}ԍ����r4`���V��΂�V����/�� `�K���|��Ԁ�c�w=�KT,p��M���fzKњ�t������6���sfY&Aj�W�1�Ɣ{�� ��B��p��G��Fbc�Q��mp�hXO��2s0Dl���F��!� �W��D|�s+�Ah�Ng^l$�oVEE���aD�9�F�$��t����Q��X-�}T�YƗ��qً�-�:�N��H���y�qE��R-4��0����8؈AtR�I�g�x\��ZZ �	�*Qn�>3�% .[!��yڡb�(>����� �e:��A]0��D+�@P6A����``�]4!9cLKu�4��3�<!?��Z�+�f�"�8����)�KD���������D�
!pp*�/w5 75R]���u����DZy�1��m��ƢUjz�~��ҟ�����z5U�?��������&��(+��eQ�^�xx"�n��!3�@���Ovy���z�ke��m�u������R��<�%�7�{}}��V�RU�Z����Hc���c����݉�^�	Z��!v�-m��A�<�u7���o��מh������<ic���"�,n�b�-C��	����o����u��AZ���-�nxk���[_	gQtۄ��$ �hԖDUo�w�n������.ϓ��(["P�EeV����Q�#Q�ރK�P�Qt��lJ��C�լ��3N�8�g��h>�<�����J��i'$t<� �����6(�Ȥ�>|�s��K����^�m����g�s���p<t�b*dL�/� �g~z�#7����A9|G[0�M��YB��@.�X#ţ�z�О�Ezȿ#Q$��Q��T�A c�K����T�C����*��p�%w��ZEƚ,p���"���z�c�A\[
W�L�RU9��q��TKr�,4W:ޡ�WA^��|�&c�4G#!NV�͚6����iJ9�}�.���oؼ��gx��$�"��mF��f�Ĝ��g�ȱYo�/����81�>&����6+�'K�r%�xy������Ȭ�&}Ŭ��� E��q��MڧD�i��Hs����8�`K���E�˞��7?���w���kLR.R}LюY��$�H�>	��q����B]���Z����:�̩��I3*�}֒R��2	�|��֔����Q�Y��'AQ��9;���Z�m#��{�S"�mKA9�/����xn�✦k�͆�����C2t�=`/�0�z���b�G�r��b�g���A'@��΃ZiǤ�O��T�YaD�"��
�O�7;(����~+�Ž�5d�P:�� <���<uNŻ�O���u8�?޴�3�:&h7���L}B��$`�M��	Qw3�;0�3U�5�^P�[�*l71��s$�	�޲��].�_e�O�~�^�&� ��g͹}�^A�/�;��e�#�<��A+$�#2ofR��u~���,�_��4S�#�ep��m������ȅhF�����=k�`D���Z�z��yR4�j��Em��g�GN���բ-�7�j}��7s��Xi^�霝1.��\n2}	R9�%���"0��Wz3���u��8�-�^�jS���j@���,�"����e���ߍ�}�F_8�[G� i�ٌ�|���xH����f��1��/@��sI���5zh���>�����+��'eMp�v�f*yPS��dH�S~�L����չB�rbAw���oQ����&�A��V2�wE�� S��F�*y��	N��1�c��3$�Ii#��X����d�1�-�̴Y�19J��.�e��>�JT��q�������<�hߌ[�����n}c��R����)��6���Ԧѽ��Z��-u�C���Ϥ�Ai/���
�g)�+%�'}�"�[d�ۉm��)�Yԩ��.�jk'�հ5�n��%�J �V� U#�~/���:i{ ����ퟳƖN�$���*���ڼ��J�*xNboV�6������]O�68����՛�摕>��~�{)$�	��.!��a�V�6~Q"�iK}y�����%��!�(#�\�Θh\/rHP�/���=kF�N��^���xWb�r��/�z;ʃ��>t�zX�4ұ!�(y�x���t�?�5G�u�>`�=@=�6�9ӱ�����Y*ջ,��h��yL��aU��U��J: �4�U
�V��AR��k`s�-�N����T�3�eq���)��E"}� #Eǟ�l�@zڪ0!,jSF�]�z��I�y��`����oF����DN�'�vϓ�D�h��c�C}%d����ٟo�d̥��, ǋ���"��m+=Z)��ڋ#����g��B�͊�v�2q���YqU�*�����l��Y�0Q*���)}U��-9�VJ�[�8���/�n�?��;�CC㊕��I�|�^���rԺӧ��U!��Q�N����֋���L��ѱe�,Iw�a��|�����̥e]0�Fڮ�C/'j��P��Ĵ@�̸\~�7���.�e6#-�u�QO����ê5nx��\^�{��Q�?�SK�K� +D��07��Ę/��BpC���bji�@6+����"�7�lܥ�uBCc)�����������UAb_
�{kک�klFXW����9�]!&�JM�.�a<�@k4륷��0[�Q�-�Jlk�iA�O�J�}�	U���̤p�F�|��.<�X����'���C�|�8��aɘ���)&�xG��c��~q��z6�֍��T��-d%���=*@q.l
���zWS�<2I�;% �u�X��f�ඎ�gv�v�Э�j��n�����D�Pp�]��ϊc��5s�"`d@b��w����Tb� 9�i\��k\qtg$�oY<�����=��1&x5ծC����r�2ܸj˧�;�x���b�CG�+h#��˜?P@(�
�sp��Xl/c���m���J�`eLe�B�С��K�gy3
�͂�}�X#UAB��e��x�7�����`�q�g�W�-�1y�;����t��m�!�6��J}��=����WZ�!�$tr#