��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ����������]w���>���[���r��7g
�1\����x��D���Ñ�m��E�8p|�(I�҉��Dw����ɔ�{��j�:znJ�2�t(Ǘ`t'�DVu���0Fm���q��vL�_�_�L�k�Ƴy�2��>���� �|`��Y-��w�v@tb	Væ�p���o=��V�w���[�qQ�}P�w��X��aV~���_��@8��ةA����,�Ļ'ON<���X�'8|Ӹ��c�0*O�מ
��[�ZT�����A2|1���B����xux�Y$���9��{!�[Y�&�aO�H�n)�o����mp�n�P��@��*�g�h�^�ǫm�@��� �����O>����̜��m� �x��"��̖ԖV���}��6�'�<�=LIY�g�X-^�~l�g)�f�)}ݪ�#e��]���)���1�-��G5���ɹ�Q��3}�����&�3��O�?�-3��A�7�|�
��Հ2Ǩ��Y�$�.��8X^���4B6_7�~QU@��� <sW �w��9��+3F�&�S�Ar��t���xR�;d���p��y��w��9�ЈU=h�\��R�,�4�l-@�B�
D(����\��%w'S	Ш�D�UW��V5�%/>
�����pܔ>E��gJv�q�jv��WQ�TA�a�EV̑|��T��*)<'Kh�iz\F�(	C�k_�FX<kn�-UV�C���՜8�%�~���zd�U��-�әN��M�对�8O��y���B3�
a�0#si6/y�:�@����Nt�X��K.�VTy|vPpk2 V#��7#l#.�{`~5�SD�G��ZZ���j�My�Eۖ�v��Ɏ��)�N��%��O�\�w�a�ز���It�N)y�L_���ShQ���>�[1#�M���2u�
�����2�̔'r�oq��)1��B��yF��O�c\2ŀgyBf������~�e_Z5������A듽���#2B�ro�g*����eH��gb�L<ײQ��aYL7����1Z�)
J��\�%��Uz���yn�7�	��!#\&9�W�萛��|Gq@�z���pX��5���
C�(zB�|}��p���ʽ7��a���8\��mDa��B������q�k���'���w�;_�}g���$�����%���]�X�m�5@�� [Ԏ9DX�6z����v�I��;�e����D����i-�%p���miE���є�����0ad�s�sp	ҹ�ڜ�uWg��@�<����C��������+)���<���ЎW�����݌���HD��x��#��uܐ�$Y&^��������k�|Z��V]�`�,r��^]����(�e�\��B��z6�u|>�qY��+�,]�����ߗ.����
w�f�4p��ra�2n�A�/Y�i�� W��?V�<��M9oc��٪����պa�l�%���?��B%Cn~y��8x��S��꤭_:���Ì�?5����e!.E� )���&itum��{�#�^��>�'{�7z�{;r�+n)�񠕍�|l[S���U�+����>=�I�h��@���o�"c]e$�o�?N�\�c�3���a8��ۆ�ƽ�3ۤ���n�Z�������Y憎�����q��Q��כ��J��e�42 �I�=D��<�TJ"W$o���+������w��D��\k2S7@T׋I��s��J�䐟x�E"��gM>�M��P��`��䀇�'M�|�假�� "���V�����Z��;�լ��$�*҆����u��?G����5����=�ؓ��z6���N��m��%4�a�*��0�F�f��q�j�����Z$9-�Zu�ױp�?f�C�C6k������xܵ0����#��:�?<�}��>�[X�g^4�����6l��t�J�0���H��v��g)�V�:�X�˸�.@�f�w���
CK�e�Q�7���s�f�m�C�$i�6������u����<^�ᤒT�v���R��s2�)aq����q��[Q��������%��z��?�ǉ-��L��p��eY87�k�`'e�~��>F�u�/װCO��q���|#9�p<O�`nW1�����UJ�]��dݺ��뇐��Z������7�d2rz)��h.������E|T�����M^��Þ���3N��O��س��b�f�e��M�Rt��ג(����Nq�kYY�����;����Q\����[9�[�a�t��7-����d�MO��tA�%��8>��0���ҝp�{~���0����PꃗH)Yӹ�w��x�$���xh׺$�f8f���^>n��H��@��i\@�9��[ƬptXp7�Q���s���vצ2' ���U�c]��H'�� T�%��AMX:�Uh�0k�v�M+��
w��f��[^j&��!h�a�P�c�����Wn,M�o�D���1\~5L���<9.�cErմg�`u�&#�̞.�Np�t.qrݎ���z��۫&�b쫶���|�>xK3�"Lfm�Jw�zІ���S�z�"B��oq��k��<GVg
5���,���|JI��� S"8 ������!PV��-�:y���S-n)��:�LB����GQz�`dZ��NQ�t����/����ti՘0�}��tTX���W� ����[���6˞�h�eMi��ol�i��KE�E	P�$��S�$#P#��E?C��}o�?�9r�I��-u�F2�%���~_�_b=�CC�� �F��V�9ppӽ�/����%���X�����I#�����q�`KS=d�����-'З�O!�$�*�Zްd
3�!Pݑ��,��P��$�kc��3�m2E�� �B���A��*Ir.[R���1��D�C@�����<���j�Kա����<Iw�4숯�AW�C����5��Vͷ���Z��h��8���}�+Ţ�HK�5`��yD�i`U��7���!eT�2߼f9I�p��G�ѳ��
2��<6�[MtQS�7(eD��(п4ǖ%��Jq��'�,�5���
�/(����d����\���؞�tV�����K�T��a|`�3����=�ӟ���mҐ�s`�y'�s�"6�I��Gf��tY4��c�O	晒��Z��PG�%@�4�
�I�sZ���I"0b����Ұg�����z�"��PW��a9	ա1��KࡴN�����"�'��Yt���մ0x��=<���5���5����o�Cc	���i�`���!�Ȕ{<�DQَO��v��p���^,����WM���Chw������4 ��?�e�t22
�5�Z B��h�T��9���	#���]>[�)���-��t��`)��sS�����+���A�M���T�k���Nڞq�3����ͅ��-�
g�s ��+������ ����j�/r*�~}7�Xy���z���0�:��bbNd�7�\�H�6ݟ����qN�A�y5��]݈�{4������G�L���"��7���o<B��C+굻d%����N�y#p���[�
�.��m-�t������.tLt�5Ő��B]m�̝C��T���Z	lp�r�r$�'�
�?O�/�j��AY,��]� ��HO�I�9g�Q���'T���A�Fx"�PTnb�d���B�����<I�+ǫ6>��uv���h(�^=��R��6��O^�����(��-�L�/Ib�%r^��$_�kҞ��~�����a��_�W�tn7�
��Y�L���.�n��tu��4P|-1��x�ȬG�o�DҨ�}[H\��E��n�9���+5~Aj��3)�ׯ���c����Cz�~��.�=|���Q7�b	b�e���,��@N_N'�.:�_�u��J
o1����f��꽹9ޏ1���hB<����������(���n}���Qh��~;UK�����7�k ��$kϫxP�D�_�MF��M U,G��]���+���_���) i�"��o���~��1����Da
�7��q-���n~�3��F��%��l͂�\��C|]'�Eɹ&��ZV ���ٳ��h1#�:���Nv �E�@�G�uqd���(��փ�b�4�I���	E�ؽx�'�$�y�Ku#x���{Jik����Y�1��Jɭ�ipgVA�0t]�T�?�Y �Sc��<>V�m<�[k�.}��&s������(;�gp�g���gh��'�<&������Ro����j��å*�A�~�k�cg�W$�^��� ��<�c3����y�]�\�����z/R�h��!�N_��nfi.���̟�7���(xO�M��1��u�#{��rϲַ��Q���h���^����qm���c�]��)Ղ�6��}�ϥT��°� }+�_1@>���?Gӵ�P��{�iiʚ?�F�s�n���F񌏧(���&�$j$�6҂M�If�����[q��O@L���g�ɫy@^ͺ��M��3��5�E���i�4b�P�dm3ޭ=����y.-ϱ'ו*o�sns��]|��������g1�Hty���\�y�Wh��Ë)���8����Qk�^�X�g�AV��,=Jf_�����_�Zc�"Q��Ä6?C�1ε"���',�^~��<p�TЛae4�|oı�q#�����q�T ��R��|�^�&s�%��eŉ��Q��KRU��EfH��m����9_��?$c''8��m��վ̳�/iײ![$���f�����'7��9f�vHē"�x��U����m`r���u"?E&7��b�\��t_�|_�Ǫ��yE��ohVvp�"�͝}�n�xO����2!I�y����y�d���f��ڷz�ej�Pxl��+V�Ǿ���{��CJ�b�Qc�Ӌ�T�P��lw]��#h�s��eվ�s��c���J/@N��v�(
�t=u���eW����}E(/%}�ġ*V�?N�|�|Φ�DY�u��s!��v��{l��J�������i�Z>3�YziKp��
������N��c��tA�,�w��v��6]�ԑ%�j\1��]W�%;a����\��)�ާ��*i�Ay=e��m8ə�Ϋ>���}9��^k��_��(he�J��g��B�!�%���Ǎz�;|[���PڐI����}G�� ˏ�����p��h��b�j�׸��>i�&O�5U�?�b
Ͻ��ܚ��K�\�@��Z�$�e�(�3��x�}����N�❲�\�\��������[����BdN�e$�7�6�`1��M�5M�m�� 5�KrMM5Hn�32	������v�	�R5��H���20�M�@�!�bs�z�^�)�6�h�X����JL+�y�}��O�sgL���]Y��}�B2�╺u�p�X?Ę*Ȅ+�Ʋ3PM6����Q%u���8�[W�Ԅ�;� �8^��RUf8�����B_c:PK1��b/4�cb�N��"�H�@c�I'�r�h��{�'��n3-^�l�����7XUҎG����6[!C?b�����N�ί�[��,��U�&M	�/Ղ^�B��
]M ��b"��U��J)\̯��Ҷ���3��r� ��x,Xs1b�	�8b��M	��K�3Q�/Rk�%��#R��o������"��n����7�HkY�WK����X���i
�x��K��R��9����^(��?[���$}�a1����S|x��DPa��.+�ގRˀX�<��X� ��f�Q�%�ә��J�C�d`����m}��9[ٵ�[�Ǫ�w�"~Kp�1�N6���1�U����7M;т�a�*S��u�sR�
(���{�#SӒ�,s�i#u
�Fcq�2X�Q3��
(���k��AK� �&�;�}4>���Ӛ~%����XV�
�+8�%T֝T�>��+��桄`y%��Q�*\����:.��0<����
2��%���
��=�	��y;}��s�o�Yʹ��m]M�F�H�3;�� ��-q%\y�?3��>XV���7�c��w+C�Ja~a��8dM�_��H���9����6 �(;&�ӕ{Xgč�A�x�ۄ^P�N;"�	�K�Nֹ|ߏ�l7��j�1L,"�n�yE���^�2��^A�}��5��3�$��w�,�e�(�����%9D�:���s*T@y�4L����Z7S��\�����~뇭�Δ��T%��a�`����4oM	č�٧�f�r��x]b�jBlڌ��U��ї�EZ{+�Z�9�M�(�=HAe»�N"�ڒ�|Ռ����fO��.=��s��vӅT\��YB��^*� ��)q��`m�Z
����ɝ<����Ш�J��G���&�d7��2�c��z�-����}i����&�J�猃Ĩ��W�2��Y��l9�w�%���yY���[TY\}_�d�Xk�����<����3bC�Hj��u��A�p�I�j�]�Y��i���7�^w�8���tu]�����|�2��r�m7TF"Ϻ�Z!���uRg�.̤l��[N:��eZ�ߩ
�`�;%)�ɍ�a1�S�xy3��;�<�����C��:�@1"1A�W�FE�p��'�Q�� ������M�?���קs�=M��$'L�y�~&�)6W��e|8�a@`�u%��KP��R��<�W����\mQZq����$e"<�C'ӳ�N5b����j|��F�>b�s	QD$�^��|�]�D�f�B�9�͚͆��)���I�,NiM:FT&��{���
�զ�^h�1�~����f�7}�[���m��I�k���q>ƶ�d�`�wb.L��g�W�q�բ��`�J�P���a�|�;d�� ���8�����c�Zs�"I�X^�CS/%2�?t��f^�0j\��,f=;������d�3�`��]��ꄎ�-Q����Fo��3: v��s�0x���4�Z��ӂ��}"������Q�-~��~~�-˙�p�r�T�jp�yH�&(L�����<�Z�"��>7��Nt�F������o麰�m�UL��r�ECƋ�(���T����V�^��৪2������G�.��i6�O�!�f�����L|�6&t�ElpdGh_锿ư��a|��ؘ�|������ �3t�sۿԮu�]Ȫ��Aoo)��P��:MP�9N��*Q��u��\@Qt����	�K�W���!w�jy=�X^ ������4�Bc�-�c��^�e�x $b�&�3w� �yn+��0[�&��D#@N 8��D0z�4T�@ɫܜ(h# ���x3)�P���0��û��@/��<D�W��k�'3�'�J;�%�r��tl2K*e0���)�����6bc��b˔���2Z�uD��v%���f��0� f0��)���]���{�8Ɔ@����R9�������@�Y}�W��V�4�W��$0p���j�ثM*����5ȝ�_~#�֫R��F�G=��OQS���ێ��R{,�?4��b���tk��LCf}���������X�"vg��r��"�e<n�R_���/� ��V;]��E�U�-G�ZvtkHz��a�"�ĩn�1�{[4��i�1��ND��Ǜ8q](�N -��-�
��fk�Z>����{k,(�X
&Ցn3�^,��^�B��+�����«!�b ��(rsaK̥���z�˪�oϡt`��i�d;�i��u����j�f�Ⱦ�Fm7�*i7�O~,i������	4mU��dR4����+il��z@�ؒ��5e-��Ҝ7e�k؋<ZW8<�;W�	��f�a�%Jw͸���1Ti�[V��v|㞢W�v��!�]�H ����W�K�Q���?>Q�.4��\�˷{�pޔ|a���Yq�VǤ���,����F\�9}�k��zZEdkg^�+����p���]�1F�8^N)_���Z/���W��N[��q�	���+-�cZ����w��ŉ%�C0�^�.�����7�	d�p�7�^�6�P���ng��>\�ޡ�쬰&E�!�^��R�|M��'R3D螷�|q�uq� ��"K�(�� ����e�݉�1�$�MjZ��鷄5ՠ����9��TS	 � �1ͳ!�Ќ�&�C��w��� o*#/���w��u��q@ `��a��Jq��Agz�ͷ���D� l�F�~��9is�~����.�����EJ�T�x��y[U��=�$����3�I� ~p��1B!������`!�
�d��聽�������;�	6�x3@*���S$���ǃ[�'�?�����]�ꃹ��qG���@�^�w��x"�d~���o�oi�lV&jze�h� �9�T/�!��mB�k�y�7|n���t#^?{�b�"���,��7)�D��x�gޘn\;�VW��a�k��"��q^i��*s�A�F�£�����0��rl:��GpWh���
,i�Ӌ�"��#�?�U���D+�2�&������Z��$9Pnj�$u�S��K�B&,q.��4,���e�K3��������\�=H�w9���9u�&Wr+_y�0u�.͗�9�_E0���{�|l
E K7��$ľ�s���\�@C�4)��]ҋ �n�����,>�ާ��74��@'W���zɊ���3?�	f���(�D�%yPE%��\p_x��ŗ2���c�YP)fd/���	�bH/���T��!^D!���7 y4`��[��vh���gYŌ'�se ZK��)��