��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�#&��#�<�����ﾍ ~��ąo��L�N`�	?|�,�r��iYHڞ�T�/�[���uİT��j�	Q߿��pa��zxX�Ӥ�T��H_ދ&-\�V
���l$U{wص����F�>ܼǯ�HW~"~f5U����s[���:d����6�Gˉ�I�3��,C�w�{J�}�XjQ֓rz"M�<�B���Y[�������1K��w;�+���t?�B���7�y�S���J�<%8vʱ�N�n��m:c��-p<�5�����*���^�|�4ζ�Ab����µ>o&�L�_#�~�{fQR-���i���d��G�����Moy:�P����`|�S�ֲVV����wΛ�KGW��=��(��-!�I����oo�����4Z�-�.��A���>�+��V�)�[�v��l��������b�h�_�$E�3g�[�]��IH���ΎqL���ys���yW�vI������j���.&�4�A'!��X�G�� ��bQ��`B�2׻�tJe�������P���.mk=�5t� ����ipq���x�o]nו��"���/N�}�SR���<:�?��l��?v�r(�w��:��16LeϝG� ��.�Y�#��H�Z߿�=P�E�m��xQTd��;Mt�.�D�=y��Z����<�/#�S��	���g��_[z�}�2��TR�TB��_�뚗�~���1d^դ��	A`$
��b�M,�[�U"����9,�%ɴ���N>{ìMo%����P�HA��
<2R:Ժ���ۥi�|��0NqDVւxmIk��R�r}�n��4�V\VOX,~��"K��3�'G8��&6��d�6�ه�he�>1��<�/���sh��P��P�mՠ(3�L�V/���S��%wPU�f�~��*�MVw::�K���dP��'QԼ'd��,S&���[�3��� 4��*8u����u�����J����*5��Hۏ<�XbQp�T�x�����{�ш�<����$F잌p�]�Vr\�i��`=B�u��+UT�J{j���c���=1Gl�oO���k�X�� ���m;�"�T2t��������]b�I^mA��ō+5�q`�)��Sj ^#�~�����o�3ePmYu��7���\2 ӵm;��P�G���W=�,j�)ao���#�#�pK��#@��=�}��>Js���.�.ܗ��	���_w$K�\1�J7/G���/l�dk$ckަ�n՟��Hˆ���$ �p!���PM�GjjE����)$5I�X�A���	�v\�SE�[M�j���`�&�s�T�28���j�u�
1W���>&,-7фo(�
&�wO����#>�:�Ŏy�ծ*��m���8�� ��[�[l���o�Pc�E �X��Yq�#e֎ [��k!;5/��/B7�N5/ꔰ<��M���{��lI�����{���?e:��@N��_֮�� ���1�T�p��4O��T��Yz�Kh��ه��n�4�0��,(#��.��´�u��O���R<��V�J�w0�^3�c�wo	�ʎN�^6dϢYC�(�-�3�*�`
�����b��� ��	���U�S�%�ݯ��	�;�����{����W���)zJ�~�:����Q~�و9OA7�<P��N��RyX�1%ٗZ�Wv�k�h���w?�|~�L�����t���U&���I���E�>��x��1���x�p=�����y1�K���\�U�'q�ːΆ�:JC�]�^u�>�Đ��h�8E�%��B��;�U��l��6	�3�?'6��B��\�.TE?���c;Ƙ��͡_o�����UM@ܫ����
�����c&I�0*�HXp���=�V�,Ț��z�q���j^
�%��@�nu�E:�!(H�dH�=(�XD^�Usr��Hg8����qb���k�Jk�� �?2E�fz����������w�B�M�9E�Y�%�}�j���u�����+ԯS�/C����ᰳ���a�N�b�Z�����סLx��A4E�������:2���� �$q�����z8:�1�Gc�,��/�Й�&���Av�pLs�1{�*��uဥ������? h��z^{l��=xU��)A��&��Fv��X�y���D���	Ҍ#'n^0� c�~��f�z�9Ѝ}S;
�+�?����}tl��4T��wx���ޑ�$h�d���W�*�j)�7�j���4�]�%'��1Xr�yI���� � q�'oI#g�)�5�l!l�fh��$,��b�Y�`�5�\;��K ��Q�Ν7Z;���~0j�]ֲ�Cg�jcjTB�Tcڍ�..9u�O�_1���E#�M4/v�
El3�Gt��,9Q���%-h���Z���_�����ْg�A:;0�����bu�2��F#wt!!#m����Hm�O��!1��b���8���%��Pfp�Hӑh��!-%"��y�"�y�Sy�̄U�?���-5�4��A8c�����4GmT��w/���n�t�~��Ԁ!�zoM.���$V)�f�j���#�,��!�����KF:r���L:�kC�22b�X���|d$���7��o�`��Sb���<��0F+��T����>{*�2�����.h���u����z��/���M�X�U	��!��7ׯ���H?�t�(�%�?�l1���
���s9�K����/�1�V�CJ4B���?���f���3^~�dBi������}�Hɂ}�=�-�㨜��.�$.�v8D��j�������9g�#4���V(h㿜`���G�W�7չ�7�[�l'1�;�q�b��LcGΔ>*����G�[�q�Hc�:U��]k���H@%�ю8�|J�O���_���CBk�m#®+�i'���ZB�6FN����p����y��}PLF�����s	T��A��E��R�`�5�{���t�6�Q�lox�N�Y_2�Ȭ>�6ND��cn�����b�a�ν=�~V3$�V�N��ܠ��h�j1;���4��<S�_�e6J�f�	�0C��*3�6P���,vYov�@�Nof�H��l���ᴍ)*Lԙ6�z�����Q[G�ڇ.'t���m�T��g+ii���>1t�zd�<��1��b�b��.�k㛼+ʲb��y�`�x����3�u�d*��oiҫ+y�����jxa�D���z�4��v�?�PR��|Ji�*ع���l@X��l����ؐ8Z��ю��R�ֹ�0�X��&�!B�ۚW����T��?�4-�3H(?6l��(�Zn;ӑ��ʟ	��QjuA�Y�K��S�������]�#v�F�:��!��[1�q���?�^_��m���jR���X�R�<�>�#���S�tCd�Zʍ�j�Ϊ�%��Q�����[���lMG4a.�.M�f��Ă��V�LnBe�C���u
y `��>o�1�>	d�(�$X4_��+�x+�8K�#�`�oȣ���=�es�Jf,WOk����N�,N�r��t�"��#�R����_A�@���:j8�})$"���c~6�?;>R1�Iݮ t��shOx�1a%�1S�x�D�U�Ùh~_�:�\Ƹ$�Bk[�f4���}O��V�R��徜�[`٬�ѱ���Wh$�$� z����ѵ=�>w࢟Z�c6d���z	��7������s�(�L��'QK	9E��������hw7���@�d�8d�<��RGIV2Zb	2��oљ���ޮVm�I1#MQ*l:���] ��K�����^�_2�w�c��i�Q?�\`Ql:غǱ���_k�-|�vg�g�7��4��#Eo�L[����Hу��p��_>��qZ"}!;8��S����z�.���F�)����!A�W o�'�}Ȉ�:w5+�k����hޚ��[
߷�o�4�YV}o��[������m�����Y��Dy�ޒ���� u��q��1�T�=��"N-�=fihȷ�N�b�T3���f4�$�O��,�q�J�,AHy|}3��iW�Q�l�ty��O/�Qp%�Z�����؃Hm�NA�E-ܦI$rV[�`�U�?a����M���K�V����8�"�������)�U�48ԥ�M�5��w:U�"ϒv�)�� �>�m�J��C�1 3�ۖ3��ft��=��P��U���|����<V�V���
�3�1ز"�LEm���16�j/"A�1`b1Y$��L�����P+��O�5��
�u�K�ө>��[�y���8o�3NuP����zx���'(�,m�r�N���twm�:ƻ�d�LJY_��<�^-�|q��ڵ�3�Bsq݆D�.:�<���6Z��81R,b�+ԛ����R����+i����ؙI�Kp��{�k��AK4�V?�b�ѣLϳP�b�I�=�CG�`��3oʤ+����|`N�e�J�Ǆbm�D�j��D��WXBUu`��g�!��(-�Est@���{ֲ�Y'�a�i���ƻ�'nX����o�\��_ �S-m�3��=�&�%� ��S�,�FH\`�����wuq6:?k��Je`+�ȃ��R�� `!nA�GӼ���!��P&�����A�&X���5щ��Na���LRXT�:#�B�!�E���mɊ�QCw�x��ߋ�D`�D����L�$mD�Z��8�<�e�M���p8���c��7OV^+��'O���=�;*v��0/bR�\���A�4?=��?�+j�k���2f��,�UF�;n
U$����DU
�'����?z�H��2�s�Y�hn�;^���:�;��t56�Hq��ԛ���B�9�G����c����p١�"H'wEɯ�(�|�du���_��[�����i0 ��9CS�G�0�D��(<��OіN�e9:Y�U������>$�t����������V�,�|��R~
j  ��3����l��lG5&��&,��=�zM��CRz�j���7Sgl�)��U=�V�®�;|?!��ʆ­'�+U�u���jZt��by�����У� 0���>�4�|f���~�Xk���؋�6Cl�G�A1��HxQ&��X 1�.��F�h����c�d�z���A!��"ul*<v���Jk-L����!���:�ҕ�a��>2��z����O��"�ᕓ�΅�����D5k�̫��5c�>��ГW��0��O9��czW�o�m�y(*�WG�p��H����t:��B��̉wiq���q��W��+ݔ�iw�~U͑�6uVk�C����s�	��(`H�9���~�T�B2a�t��N��d�;��~�
���-A٭�y������S�P+��%8D�򣵨(F[�����׬Hr�Z�/s�.�I�pp�Q�<L�1�H�S�k=?E������⟺ِ�ƛp� `���.Rl_��t��y��XK�+�������&X�����;�=�z�L{�W9��YR��B�W�t�&Y��24�,mU�&�l=��62��'ߞO�N�I�®��k�<��S��0�s�
�rQA��ω�����4e�3R�l���D�ZX��;���Є�
��1�;�ߜ�3�l�#uhP�#�S�l A�+�NM�Tr��� ����l7�9�gW�˻����}�Ad#���$�������}�Q���HW>�ԓ}R���l�,0�W�v�Õ饜�_������aqh�'���^���� �ۇN���h)��_���I�:	-��&�P��橗ƶfW�"*AYG��5��p�f�3�n Gޘ��[ 3�DHc�����J
���{�ɑ�Yu�nH���B��w�EF�3�m/��UgA!�����_D�$؏�o�Fzc�D%[�k�S��j)�O�3����ϥ��
lۺ-��h 3&NL�r=w��~�©H��]���o�et�@m���&��F^��J�捤/�G9�cXn�9�K�>����q2Hن'�+�Szd ?�/�צ?�2�΃���a�e����k��I�z�w+�HU1�� FHwu K���^���9K����V�G�����	�2O�|�]tT��<H�xAԞ�NX?{w�X��ɳ��!=)�jS��/��,��-_m8���ņ �P-���"��*���S�Ng򜩭���/B%Y�Mղ�_���⦎e�X�5w��G�M�=Fۗ�v�Ώ��`r	͜�%,Ʊ.yA~Fc/��\X��7���O��sPm�%��t�֜�,�������qM%�w�BWbb�L�ģp>a]Ĭ�	 �F��Y��p�i&jI\�p��Uw�t��B��|[y>�D�#��U��1�«+lx�vP�0�^zt���
�x*��z��a��\�RY��_Tʔ��6�)�"26'�*�j����]��w���=Ux�b	�y���@Nm$�B��N^88c�wQ���Z-A�t�
��q�����񩳾�Fk06��h\��Ք���<Xf��j�J��>�t]��0-�U'䍡��f���L��w_���\	��OV{�h�X�N�6~�E}8o��N�]��륐�#$hI"D�P�Y�C2�2� ����7vy�dU-o]��y�ʐ�˅>�3���C,�/���V$� .2��+z�\C/����n��uF�6 P�x+�����ZǙ���ゅ(�����E���:�
�z��0R���( &Hg}͊X��o��6����l3�?��-�Y �*IN�w�tN��z��N��n)�kk#%G��
����! �a�maI~��)C� {�L�<5���#!rż0i���F�)#Sl�q�T��n�����n�l��I}�Mt������k�m��{D	b~��Ћi���� �4������S�ĠW�K�n��:i��'��;5(�C�$�D0y���m��#��lLaĒ�1i��JCP���P��ݝj>(����F��t4IO�u%����Z�Gu"�+� /K� Ț^�IF{�;�fx��@�XKW�;-2Lc��ߎ }�KY���R�LGy|� z�H�-����9��E��S��Q���
\�%�m<Fј=�;�iG`@�����yt%������K���c-���1�����mK�w)���-엪�ʢ�����j�'#�90�㢭׸0DU4���qt�Hr~�N��5ٹX��aRr/���Z
��,Yb8��"�@���J���=�m�x�~%+Y�~����]eM��?�zR�?#�$!�8���?��D����h!��b�~����O�q��bփQ�l}$��)���B�ev>s��i8q�Ƥ�E ݂f7�P�H$����醕��8Ԓ��K_ӓ��=������J�r�)��F=ҧ(�Q[��ڀ�z[�4�P��B��3u�`"��Σ��!t[�K�4^�i�h�� �7;��L>��	Y��P���Y�{@�}�+��b��W8�>��*�F�8�����87m��
���[P�K�t�go�ʿ*����Kf�ӻ�!k2{�~��V�ej���JJ�xS�A!��Ld{�{؅�G�����*/�16��҉@T�T����z�=���u�1u2Lhr��WB�I�qo����~�h�������l���Cn��\_	�$��7�zM	bL�S $F�a�k�<����0W-}ӡ��b�A$E��i-����.!�s�u�C��FZү�~�v�bW�O,`�Q��+
<�4�veH�/(���"�E1�dI�.����CP��9P�0Q樱C�������r����{���>��Z"E�?R��S!b��l%C��6�V���L����Ҡ�Ճ
�{�ꭝ�!�R�����<E�~�Za������c�dز��+"��/P�Oxl؛P����;�)�i�l���	�����L�hq��}��Vf�Y�ڳh�Eس�	87�A�4���\)@�T��N��"�ҺU����ȅ�����@AT_A�+)��!��d����~�ٳ�q����c�`4����Kp��6y���Kj��s��V�?*zš��zz&1�	�V!�����%!��*�^�nyT8�k�Wwj3��Ε���)�Zrш���6ٱ��ʿE"5,@��.L�U"��qS?��j���J��>��`�^�vʰ0髒-;\o))2+�/����d������uHNf����4�N�+YU���T���޵��~���grb'dI"�w��$�}@����ު%��TL����KD�֦�[*l�<A��%�U���^k�NF�ۙ7K��Kl�v�eB�!M@=��+��W�Tl=�����#�{4� �/�Y/��g��/�ǅC 6�KyjS��%|c�g1��-]a��Qz����|�R�dg��A<�;Q�(�>�W`����$�j�y�q���?g��7�jא'��|���1=� �[�����o�6��/�^�IB��ʰe;��ؘ�c����WY7��b���Am�j��G��&#?k�e�v�2ȥ9��<�R���\,T�>�p�|�!]�[$��c�JVH�R]�-�C�x����$pw�����i?��d=�ء� J��z�s/�5d�fY>"���÷,2����0��N�ڛ3U�(��d�#.�0F�C!Kr<��䇶Q���x�(4.������5��k��C�K��PR�ԫ�g��6 ��Y�8f{�b�D�� ��*u�kC�J�P��pW]��1��ct�
L �N�8��雍���p7{�S�8"��Q��)2����u��d�F$��R(�'g^��S��#�k�����_�l��S�!x���V4/�����vJ-��8�H:)3=[M��T��%���XS�,bD�5W��I�O����~9;�.x���M�|+��k=~����{+%7�L�
G{G��+%)+5�'�������ߛo�?�������`E�3���J����z��j�hG3�����u�U�u&c��.X�ɥ�wd��p���`�dF?T��"���0E�/�_/�P�G�;�4���u�ikKr�8Z=�5��:O�$�r��
��d:�r4>��2^��s����ؽ�8�1�{�J�*b��}�r�Uz��2pBE�@��k�ݝ4�W�{����G����KE�n�֐�)��W4ڍ��3j��Ҙ�p�R���~�3��>��@�pO'��,��s�Qq+#�@�8��B��Ylw���0l���P@���ƥ)��b��e�s_������ T�1ݪ���S�9�݈F�'�����Q��a��>I<�����*YBA��Ί0(�D��E,�L��D����a��]X8��O�w��i׵wb���!�p�}�M[��N��Os��6��Q?(F�q�ڵtg]yP�s�~���b�̀r>`��W����*��3#����A�/27���1����wX�kŹ����N���<9�tIT�Q�'})��DyѾ��ǌcG�����n���ՖL���8�
1�����=��d��!�c�����8��m7��\�T�%Uߓ{AF�0G��������r�?o��Lo�j1 6��k7<���|RP,]B�nV�`�w'�S��Ny2G5�zY=�z�*�Z=+��&�>- �c�䔯=�3�oAX�˽�ݨ��Ctδ�%�<��T�dٜ�#g�s�?��"d"Gk�IpŚ{�c��qQ�|Q�2^^�ؖ�g��K,E�pn�����`���+u����R���U ��*�� ��s�M����T��t�j�+���v՝���R�M"K؉s��]탣=-�{�gC����#��;G��w�v�v�h��Jyw;d��3VuC�h��q:N�h�lܧV��c^9��G&�l���5�C�YA�B3	5�&263��_��E�6��#�j%2�#?Z"����zOf�طt�WAռ�f�MZ�n�u�Ksop]�8��
D��<��c^C���00+��@2E��U)���ę�a|w.w)��.��DS ]u�S��Dc?���Vt��lJC�T�Ԛ�ܢZ��i�����oM��r}�nzn��������}I�,c�&���:�A9�*���& #f5�h3*��[ ��?s�����������-���"6�}Me�]����b��w�jL�yٝ��1�)qk��d}�f�M������͘���t��+�5T�-�p6�+�^��vI���]�6EZ��XG�zO�,��~Udav.v����Q��V4|J�ܣn1�KK�}U���`��d��xh_�@TO�n4��lUФ/�g�EU�@���2�x
�L����DX�"������2��G��uWѺ��-'�:5]bҊ�M��Rx(�?�ɥ��v�-]���T���ئkK��XZ�'ϫ_�m�7�<����A.O�ȡ l�]��#_�V�`ڥ�!�܈�a뷚4#kA�wi6['t�,	�ץ+���O:�=� �Y�n��}��I�p��x^�>W�Mg!f�	�qd��H)�8O�/~��t���hM������3T瞷0S��d���%�JFyd�K�|��ky0/��&,���v�{�X��)�Xh4��D/>����z�Ҋ���ƞ%��7�p�e�}Yʁ���!�7}�/��F]]��qu0� ���͸�����g=As�˫Ut�dq�ֳ�ѳIN�-��M��]��7@?n�Q���̢T��jzؗ&���W�x�~L"��)��̵o��i���k�:��-u,FE[��|u�c��f;�����N�y�l�+,������Xkc�|�9�S}\
S*����-�=w�a_��Z�Y0P���Z��+��R1)���6P�ebÒI���S��(��	�'���b��\�?� $�G�����o-j�qZ1��ŉ�(փ 7��h�u�轼)�S���ߊ���Y):˰��O����4t��載����ْH�-���]~*���颯��C�x�h���sU7h�C9_)��p���g� �fM��Bk���xN��v�{{�+��[�e�V�;j��a[��z�5��i=���Q�?p��:�1�{ϒ7E�3�Z	�B���t�
S���lr����Tt��5�)�ļh�D����o�[V�t���y57�}{��*�O�mU%�)�_�w_��(30���j�E�zn�ׇE��ւ�%�q�9M�L���G|h��BW!V��]u:L���,IK�_a�c�l}P�2�ܵ�ލTI���ɾ�Ī!�@�� ��|�
��F#�1y�@��5Ӂr�VM85Pԗ��J���L/6���O���9��</��ڑ*��4��l	�tNG�^_�p��(���q��nQ5@;�� �)UE4���͟U�H�yu���[|���`�c��w��`3��SZ����t��%1^E(��E�FK��Մ����~O:T�C�)?��I���F�y<�0�Y�?L�B,64�.��j�͏i/C�=��tC�����C��&5��D����D�@QX%����g�t�h��|�`5�{k���3MH��>���C���U�� i��b.����{��L�;L���Y��=���<)�P>4��9�R���fS��s�0�g��ߟ7��z�u�k*.�+��˩���t�`�Px$�i��\�[��a����n �p��ͺH�t?���-TP\�	{��n�z��Ͻܘ���̇L��kC��L��Q��g�L{��1�3l������1����na�A�j���G�D9PJe0~��^�����jd�S�@Y�a��H�ݓɫ�e�юqEh���X�%�W��s�X��s�
Ĵ��r�>B�D��KSE�D7�]� #��X1ja"d����E�#�~�7�d�m�����6�,m��.c��ӛ��x��ޟ\l��=
�nBfN����:O�#�?�ezp�0����\�Z��g��7�yUv)�S'� �Pl�ݭ�X�ԐC���塹���	5/'W����ȥ�iM�0�e��}�ș�i�`�������|9�^~����#"�Q�5�{/'Y�bd�6��!�\4����땺3lH�!�Иj�j~�X_�jS���q)��4f	pJMy�m㴳��h�zI���>Q����Ku�2���J;Jd�ʿ�����_6c �d�W��с;I��&QW��`@�Lj{��`h�
�/KfM�T�_�}�F��꽎fҘ�c%�$�O˴j�:U>3���` ��Qc�?����z`����<��\TG�1˯��]���;��I�%�4�o�f��>�@!�u���R([3�+d�~[:���3ݒ=��Y��Me��rN	I��W j���F���gУ_�e��N��6GN�pI^��0�����o2 ꛢ���f��� ��q����N����ӐպS��t���{˭��m�e__d�`\%��~��(��U3�n�$�稁���&�ؼ~`A9�-qaP�i%R!����㞔�f���	O���ڒ$��wX�M�<�.1'�@FU.,f��$���:�-CET��)��<��F6�*�Oj�>�n�]?ތ|m����ٲ�� ��
���ed�5@�XNq�UG��7L).�tK����1)��*a��5��i���z~�!?�{`M5�hNe�_�4�Z��S9�$k�u$�S|)�18B&}wz:-�"*��{�ÒB����i�Ġ�YM�4�/���F����@I8�X)�8�SU�4O���. �҄����s�W9e�V����Z@�{�d���1Wߥ�}*�6�y�G�h��W��w�>�YhP�}/F��:�LyE��{D�PLp��m��:��#+�2�3�|3V��y���%�r���>�,�&V� e
��~K��6<ݤE��@�_�&�������_�(' J�H�C���]�}Z�6��Ͳ%�/�ܽu���6sb�u��d;�,/��	�g~���|�e�E�EW#�g��:�*�`�UaR�L4td���U$w�M�_ӄ��L��%Y]��|S�X�>�E�=pE��q�S|�Sm���<����3,�@<��U޼/;�OƈӌNAN�mm�w��I�'�-��2^W�(�s+�#	��3�`[���9� ธ�s��A�[x������냣Ok�94��sh������
���A>N��LQ1~MqȤ�9սi��*@Z'wV�=��- ���8�xW
g����Fqo��x���'__��B�U�����{H���W�0#�?!a�^��Z�Q�����d��F�%�g*��g�$�ިO ��&��*:;��ۉ����P���~�lǴ%'#z6щ`��2(�"����ʵ�f�+j�#�T����/H�,�b�]�e<"*D/Њ,[���<X�2�W�sR7�.~-8���_�P�Hp��N��m�T�~12i͠�x�]���#���<P���R>�{�8���&�'>�&�f����}zKR�*}�Yӥ��"W�'�X���>�J�,bw���5��+_�G��E�RMr<��1���}���r�䢖���]�H�6<�P�:��AZ�
�304|��ى�v�W�T��L����FB������s r��fQ�C�s+�c(���3�����2Ku��֌xԎU���pO�
T�o�=��H�;��Vp۞2*��'7����:�sʹ��Huϧ���Y���wW���h�WI�(�9�|N8_~V	l�H�#��.`�Z�P����9�y�H����3�-�ј�E>�YԊ�H�%�c�n�XP��Ă�<GĊ��%%��+�픔h02�!#����o��q	d73zw���/1�� k��*�e���*�U�!.�L��@uVa����(�������q��iX�
:�K0��G)����s6�g/s�uR[��zfҦcI:D�7�ƀ����p��95�8S�=|ouE���Iz��e��XprS��0�4�d!/� ����oN���F~���� �e4P��9Lq9��5�?�=P���ts��.oc0��Ъ��^}A���t.�!�ugX��2�O�5gr;!ò����eE��@�\w1�%�҈U$�4���Dϛ�v��!s�o�A�{��suP�X�=�צ��ڑ@���xh����F��Ik�*$̊�6���vQn!�#��P�Y�`G�<Ӊ
;R�cl��m������m�vF��悘�� �:jm¨b�u��`NȬ���-����o��Dz��O�B8h����"�-��_�*[�gH�y>�?�6��ЃpA2l�M���h��������b{Κ��8Vq#� a�|�v� 96�9dn±6���c�$v��u#�W&��s�Įi���>��p���wؠ��"���F�58،�|��P>  뛹s>;aa��t�:��B�&�A�z}e���W!�ɫ��w��z��Ν�$ۆ�8�f��/�K%.y=�ϛc����8oc$:�FP����.\�c`w2���^�0;b�XO�"�K�V�$@+[�G���{Ÿƥ����_�ZE����t"= �3�7�?�̖�0m(ɾA�dq�p�K�ҡ�9|�JZ~M��oxS���ja�g*�7��Y/}jA>����]o=,��b�?j!�|��5�i�S��Z3�6��P�5}k�J�wU�u�k	2�)'��sJ6i�~	ǵ�9��v)N���uFk�$l�0;����C9�ki-+�h�:g��m�hK�������'�%���H9�����8�.��������(��a�H�d��a U��B�ٶ�,����Yʤl�w�ly@��wI�բF����פt�ws:�M(�c;��5�o8ȯ��𪉂�G���"	����d��1�>��ɀ:2r�2ce�V�P��z-��Ă�٘T%6�,O�aGi-��eړ�*��j�������>1=��o��SMr�GT�:���:Ԍo眘=-]�.�)R<섏�6��{Z�F�ǸkS��k��������Q#ѓ���C��̮	����7�>�%ʶM����U�)�U�`�ɤ��*�D�����c]{(;`n�y���2�bO��� 0�m��Pt2�V�{�l�A��&I`[�$q�w���d�{��[�hׯ��@�K!Um��� �AMO�-��Y
�n"��� ~V������a VYɇ\�u���=��	�<�X'�,����K����\�E��޵�z� �'�C+��Ҹ��t3�G��Lbz	�,@�Y_	�_5��H���+��R���1V�FP)��P~���ӕ�ű�x�@���E��}2�5���0�<��9f	Y�E�#��x&��5Y�0���̫-���~5u����O�V���z����@���wY�
^��c9gz:��m�;��b�/�{d��u=���u�
��'s�'WE�ְ20�q�t]=K��cqC��w�Q�-/�\6X]��J�0�,�/ɼ�L��R�M�$����X(�,I$�<���������۸x2��5X4��>�m�Wl������J�O2������ߓ� N)��X kճ��1K���1�27ò6ؒ���E�ݎ��L8d�&��v������^.��\x�3����=��> �&8\���@��+Wԁ�'*S�<��d��Q����q�2 �tVA�È�����(m�drG�aʽ�S��.�R+�����A��oI�i#�[���A!�ҙSyG.{D6������?y�A�wr܆0�!b�Vh�(��?3&0[��i�p�f�|��/��$�V�]���5^�ܴHuKc�c����㞃��^x{�.>5�JT⃼�L(����Z�'ǠbZ��J��x ޾E��ߣ�b�r�q)ٷS��q���03%��5^������l~8u�V��֟����W��^Ƹb�>u��S���tV�Y06ў0�*p�7����@�ͱ�
���,�s����Iҷ�[��}x�Z?�e2&RWt�����)N����7.�F��2cIʹg50|�ӋW˪�	�H��ϡ,���E?�꒗6�2j�����k��?8�Z��,�y0bU9�4�s]�o��-�l'�
k��c���H�W����O �{�sN�T��Ư�K��r�~��2v�	5r�*�M��9�8g�M�
7U��Fe�����)��<�t���,Lm.�p�Lf���T������t����Ё���
v���3	-��j׎�I�g��(8���T]1��: ��X^�j:�6�tno�0�}��r9b����ه��������~ha�K/��D�-�C���Ff���]�1�,[��e��:xl_P	��o!�&�1��{j0�%�@�X��c��KH)q�Q;�} ɜ�������&Ǣ�<)_��>1n!�q�=���ܤ!Yi��0tN��&����%\���Ǩ6�5?,Z}ԙ��E�b��*���5��pD�5rri�=R�>y&o��Pɻ1�E�)�mTR5衢�O�-��E7i��ϪkYfz_����kq^�0:ב��h���o�o���r���vM���Eݣx�-��nڊa�\1����&Ys�W�f�W���_�!B�C��X|����G�I�4� 4��iolx�ϝvps�����[��]Z����r�����w��pƂSl���=0��jj��gHq�%L4�gC�{���u2?xP��l��5c��DD��B��I�3�Y(���.(Za ���)�.�R���s����ݗ@N�ѭ¾�d4�;�@�����)�дn�_�B�ŧY���/���,�ƞ�$���6�V�I���B�B�LM&��F!(�T.?�ܟ�����}-R6;�Lp�0��� �}yS��͎�W�J7��Z�  �u&��r��)���q��Ae�H9}�z�C[28�sQػ��� 4Ѱ��FXC�����/K'թ`���y% �����cC"�t�pu)�R~V�wFTIS��c;�3�l�5�&u<JBF*>Op6�d���y3������4���y	��7H�7#B��� KO�9�*�$X��]`���?�n?�켨�yl�;�I��"��o�|?�ѽ�2��{�U1'л�
^�^��N�}������~���+�<�� .sR!�D�	�ĕWZ��U�x�S�FG�tMD���KP�N9��}w�\/C�d�<�ةɧP9AǑ`���� p��Ϣ�U���a�`TW���|�ʿ_gC@�����:�\�����pA)����g�vD*ς�򢢼��AxK���|}��6e�:4NC>U	�.s��c?��S��Al��]��P-ad�A�����z>Jl��/��!����m�Y�O���]��sn�����G�0�$�v��aU��]�7y_8���p�,;�B�/R�r=�a���p7�X@����~�^ Óy	 RXi���2�<�M��Pq��*��0�#�O` 4k�a �X[2����{��-�)Os	����:���z_��T*o.��nj\zğ��>�$����ݗ�_�W���{hMI�7�.m�����]z@ϟ�o5�dA�����`j���,��}WhBj!Ǐ�ܩ�n�O
<ͦ_��K�?��X-��8_�H�L"Ĩm��W��9�s�;%��x�Yza�^XgieO���}�r����mg������DX�w��EA�M�O����Tg)��Zi�7J�t��I����x�����ӱ 2�{ن�3��'� B,|��U%�����*�I�g����>�y~�%�s^�l�����Y�m��4��B�B����	���>p����9��ŋ`�<�h���}j�N��s�a�}��34W���K�Ņ��W�U���vb��v5ɋ�������ۯ&M�����{�`��2��mo��i;��s�]�E�n%:�ֿZIf���F�� l�����L2���.E�����ו����=����a��L�/��0*�aڹ�_�d�+���g}�"����1�$�>xH^N��,�J��A�I߇Nc��9B�}Z�~�ˏ�ņ��o�z&�[�m��0����g������S�p��:�U���4P��^SY�n��g�1�I!j|8[��e����16���7Z�C)Ē������_�h��{Q�jS{$��
����ds��n��E<+�J���������Db�ä�~ǁD������8�#q�d[=��6��tH��·���7��
H������Rϲe�y����R�C�j�4�N�>и{��9���O����4����	ƴ�\��:qf�w8�t	��5�?D8e����$�ZǑ�i<HB����h�eb�:mu�v����������l�(��~��\���84��%A�u�il���q&����`mt�~V�F�uE7��d�N>`�!�)����¢�8c$K��c�BE_�Cb��z[&k���������� �uj!�&=Vеÿ!8���J��B#0�4��ʪ6L����2��~�͕]���J��#΅2L�u���������l���km�S���c�'�';���DMt��/N��{!L�CK�oD�<����̘�-���7����6�sf���v�:���ͩ-�*�nX��� ��qh$�R��X8�oɫ"h��;���s�L�Q�
o3�8�V*b�:=�	}C�+B�e�|�{��Num<hZ<����^e�9��d%(�c����-���O�ա-��|��_�!�m�#��}�HNל��$��`���@�3s,�A&�n��S6���Ǆ�O��V�h�P��v�	|��ai7�c�	�<��Rk��;���]jG-%n�%t+P�[;�~l\�h,��kO�e�χ����,����I\l�P����n��ғ�+�򦶲���m�ْ!��>�;jJΚ��3*~v�sG�B��ո˖,RH3S����W�L>�(����(�iߵӎ ӌ��ؠA�#�<,ڻArɟJ�B8��2�̝��(�_�Kf�l��
��eM����B�D��2C���)��]D�}ϻ�����a�>�̓�
�$w8��	�^Һ�#��;8Tѵ�WG�+�� u"BKz��4j&lް3�݈�ǫ��0�&��vC`ft�����������}4�����0C�,-ki8����;:�����Ǟqړ��.<��*��gx�z�8ц ���BX}��e;aW'�-Ϧ9v�#�t��1tL_�o���@
_�u~	�{��,^��3�a�*ݧM�X��I`!�,����!������`X����s��=id�&s��p��'�+����zJ@
j�ʖ��,�7��{'D�@{���5��@�}Xrv$��3�?Y_~qk��qWh��bc�t���ʟƲ��9�;��Q�!�.�چ�YjA�:��
��g�(����^���z�w@:嫪	j��~� �u��u����ٗ#̞����3W���[��z��qo��s�t �-[��y>��y�s��\��2���ߓ����(�?.(ڑ��|Sx�S��ȟ;e�^������[��c��B1;�$Z�*���{�+����R�AP�7�Id,��*X�#dr��Z[c�i
���ț٥��)�8�CH�����G�(�g=�1�,��Mj��C���E�_C1"a�ZN�f	[@��l�S�"|���3�՘�T��������@��.^�x����ׅ���@7q��� D?�f1iPd|%< �>�=Wưi5||�NA���1�U҆$�2��kO0I�aE	�<�o�5��&��o�`������r!��.�nШ�`Ԏ׃}�,w��,�M'������b�D� �(��O��z�X4�2���v�e3f�W/ږ�
��?/�C��0W?�!q �(z9�n5>'� ��c�J��$G�c��~,{��)�`���l�F�1����B!\���4��Y���+2���|�m/)�N_h�;1-0>�I����'�ɼ��&�}��5���A��E�J	�}R\�(�nd���Էޢ�8w�B�׾V��p��-!k�!��w�>@`�&f��A�%�)�3�|4$�FIđ��.Ԑ�C�ƒAMo��uD��?�)�(�y|qx:Bn����`����;�w�©t�:���JcE��rHk/=���2��^HW\�kc`�ٻ�O�2���k$,~G�\f�u�� �$�HD�#:~�"�拱g����M��\�#��c�E��3��9u�<HG�^V�_�1�m�n�����F}�{B4�2��aU�~�-��#�U\�����r�o�2#벫_��E��+ӏ3��(���`U�IRZ�r׮�hh�w"�U���D�gۙ��|)���q���k�_������=�'���J�M��X�mf����K�d��g�P)�0�v:0�yh/�bz���E��C�����fIli��:`����E�����V��.�d*(��C�)�k��a� tf��>i)<���Y�`�G�$u�-�)�HZ�u��tDp�2O���|�+s\&��o�����e��>�W4�&�hS�A���f�ِ:�r��&R  �5RA�Ri��x�5�V�:�-�p1�>�PL�V� -�L':��R�0�K2uW�]����%w���������Sh��$����	��y΀���^�Ue��)��;�M��}\�*EԨ
Q���W|}C���b�TS��7 _�j��kʷ����4˥��M�i*��Y��ET��nU�E�MGbr@C��t�^�N�,{��0;�|��G�1m��|G��f�Y�C�������4�<<9�ζ�+댡��� ����Psb��B���h��?6,�>Ǣ#cP!+�9k41���K�5��,:��F���g?��Lm�f �W\1R���%�Ѡ8�)�� xY�C����+����8��mG+�5�UI�*��l=^�0g���Si�:��41m��W�:t*��2��(>���ܭ�z.1nNIZ��`(��v�*��o�5^�,�����.ڢ�=���6Zh���x``��eB�&�zl�|�#��ąQ$���P|7�+Kv�$��7Q�-��u�U�NB��xȦ��~�1]��>�¾�Lc��L�w�g�n�ګ�$��7}�{�w�`�����|=T�Ԭo��0<��.��:9�Oi{.�6�4>·���ҳE���Z�C�O��`��Z�P1���];nb6�e3S�	f>/���0�Ms��}|w�[oi�-���d
�a���	�_ҕ��g��ڜ��I��`�F���z�dVЃƶ�~ў��$�$:��,U�QV���Fӯ�?x+-Y�j�k��_�\{�j�jw�g��
e,{F���.����0R���j�e�ADdwχ����63,��zn�*�0M�l]�٥$�d��+Yl6v2��R���]�f�1�#I|R�O��W���:�Yi�Ki��_�>]�$_�+�g�} �l;�	Gq�[���w��a���C��<�Q��^�*��8[��9ـD�tHS{�!�����{R~�0)�t:��4��θ>�
1"�0�(��"�������n�LJ1�t<rL���@�rvma�&����pl�n@龦��>*|EV�-l�&zS��7���(�J��z�>��cG}��8]=�H����qp������	���]��:Sg�y��L�T�0G)n��:���>�z�q!�!�?=L��n~%A���҄��R�B�!���8������)�Y��G�u���@�o���yk�T�����rg�����#��ӭ��������o�82�a������H�<���@���������Ry�u�����V��ܹ��9,��lb�-��U~ڴ3���O�r5�[~��XF�w�lW���y�Yo�Κ�����2�� 2�INftu�(�KJ#�D����>�n�\-�ŭ_W�Iޔ��|���F>�&ZP)�J1ᖟk�J��z�P�1�H��64����J������z�C��D��m/��Fqy.��y �d������G�y�G�&����G����ƭ(+TP�#�n�_f`"�����8�*�[�'���	L�ma(�)3J������N�l,k��aQB`hAZ���⣇)�t���pk�R�]�HĶ8�N�='�qC�˳���6񧩶!&r���1;�K�o٢e�i�1��5��Tz�w�L���0n�B��?`�����;�B�CWV�����MF����U���Tn:JK�V�P���8�-