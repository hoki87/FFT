��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#���������l��U�~�׏O����j9�PY���`T���x���s����uí������P��"��b%>�1eτy�<�gܰ�N�Y�	� {��I�ɍL�ݫ�G�R�k��Q�!E	�5E��.��:�͂2��y�m�-�.E��i�����YS�
��@�H�ۼ��nD��Y�l"BU�.TԊ�=�-�����q���Ǹ��j��ԋ����tr�a�ٵ�]�b	��%�ɔe�)rYOjX5;V��R�������M\�	D��ҏ����9c=�Vͼu��Ro�P�Jf�tRvsY��c�"n�XO��	3g���Q���^�Bʹ�7gQ+Г���$�-��t�8�����A���<����l-��*�|d0�<-�{)�I"�>N]�[!E���3��SWϣ���鲈�ƅl�a��U�q0�؛N�L���[�X6~�.�Ţd	�E����x]���]�!��5;���Ө`��F0�+@,r:Rkf���s���c�AE�����8"0�6�eQ��q��^��Z� �L%�&��~�H.��r^���}���SfS�:l�J/k7�'�\�w��p��P[�Wi�k�A���{G���C2�>
.�k�v�,g�NZ��)��[}������nf^�Sh����В�zb�2�-o�-�C�"�1F��%�x��:�,~�Z������qW�BJf����꺛�6�8��ED�}J��1���#}�g�R���7$��=$��|���OԘ��o}&kݾ�juח�ԋ�ի�"��u��p�@�25)4' �Q�TAJډM��'�=�u`�Tgiq�iI���l�q&?��1���.HF|�?�&.H��0���<p�����k�[_�ȘD�����*�Jq�ˉ5�Lk�kA-+ч�YvԋI���ura��`wޫ�+��F�Me��ǝ�Wm��"9����� p��Y8)�*9"W�e_ >�ËE7P���z �w|�#�	���߼�R��Կˢ��	Q8�����Ge5'�r!�@�v��m�;8ydD�Ï/J���
��bނOo�
 %5q�G^�T������(D����d��Ѻ�IK� 5(d�)�Ĥ�"��kT��1���)C�TlB�W�N{{f24
�k;����N4[~�����g,����,�>�E�<����=���r��ӻǅ�r��F��5�J�x�
�N�ހc;zM�3������
��u���9{�%�h�(yĚ�O��59?�j����vq� B<��ፁ(��B�����ć4� �w��A�	�-"�OC��j�2e:!�m�d~�d����8�H����4ϥl��ª�������.	�pH��bX�Ϩ��+$��)ï�>@*�k�]���5�X2�0}��"bj-�n�V��R���\P����e�5-P�J�ç�	�j�4<?�ڞ������`	��}W�HN/l��;y�d��@�8�b��K5ɳ��p����,�<��Ƚ����M�_"Á`��C��K�	?JU��أ��s����ݾ��m�\'A`�؇��ʼZ٣m����Cm:���p��Hp���o�,�`�M�-͇��Ɍ�}б8w��Y�&��?4�G/>'Z�cX�]-ѿ��o��<��Ю$9�Bhܬ�z���Fxz��FK4!ָ�VH�
s3K]/���T�u�C�9X?���1;'�!K������;a> W|���nŰ��F�f�d��M�t�^��ѽg`x�<��ŠıT9�#�u�v=~�y�?�؞U	ΟW�۠ћ~�`�Y�m��"�B�8G~	V$�&���oO��0���n��5�������Ue9>�Cؠ�5�g@�f��T�����O���M�o/�8�tQW����Sb!K�@9�P�ſy��nd�t�DY����gq��65�}�sSp���g��x����F�Ə�%:-�(K��|+e�-
O�\4�2�:b=�.E9|˯�?�W�o*��-GsT�ɾ�+��ڈe���&��=e���5VP�mQ��~7��o�5�d���	��MG\��Rr�"I��!|�8�M��N��� ���s��vr6��y�v�"��+om�h�@�˂�9�z�j���c��~�JT+���F��@;��Rښ��kSSfe�s�6�������cf�!I�-ݭ$֬�Ҡ�/B�Ŧ��W���4r7�:����/�w�ӑ�nft�9���9CB=��m�t��G[M|���2�h��o$�	2�&��Ǽ�Sۤۊ�&|��n�`����r�Z\2ɥ��t?�"��Zw����D������E\���Qz�_,����W#Q'w~�|�ߤO:!E�v(����5������M�r~�MI��xnE��kK=�,�'�����̒�RIa�i����aLS��Q��J�x's��h|F�ƆDGZ����p�$�vA�0G�|�V�M@x~��q[Q��Z���J<�o*�[��.cG�b@âI�N�ħ�?��=1KZa;QD�怣P]�p�#���U��L�l�f���5�k_ŕ��_�1TO���qX��� �*P<�q���"�������缦��G�B�w� �p30OH�6G��n�H�' <?w��@�(h�c���ڀ��\K���)�a�$�ȠJC	z�<�ö�_L�,�l+�����B
�\��ˮ�o�J��쵚s����ka��E�7;u���1z�H��ɶf�	�je���b��%4Rf�}LE�6v�'У8��C!���Ν��*Eg���)/'_ߤjH>(F)j?1 N@�U0,�9\'�ٶ��f y��c)Vt��}0�F�DO�?f~�-;���U'm��Z�J4�" ���%5x�#�J���1��M�V!ӁW[�(�`�y�H�/>	�E���L�Df�KS�%�� �ZƂ�kmѧ�	�]��o��1S����<������n�3i�����gMʹ�e��Aܕ_�H6<$�o��&�Ȏ���:ݤ�{L��FЎJc��uӤ�RʸJ��F���l�m/�`BZZbWj�|�N�Qb+�H�����7"e��؏+)I�r)XF0-�������K�J^�Zl��^wGo���+�ÀuP�N�-���w���#n؀����b!��|���vԭ�߼�4�BM��N���n�ܿ�{zv���{�Cd�1&���Y�S+}S���HB�}�n��.L������怑�~�a��~3A��B�i#�����q:y�og��f��.�����=�p2>�$�y�Rr6i�2n�,��z@�j�c����ʩ^�%`�;��Xb�&ޑ����ar/���GKT&X��XSMLa�������
zq`>:�6��S$���AtH�u������ur55b�)N2<���KPjj�b�9 �R#0��X�)p��I�3�s��Y\��q]Q,��o-�'�>\���=��qW���i~��J9,*�95^�]��QР,����=&nu����{||��s��VR8����d�6_ޙ��^����Ub�O�O�>��)B0�#d�E��=<��XɄ���}T0�
¯��c�%�V6'��'B���m�A�"�Wj@h��}X��
�̂g�n��v�P*�%0摼6�u0Ҡ`��)�_![�2�\�M:Pm���
����)�&y�Q06.�=-�`�������������P4�~4�D�:g���.�.���t}�id��n0dq�GՂ��x�Mw�#��짖g���>�<������Sg�5,�c	�l��\A@��A��$%�ZΗN����sSz�2x�Z
�<�	�._����
��)'�uh�Ѯ�ϣ�Ao}X��G�HD� ��y�n�ڐ�cKbz��b M	�//�ۈ��=EJ�u����'T�*�ң.Da<I����6Ec�Z��j�O^6-�����e��a�YC	�O8�Wz"+cʛ'"�C`���� �}��8���΋�n o��,�8�)]~@��p}���<Ҡg24z��>z,���أ��soƩ�]3+�6E�����mG�\��죜v����yZ������H-	9��GdgDa�z.m�e�0��^0;<�|�2��їmX҆�f�3O9�f�����ڢ����D����~''Y��@ڔ!Iź;&�3���~���T���N;y���M��8~�?�U��v���5�dҭ�Zl�W#����O�z8 �z)�>��c��ɍ��a7H�/���GKA�r܄���B9���2#	P=I�rs��ܟ+�y9B��׊�~ �A1%�����O�	D�r���H���[M��vy-v�81�R�� d�g���+���+�:���1�P��G��3����U��"H�>�n��W�����b(q�AH&���$O�}��9̥�̤3Y3k�.y��\�mvH�XuE@��I��3t4�=@���I��H���b�:W���Enp��q�R8�}�.��b/�,�p�����8�{{���2R�0���M���_���kT�Ԋ�=E�ѯ{�I����x��OBǚ�t�x��O|��G�sҨgs����x�`��ϛ���IS�x�h$s�V�#'.o&TUN[Ya1�-���Lϟ_X3������Q�j���I�t_9|��U0`D�����v�V�z�����Bv�b����0��Jej�@������ z�j��КO���xM��c��j�]�G�X�#P��YX�c=��#k��@	���)-��j(�
��gn�T�/W(1L��rZ]�(��r��S������Q�5(0n�sl���xT)�E�8��C�a��D��le{���u�AMI�o$��)�����M�����ϱ�iS���ܯӭ޹��>Ҟ�GW4T�$��t;���4���Sj����fs{�Z���"��2���O��K�n�UY�� �}�:"/Ȑ���6�vJ�7P�c�����vp��0��u3[�q�K.S�g���ɂ2�o�;�ۍ|��N�B���L��r{�6����2-;6�ò���VӖX���yr'����|�L�6��ª}�2v�ɬ����mv���P]x	.	�Ƌ��Ȅ�I��b��c�h��z�g��%[�$��B��2�O:� e���1$��CLjo�m%6���+iu����'�<���|7rU1v��̦�U2/X�3�����������.�;�_�5߭߹�K�j|��˾�נzFhs�5�fɜd������eyP����4��]FH{59Ʉ02�e�B��I�Mm+��.F�uo#,1H19іߊz�DK���%�{.u��er?B<C�Ǿq|�,������&�{�К�ѣ���l��`���b���d����I�/�V�t��[K
�FR�.{���H����E�5�q��MJ����U|�>��L�;R�������I"�R*h�P�+���F�����|6$#�؟��oN�Ju]�8A$a?}��^�xKn��K��e�_��QQ�.� �~.5�M�Ep��^����%f>����DL龽+Zx�b}��?��0�_D�(�j�9����E�!��%2�-"���'���dm�s��|�)( S?���J}�7�w��9|SH�6�i(�������"[�;aʳxbc1���Be���ի[#w��i�d�+0!�l=[;5%��� ȥ�SJ:Q���bs�w��AS(^kj����*&2x*RqB#��.PL�B8M���;��=��(�
��w��IS�%����IE'Q�m3z�'�fS���t/��T���v������èo�J�d{���f�k����iĪ�r�%n)k6xU?���ዖ;��
8���5V�w��e�0w��)vM��'X4���8;{�y�j��+rkĵ�-`����N�9���|�a���(ݱ4�T��SIn!P�adr9�'��Z�I3&?_��^$�v8�:�T��`���g�� �)\��	��;p/�bsv�+���K���r�4�G��)��'2��5�W���7T�U,)��:��51ʼ�q�ؽ�t)�ۨ�@�P��ׁ�.p�v=oc�8�4�i��fˀ����N'�et�͔SQ�O�&�}��N4.�~��d�/rOg�f�_@=/�Q~3��	7d���:�j�ZO���M�1����i����k!`�픬$l|��[���(�O���A�yI�f����^�k���.����d���).3��M��.�3�4h�#(&Q��@�9��+A�i�z��7�M/1H�?��(�j@jp��G�p�3��i}�/��M 
=E���$)	�d72����)��b�y�)�{���a�*�Ǩ�''j:���'���6��]�/ ;�7�4�2L[`3:ӄ��o����"qm>�k���żݏ�Z�r���~�U�������({l���Dq��}�Lc�"0 �U1oᓵ��u}z�=5���t��p���������\oB.P72)���3�HBkj�Ī�e�rc}]cL�R1�RQ�N����R1[Ύ<��7�Vd^�I+#���b;�E�f�Arf$��S&�"��� �1�|�%-H���p���ۻ*���C�&��wS�%S��;<���p�H�-ڤr�d��� �?��7�3���3g`0��()�v�.�Ԇ�ù[���95���^A��$��ݢ���>��#�@�l��]���ga(rR2� ��0=�΋�>�؃�읣M'�R�J��4k�楈�bKZ^H��9*di��71��J�?&*�<�+�.w��«`1���� -�&<9�iĤژ�����s9qK_٢Lk&�����E^��5Vײt,�1^1k8OV���	�,��ӆ4/�:	k��J�t}<Aє%�nc����X�y"�e� 0�D�J�Z�䀻�7�`�����qo��cF�D��q�eσt[8��Jf�v��|V��\�p�?ޅaCf�WP��_<�)t��f�,9���4T�i��S-��[�$�,��m[c��R�����^Б�_
C�yo%}ը�"[|އ+����Z.P�T���d��~C�p��b?��L�1�Vu!'=�Ek=���F�y��i{F��&CQ��uQC�c�L��� �������DB�[�fQ{%���Yl���)a<�PK�C��<�x�e���JX�q5�h`�7GiP� w��J�,����E\���PG�ߏ
l�y���f��.�e����O��}{�/�p@Uh/�/iY�"0Lw*�<?���!kD�,?�k�ӽ?��� ���`�`��/�t��Z�����c�lqw�(i=K�ӉнD[�<�k�� ��qwl�&5�4Ʀ��?I{����Z���[�[�
���N�6��W��n�l-�� ��#�$�܏J���o���Amog>��.�i=�����%��d0K��%�q��
:�Bق��	��;���Q����<a���S��E�wN=�E)7��K�QC���昨�I�r�X��mϚ5���w'�B�&Oݓ�i��0���6='�������RVf9�p=��͎�K;�i��{�� r�i�C������|X��o�"��I�46�'������Eh���ps��?�iy�U^)Y�va�|���C�23Gb���hf�G�B>�T֓���ߝ˃‐|M2��c#,;m��2}}7�2�e���K%�'��?aF���d!�n<Z��n��x�˼\|W��ն�軬��uF�Q����D�3���@Y����(_#�4���ֈ�(�E�:����	b�q�==e_{���88����cP?�i7�'Qlg8�z-<��2CUɏ� E�s���}WLMg�Sݟf�! �P����.����v3ִS�	ҽiq�s����4��[�^2c�9T�`�L�V΅�A�k*aN=8�M�t�I��^���	̪�T��y[]�ur���9Df�x��2��'`��Hu��YdtC]��>��f�/���,�$���״��r���Bѯ.���`ࢱ�q��8:�j�	��L4D�B�)���r���t����/�3(O�G��=Vp,�q1���psR��[���!�ֳ��M�4\���j�E(2����ZRt����&�C�t��Af��䔂���6X�39�9�
+nuY��y��	^1��<��Q��\L���EwG���@ɠE�<�r�J��/w!���@�~�����pf�n8�z,��N�E�����c��+�	`�RE���.��w���7��5^z��5}3K9GfнӵRed��x�}\��T�7�,���cs�[��IZ�].Z����ۻY�1��'mr��K&{e��F�e�K_˼�K�!�66D#�h?��}��*��z=B8��U>�=|���A�hB:od�lѷ$f)/�s
WS~���#�{T����Y<�� LC���A_�)�UjW��jCPsC@�:a�Ӷsqa�eb�<t�-��$y��ņƻ�����#�J�2��Z/�p��~F�u�)�VÊ~����몄���'����K��)�QB�+��9λ��M��k�V3�n�V2���'�
}ĉ֏J���o�$��3k|�@rg"�`���y0B�������L�
�6=7~7A��&^����b,`7�<]ϥ���ے0(�Ch_�&=.��i��S���C(���-,�c5Kzc�}$�9Kf:�3z��Z7���K*�)� ����`������_�ݦ2hhe�Ty1
ηO0�R�1�9�d��n�>m{�f��t� Xs�>�c�2M�YqM��!����&����i�0�6m�T�TE����1��W�36�x,�T��s-ss��PM<�ʒLUV�>Dx�y]H�xrBC��ձ�S�Â�p;���h���EBw�����޻{�i���=��۩���/5
���Vq:z�/��/Эk���T6H�l<�t{������]=��Yr���&�r9!��Ϲ; $�\�\{e����y�}���ξ��wh"5t��ד��
�3�˧������#j�Hi=��FuhG/1���%��>:Y��9��⫅v��yH��O�6�����MQ��֌��j�S���R5WẏX���8���|��7�zοd8'��kl�6�lOVf�"�H�h,�b_\ԯk������=�����eX:�V/���
�?ڜ�87	D#�0�7�/�e2p�\�a�[om�j<���CI�	�ouʩ�/ 8�K�N�}U����;pY�D��j1\��gP�Ci�v{��gH�U�ɯ�(��]z�ĻҊ�'�3�L���Ǖ$?2�3�{�U�n��3�U2�p2mZ�����z؇�M��gpc�eE����i�t�5�0������!�
 �)�Bf�-3@Wyp�<tO�iF/I8��*
w�A1��n���X G��x�Y�lS�q\Y9^�h"^]&�Kb�Ѕ�w���1��Q#��в@�<�?�'Z�H^w[j�ue�c���ӎG�$D�,���C�[�Ր$�k��(2�������0@���RI1��Una�Ԁ�#��y�1���愸,r�J�SV�A��YPhVF94�T�n���T�f{�k'���A�~vN9*��w�|#H��K�I��x~���F�|#�MG��L�>�9o�"��9.�m�	�p���O?����`X������l��	 �(D�bM>���p�|9�0���6@ºD��w��Rd��yd�a��]8�QM�ج>Ȏ�L��2��9��em�����Ԕ"��j�$��|��}���p�o�5��ď�L>��v���,��c
��:��(;��4��q�_�O��a�Է�v���ާ�m��8��FV�I|Գ�����-�س)՚��~���rW,P#D����+:'Sd���eI��x�!S,ʕ�S9�}<[%��e��^h�,}ĉ��[�
k:rUD�\����~��
��G�ʳ~�����b5��J�W-��~��. ����K۴V-r
HNh��G��TU�^�;�jV�����,���z�U;#�� �[����d1���l y�Y��'��� �s.�����X��\ю����.��\/�P��3Ҏ	ؿl��|�n�42���qҹl�D����-M���`�u�GH�̄54tn.Yz�5:W�b��*��(8�5ϴ��@�N��X������?r�+9�*���ȼj��Ʃig������a�zh����v퉀,O[�8� �
s���Xm��jh����σ��r���))}#,j��DL/��e��m���O�U�B"Φj��&�<��VzV��f1�?C':���g�;?ɩ@�S@�oӬ�׬�DWM���Hd�������+D-R'�zv���1��&�3��hU\*˘�v\jg�P��1P/Y���(�I��޳�Tb�opz]0]&��M�9U����y�/Jس^�<J�<���J<�q�I�I)�7=����T�H��$I�*�
F�,���u�Wx޽�0�\�9�@>,�Qg0���X�&?���T��)�|���Y��!����
]rb�X%���%O.�wd��ء/(��&�T���gR�+@Z2�B�)�6;�[������I�f�wTQW������& r�2g��u֖o�ԸyS�v
uN=%��=%c��{a����z[O?�\���_KJ�iZ�9\#6��t��6��0�f{#z�6iL��So"�WZ���:�EG2Qd���f5c����(�g�[�+��K�o斒,~�ކ����Ek�=Ec�)���?Gd8˅����'飮�|.��x��d�mw��M;g��D��h�Q.����w��s内]KB3�~�\E��!�H&��2tOG�U�C��TO�tq��;=�{���x�m�)0�?�*�'h$;q�U�Dy4�������tc���+��M|E����f�N���)R"w�d����^��1�42�_�ٹJ��;��<��i;�B��7����+Ii�Yo��f'l�v@�2�uDx���_�E�&���)G .T���-3/70�����%Y �8�̕�6a��{��R/ï,@drN	L�	d�0����
�/@����fw�ڗ�:��X��ȼ���� b�h�e���|���.U�r��ԋc�t^���U$*�xk�B��{!����8T�ע����C��5���D��\ �wYIڎ��|֓r��[E~e��&%]�%D��������?}a%�/��ȏ��σZ�9��M�B�_����d,k1ʟܳ�����j���q��"1�e�p��!��:�V��^OT��:���! XjO���qM�d
��f�YiA�'b[�g��&����4��f���:��/1'��m����"�vh��$�5ol�t~�VjB��;��-{]�a}�m�L���A�x��E��Y�9o����a'^{;v�Y���nh��)���2^����>H��$t�bN��F��;릗z*��7!ս�n_ꎟ���ဃ9\V c�^?��S���n���L0^&oS�v�$wt<�"QGG�t�5�<s�<U�[Նn^Оf`T@<�{�I�7�>��p�F�/�]�.3�/�.��wC4����	h�I�hl��<�ݻ��Wl\�Н !O�6rA���5x�oy��o��D�u��cdx޶��3�*|=��$4�D�Z�c
�R���I�x���:"+%b��5�<�:}c�{�
���gv��D9>޶z��P���C9*v�ט��J��t�j?`t�������u����뻔�l�/��?*B��rl7���7���F�ޖP/BST/gN�`(v%'yN%q�,Gĩ߱4���Ȉ�]]�@��	� R���F����NF�0�`��=$�h�9�U�0��d$N5-d�R��Yq�9���lx���U��hƉ�ՙqj�M���!���9* ��-6�&������f ��&O��~��.ہnM^�G�{�����>z~��
l,�����j��G���)��_$�s�A�����$�f{7�S,ɸ%�7�}�N�q�MeY�A�� ��ڧ��Ƒ��͟�;�]V�J{�_y|	jH�׹���� e�$O8i^�� n]���� ���?�C?Q��,�y[>b[]�P0C>�e��>�M��ڧ|v�d�'p�z/X%��Jҫ�kD@�$�|v��VЇ���!d$j��*�8
�6��d5���/�if��4c�省�O6��->n��T�"j���<d܀�Y�f���L�-[��%l��+Nrπ��Eϯhc,�w{��	���	�����1D0Rb�ls��*1#M4P5A�Q��DB_K�Ę�Q#�w*ݴ(`�$p)��t�؜��j���	�0W���" ^��X�>����W.�w98�:B���'~@ȰL�?;O�L�ߔ�1�Nvۿ!�����S��p�+a���~���Jْ�m\��sߛƋ]z�$�x�#�?�,��U�vt�~�e�p�������Df)95q\�|�����Ӝ�kK���R��e���3�Q�tK�;�ʕ)xB]�V��;01g�t��^n���q7��N�� �U�F#TG�;�b6:a�&X��1j"K�N�q�3,���JIV��r��ƞ.&��WLX��g�mԬ��8<��qv.17zh:uu�g�]����\$�yC�6E�%���GR%��|V����TF��l@u���I��m+�C�q��-���0��-�6f)uy�`]]䀗H��}�U-�J�|�`Joڥ��O�;�)7n�6pm�V�H�G"���i��N�g��r
��BB���`�,��+�r�l�ht�DE�OͺT��9 k����=���`o�a�9W�O+������PR�>w��Z[�1f'ןm8*�Ǘ��O+��3�)^���"�c['�V6&1ԩ�B%U"��H-�����,��M>RͰb��p�ހ�� �9+���eG���v.J8h�3llM�V�NW^l�%8���ҥ�<�S������^�<�}���hZ\2�r�E��U�(�$y�ά,��E	iez��PS2�"g༭ Z�Tv%P�C��Z��-�kⰏ1�_�y�`�P�B���m�a�}J��E�Cqԟ6=:��^|��Q��TW��t.SÓ��M�ʸ��r��rP�3ң��'�2��0]�4r*��D�9�#	�9�b�:��s��sq[���ɀ�ee���/lfn�A�����1V�:�P�P^jU0]�'i�X����[�!!�t�d7��V](�ת(�R!7�D}��qE��1��q�]�p>��-��M��#ʏtn��ngZ��a]���2׍�j�Y��� �� tbi;.`����xI;�����t^5������7cKnK&����j����~O��ZsFR7��F�1��SƝ��F�[�b���9�	/�2�:�zRBU������X����$������K,�*_e1�?H�l�3���0�!'!�sv3��hh:MjXl��X��b�ؚ�0�V{�B3�����D7�r�*��IQ
X=p'�n?hс���� ��÷+�]b.z�|z�}8�T���{�@���ھ&T�A��%�PT 
��xw;�+������H=���k���)m���ާ������pZ���&�]�R�,}� �nF�MM��1��{��9[���~���f��֧�ݼC�?ic���b�Ɏv=��Y�
vbN��r3���d�յ�I�h��@cy!RJ�����crm�oEuP�ް́IPu"4�&����=���wƠv
��xM6-�s��{
5ӴM)5Gx8����1�7�'*��7����T�� ���(8$@5!�-�)�*�a�?�餫�8Ad����3pݵ������ʍ=#��t��E!�@/ʼN���7���5Cp]�g���5\f��8��In�Wo�C�9Gl
�9��ػٯ�'嵰�WǾy>��Ϻ����"$vqCջX�#��u�Wۄ�:��A��Df�a2��1%���tء̷�)Nb2��%4��VƧ�S����ؔ,@�_���x�^"&~�;Y�z(��`���+�h�3�IJm�8���~��P�����˴0���Ì�?$,���W>�W/T���۵�2/̈o屒- ��շ�����
{��i?����%�r�'�Těz�$��h��էH�j�'�4����/��)ԫ�!(FV�
i��#�8C'��/���g`��z��\g�`�gh�����K��ߌ�o���������C�Ȥ ��Oc�B5b#5W�B|`wP耱����,��?"�>|�Q=To�'��X�煪��/�`�������r���n�r���`'�Ǹ`o���[É�p�[���3�0��&$C���?��
⭵��m�xE��5,e�yРZP)��Ω�#o��I���<���Ň�B�^�PR��W�Q��B��XT���7����%�����n�����'_ܲ�%�j�9���5sP���U�ˋ���
��kx_���t�(y��I;*A�R�Z�7In/�БsL�Lfb��φ�_�nOh�X����\X�����0S>�K����~����3u�}}j(�r���K&��@�s��NS"���P1|C9�t���8ov_L�ξ���<�z75S�W)?E��_�or�h�7�������N�U�
T�3L
9�<� X
`���zO]_gίb5�?���A��Z��O���>�<g���si4/���V4-1Gd���d\����:�0�Χ�|��J�%�N����?��Y����bZ�����ђ��ī����z12��q��3�¦�os����S��w̼����:�hY.����5�%��	�X�t$�F�{��ynj�c�H�3���'����&�@��Q�%�[1r!߉���8�h�ا��&��
)���|�j꜃W��t�����_c�!��[��HP8�@��m�O����V-�[S�87���n������0:�ݭ�g�T]��MU �SI6 ���;=��*� ##��Q���-��4�e�H.2CیL�-��䞥t�>��!�&���@E�gB�#��9�����2�����e;��@ƕl�`r�CT����C��!M�Qh��A�h;m�����G0�z��vZ��R�L;��_)�b���7�$fi7�j:�vRs�G��pwX���{VRS�X��+��s�8(�Wz���ь��j��ALن/<��X�±\Fo� ��;W��� &�8���L.>��`m���
�gU;!n��}����:��}�lF}�êYt�
)��E�KNq!Kw��߿!�0�|^�}��W�֐�@;B�dJ�+����u�*I�q�&��h˩z���>p�=Jz����9����[��&`+�����^�H�[Z�Q�%J��/%�랴Q�X���"���Q�&C�J�¿C�$�g�3��]/�w���{���;a�PB�t�+���?�r��h�R6�%
J����o�*�s��MVau�VI'(��Ӎ/,[)�4wkl�b���T.�ɶ��L�yt?5�SRg�A	q	�߄%Q�NHo� .��Vc���3��CT�����_U3��"NQ~�oU�c���������מ�%(��&��U3��q؆�����>�SWm+�V���8m�j �Q#3���PД^K�0��Y5Q˞5Vʻ�㋎���e�mN��|���N�<O�1��*�����<
?�	APq��q6��bT�V'���1��K��YB�_9Ɖ��<���e���/V����k^�H��b�+f���(J�Z6���a����N���Ƀ��@���3G��/�T#ͯ �@���+s�XK��M_�P�R|M���[cdTjxY�Uܐd�����i��ƅ9��}�#��C1�����$�7���bn2�М�]#<b��m�;MQXk�I�9�7y~�憶n�'9/���Bm�A���@��!ćB 3dX�3�e��e�vY��-��tik���3ђ�0����77�K^+}��V�E3��B���%�uz�}LF�����mҁĆFFёP�C��򔅄4��O�p�+� �,�Z�,��v#ah\	@��ESt�����)��.�^�Gz�	��H���2��8�I`�L�����"!�Û{���x9'��i��S��4�u���)sm���7�'����l��{�3vZ����_<��L��?h�%���� �"'����:�)���7l31��Lu�U�=�00�w��O^��(��R� f| ��NNa���C���E	ѡu�/f�ؗ�j�V�߁:͒��r�BX!.Y����1Ta���3�?�j�b�t�Qс�|��a�)���R���D͕.�q��g�7� �|xj�nϚ����}q��s��d�5�m�lhT�`���
X��<4wS\+%&0��[��}:"b4P�M���?A+��9��R�1���QϵX�v3=���1�o*�sa�t]?��z�@��^^���"�+�rP�1�ʈ�]��QO�S���	�Q2yF2?���|�K���/#.3|YP�>�<�R('五�ᩰw���ҝ�(�Bh��r����b�$6���D���oB��ZW�4���%�i�U��$?���[�f�Y��{F\H:�6�.(��r/��=7�g4����F�%!'+�G�-y��'[�����@#M"ϓN!��.:����Z�L�t�Iu@anr~[J�����YO�ݽ�hO�C�O::ԩ�b)�Rۻ5�;�ox���Y�� X���R��y�#U]�$��X>�T1�r�	�����-�%|�X��@�̩�����a��(p�@�vф���f-�-5�6��t7���S[O�==b�����5��k�Ξ/}N��X>Ԣ�+�WX�l�fp=�_hʤ��7�-����0��\O> Dj	�CK ���}�mE��kI2t���r�/��C���4���� �@�+fӝy�y�2[$U~8���b�p�:C[��$=��c] n0��k�
)P�;����'J.
�F+GP�$(3߰�.�o���	�rԎK��(����q�2ơ�hꅾ��{3���]��65��_{Q�-�k�u�yb�����l?\�J�R|5��{�B�����ۭ�ɼp��n���$dXP����,8���tJ�W�E����	�$� J7z �!:�}���;�=z�q<�R�
=&���U�>u]��9�WX&O ���0�ʆ�t��R����� �K
M��Wa�χu�O��g#� �kh��Xy�8���Yy�,5��q2@��%����:�u�H�HՅ�"���a�\��{mp�
�T&@H:d��/����SA�4��AF:���e���;�l�'�ڌ��w_���ұ`o�Ul�q�������ݲa!^�gP���rmlh���t�Y���dc�\�Fof� ����:נR���%8����]�2�\D�����d~�+�~�A���}�:Bk&qS��0넫���Nsy���r�Q��T`�/8�1S�3iZ1 �^{HT�v/��������5ރS��h��t����[N#Zd�$y���[��4��c ���\&�˽$"P��ɹ���8�
Eժ��4�u�D��D��c-5��D��p.x��On�!W�����)�4�H�/�<�T�%U�S=��;�¼�ߪ��[T������������^�-ez�-W�b
K��4�Qiha�u��"x�(��p
,�dy3�y��}�\�������X[+ފy�s���g������yV;Qp5�ҡu�p���d!q��	5�ʃ�A^N&�xS��zr��5Bp�Թ�0��,X���UK��4�1+,se4�\
J���*+՚Kd���!�v�6��9C�R)m��[A��Dxo���/�=ҭ�Q����-��r�6�L�W�~*sn��厰�+M}-����	<C�Xy��)m�Ar�j����}�n!�*�>)m�N^��
���ek��I<upmyZ�S��c�:ui�Tx�sGi�K�8���z��B徠�Rǵ�/Lo�T�i&�˥�W��o����e�ݬv> ���df���OuU2Ah��DkX[b�qg^�]LeA�up����گ��v��ɸ�w�R���7\BX;C�K�4��}eK_�����=p�s�?� �Q��2�lO�F�	}dL�:��$ V�9�Ƨى�8�z'�|��8�V�X�� �䝙 �b��	Ɵ�o{;a�BHq9P�"�}��1�"��V��4�o�fn1:������,�?�?h6d@&&�,�2C7_�M��N�0��/��K)zJ�L�	����&w\�(.���\�"��f��:�Y���_�ƭ�W���q��Vs�c����uę{�tJC�$OO��S�����N}?5�k{��9o6Gl�����g����T��:�,��#$������O�v:a[b����,�I��2���6ݍ�Tй�$�A�<����8�I%ڛ�e+� )~��� 3��]���T�P�({��<V9�м�Z�ј2q+�a���|s�KA]���qi�vZ�{�c���-1��>^��ݎK��K<cJ!U8o*?�G����B�nlJ��I��6r�rZ��"�U�N�äD�!��C����	���:nB��Ed&>�}1Aެ�i���Y*����B��pه<Z�?�Hu�
㑥�$봞(���k
ofr/��Q��b���0�ȳ	6mDU5H��C��S6����������n,4w�Y��q�P�
��f-�ީ�w�Q?��N^Q0��E�j9�p�H�@Dis��q����IIo��b_$��A=9X�B��nR�Z��>kR��y1��s�#�̔E��x���� #xt��9"��.s�[�[���
�:�P&�D����#{MI�=4B��&0�I�C'i*/
yZ���v~����C^N�@�^���I�?���C�/��B������k/w�:&Ơ���{�?sX)�����.�_*&ᤎQ�u¨��k����$T��Iun;�cS翴r�o����Ia�y���ڞ��#����h��Q����`�E�L�#$߂\�������I>
��Ğ�A�as=N.��A��'E�kIa8G��[�K��$O�KՔ,��^pgw�@!R�}�&A���WC�a�u=۩�V�t�F��:[���U5�{Aա�c|�_ )�F��=��*9i<����7ZO�*pP����eD��?����!}|kOjÞ!�D�{qa1�f�Á�9���K���u6e������v��:ב�7��b=ǁ���E�A,A!����6����}����x����Y&u���^�66Z48�V6�j@@H�^�A�OS�������̏4L��Q�2�`켨ҥ&n���G׍<D�/�=�!�����Jd���y��(ZE������n��BA_2�@���? n2R:Hڧy���-�+`b��	��Irt'��o�E�:��o�9�;ḕ�8� `�J#�	�F��V�y��:���⟈�8s$�ػ}e4�;���(^ &z�y�0*�	��w�����Ҽ�t�\&G��6O@��<惶��q(��F�pI�	uk?#,��ʙ�I������0\ؚ�'�Φܠ�j�Z���\2w��&��/�?9�����Hi#���O{�1����H*L����9rY����'$�\�]�L%�V���)z��RX^o��cTn��+%k;s��ktB��&?`��	X��UUIV3�M0��,�r���x�5#d�5V�����S�BN��g�W�� Lߤ�~��b���&��y3l]�0I���i�Ofc��ᚌ�y�5j"����n���){�ñ�]� �ę[�7��\���5�A�OX4M��H�l��G�05��wn��hHw$�����
e�:ܭ|Jc��@�<dE�.e-Do.��Aл�{+��JZ�b8&�ɥF1�m5�p
BN�EL����t��H��`��2/�d��	�$a�����(̫�l�kC����ag/8�ӟ�m��-Z�L:�:�L���05BQ�<�(j��[]>*}�j�C����j��� ڒ;��v� NJ~��/7y%�'�+�U��E /�,�]���E��s��#s�Y����~����(��<a�]��I|Hi�=���dt1�O8 ��/o"
ˇ;�����L��P���A �<�±�nw�Ø���>q/�X���Nc��o+5�X�X<\_i��q �e�I�}��صN�W2X2�%W�v�Jx^dk��}M�~��IrO>�/&�$k�*^?�����M3�֡-�TF��<>�C3����#f[��ut{�X�(���r  m���gM�G���I|��Y�6\��G%�7���xN�ϴ�/v��1`>�NR����bd�W�ش{n���U}Q�Z-[I����!]� 4�o>;_C7���Q_<�p�iR럣F�����!�l��_��;$�[�������ӛ��	�)3=�c;ұM��s{�6�U`U�5��t���bb���T�r�2j��K�
YK��EX[���ьP/���\D?^��0����1���V�iw���E�d�7�ޑo2/���Om�?Dݭ2�7A/ؿ�0x;DzR��mj�3�����q�����TCJ'=�C
�@8)z������%�\��_�Y��TǶ�V��Q�8q�iOߢ��p�+�5e���3���4�(�5�������H3h"����[�t� �h�f.�䗭5{�%[`Y�}Q�����{G�M�v ��l����a�>ˉ#���E�w�ha��v��:�ښ��C�Qk�o7SvY
�U�Hf�r�(�:��J2��8d3�0iLp#�@G�yD��􉯗�˚�1�W��ǻ:�_���G���
%�&�9@F���,)���|��8~�7Nm�:z���q5�5~����B�fv0�:s�t~����H�&@a�ў�څSw�z��)I�ۢ�ل����,���s��P@�{�#��6�2� ��P�ƫ�w����`��ޜ���d )������/g�OJj��R�/�w���y�2���Z��畔��}��Lh �[������Kj@�m(��I��XZ��>��C���/%����6��&�8����k'���+���A�����8�T����15����^�.�����M�H�,���k�T�p#�˴�W�[;{�����~�2R���o"�w��_���5��MQ�7!�g����{I��h�s�� _���bYU� ��DV��ab,��"
�u��Yf����@0�m0�&�U���=(�U%�2ŔH��m+jQ��=���%/ݻ�G�:�C��Z��"*�A��Ŋ��H�$ç�VJ�s<_(u�����F��s"ٿ�J��c������ˉ�E�o�L��}3qX�Q8�)BM |����W���h:.���H��ΗH�?{���2�%�-/��Ԅ%�P�mb����v�S7|�S+��WT�v���3�wM�%r�"���p��ش%'�emkh���hzu��X(���\�7 ��s���kc�l�G��Es	�DNV�(tE���j�ʅ��I
�<�/O�����#p%5�7e�O��)�V=�4-�ō��N䲄�]�?�a2L�Mz��ϙ�ԩ�h��ʝ�`$k����NM�;�;CzN��'��ͧ�S��i��M��#Z"%��K��`��g��	��]�4���ﲣ���Vq�zF��Uq-���z�1䚓�D� ��:���܋��=0A�!���$/
Z�?���<�y�z�5_=ѕIu�ٹ�ߵ �G9dن����7YK�\�������r6� eeФ�ÜA��u˦f�k�� yg3���,	>�uX�ˁ4�����;x�ǘ*u��{o&h�¢O5}����ػ��q�bO����]�-j��'��J:�$��ۃ�h�ɯ�p�nl�Z��b�s�n��k�y>]�d��"nH�Ze}u�:a+xy�f��J7���������25��s�>�S9�
\/ƒe�������W���J�4 k�#����jᗃ�&hy�v8�T�LL���p���~�,?��]���mAF"VWV�Ҍo�օi��A��U�|N��)P>�!��V(����Eo�p����k
��Z�s���.#��9�,�vK;����1�feT=I�Kg�6��Nn
�L˘{^S���;�(���,�i�݈X]{cA�<��|LP\��1Y⤁q��Wݤh�w_�&����Sb�mlF=�ۥh�p8#���D��ݚ���֔u=����7������#>P�ѯQ��<��|�@�Sͷ��v�}�Ӄ2�}�8��烗�6C�zWs
�<h�;?z��dsW�X;�BM��ep�/h�~����m;��|'I�����|�|�\&�÷ڨ0�S��O�K��$T"O(��a!�Y7uMrUU'��)0�c���F�f=��q���\b����Ƃ^�҅x-�?K����^�8�zvUk�9p��x>�$��P�N�cL��aT�&��u�c��{�����Qf��(	$B�`)�����lO󩁢��l��'����xq��k�
m��I������1k�,d�ċ����M��?�l�;�4?�I��ؽx�i8��O�z�:���x�s�7
:��щJb?��ll=���%�,7��ʞZ��E�����3�g� /�wd���1��A�P��)Uk�~Ge����ˮ�'E�!z��Ar͗祕"L�O@�b�_\?ٔs�Z�������w�A���EB�~��$�w,��c��"z2��!�x������(�����l�Z��0!�ߤ�i���+?>���|܁ԎD��fi�lFl�2��L	���H�/A�=?��HG��R��1u���L����KI��* n6p�Ǘ�b�	˵�`i���XDZ7���C-F��_t �:���H���4r������ݮ�H��
�yN	~l�
���Ue������e��M�O������7Sq�P��0�T��P�#"�K��K���E�� ꚝL��x�V�� ����&lC��w�C��΋�ǕDZƓ�O��N?���,��D	�<�����|���V�M�݂�|9:TSմ\Z$���C��9�s��&�<�>[���uD2���<S)�yO��� �V�GEK�!��ς�i?]��W~��MR�~���'��l�5�G���:�Ծd�ܕ�A�_r��]U�%X	CIJ�w|Cr0	��?k�f��u�]:d�ݮ��ؽ�|ni�2|xf϶W����m��%XT.�����q��ü�fy�N�fDd]*�:� ��������0kH�:�N�9����*������MdC�9>H���F�Ife��O�*�~f�^س�j̲|�R���%bW>o�r����>%T��h����N�C]<[ q=������o��x|M�rS�A�4�� chw;FFgE�+'��Pgk��E�µU:���-�u�v�`{�W���)k�.�9�s����`����#������ύ�p�W���謰1- �4�D:�vsZ�~Or�vePX�]���cnvYG<��d���)L��Sl���B!@�&t����-P�{WKzC�Z�kl.�'��d�c�؜3G�[��[�J�޿)�ƪ~�B�b..�֜:���d����6e�z�p��Ҷ�J	)�R�U�����9(<v�6+V����2��i�!WՂ��yrϠ%� ��'���H~�,h���*��+��zAm2y[������{�L��s_T�Л`ls��:�k��#`��m?���p�K�3�N&��u���SWR�h�[�Q}���x�3A�#�����,tD
��Օa�K�C�U�㇌���zr'���N�/�e�FmK�yLr��K7�:/�{��W�r,WXM��M-�	�Uu΋�jdp�+}��T�2���DԻ�9c�}9�𙿁fvx�~}r�����3�]�<�r�y�9-{g��5c��y���5{RS��8.�E��=��v]�OPe�?��Y�
�u��4v��d���l�����`�.b'|/8�eN��<�J�@k�h�=E�[��ʖ����;?��W�� =�G��'�}v6������>;(�4W{�������mݕ�I{����/�k��a3�ý+�쪅�Jd=g()���d��O���;L�\���u�HҨ����z&�䩡�Fv�gV+b����i,� )Ǉ��ʡ�_��u��� �aT�L�)��	�^��i9��l� ��������s�CX��D
Be����OW��=w�[ť#�2�_���۪8��*��ͳ�C�6@ ��~�	�ԉ�q�{b�@�tB
�ނ}?�.��qD�=Q�ft_�x����w�'�����'Q���!��h
~��	D8ۨ���Jc�����������Q]w��W�$Ki�R� 6{:0$s���>�uem2�GN���.zF9j?X;g;5�f�9�$&�<�Q��������$jo?��="OKj��l��r�,V��FK�|Li��>d��|���Lqa�$�F(+@1�c�6�K�D�a�E��U]'+��/�� �}���q[��N�r��Gt��J9��bMn�2����,0Q�I(#&�b~��w,/�F ���،Y�ډ��줗�(�G��L����Rw?�/��*$K����'�b5SR>���e��L��ö��H�a��pA���yQ��/�T1	?K᬴�'/���Rh�I� �	@d0�J�u��e#T]���t>�?�»��s���
M��O��L�
^�s4E+�6y���vD��޽�������L���(�:/3��daUi�9��>��d*�(޿�Q���Ӽ ��;�W�V��F�qh49:EK{�)=�TȈ��4껨�٨�O������E�O-�>'Q���x��A�!�m�=fԊ
#EGQ^O�OFN�Z��:�>��gu�Ӯ���ۉ���o�tt�B�B|8�f�jWO/��"9U����hxID.�:�K�̀����m�A����{�%T΄��,_H�'
M�i���Y^���|�KLT4�{Ù-n	2�;@�~|{zf8ry�����c��}��Mo����5k�!~�6�_�>�]���)��m�-���|�1�G��fB����P�1�v��0����J�E(.#i`m���<��ڔ���=�q[sˍ�W	�`o�d��O2}Jj!M־G�Qx�B4^9 ��C�E.=w�p秘�\�Ŋ����j���HM(�+j<2�-(nb�"�^�K�ޅ��+�+TG9��xmA�Ͻ���<-��a%I�R;~��8�Ik����u 4	4Gu?��[q��E�[�`��[����h;�������X72���s�BW� ��jՃw�[�)��$�����:��$o��`��[W�_�m��	�?�Q�_
���>���>���B(E��F�y�����n�[D^d�>�����}�h5iM��=��t�}B��?�[�#U���Г�Dl��=�	�U�g�@������#�,,SW�ac����e���߫h���gV�l��t�Ö�h�V`;v*�L��L��_��ǅϰRV\`�|#U��V�M�·�
���㎊k��ԋ��l%��`�i|!��Ol�óL������O���o@�  �n��a���>�;F����cn��tf��ʽ9`{|+{��_�v�ͽ�7������/��9��|ǎ�aI�6�A$7�)-x���#���2��?�qZ\W�!rվ|<2x�$$M�-c�Twg���Ġ��RmRMʁ'���u5,]��Ƚ`�-c���۬�O40M O��H��2 L#��|f�`d�Q�ۗ�I2��8��t�r��X1Qn�k��𡌫�����p����>�=Q���B����L��ɳ6��"�C	���TJ~#��嫏�jA���Z���9=l*�)�t��'ezk����<(�b��b"�Ex�����Ԁ�Z�kC�["��4{�r���ǌ�x;�3&r�)A��@򸆦7t�.�
A��l#2B{ϵ����e&���o{%�ۿQ���m��.���8\xR�ef⁇��vK�����浃��SQM���	c�P\�~'@xș��;Ү���V�ՠ�9���jɼE�]�W�lz��}�����I�uX髹��=\�n+��>r� �ٲ-�����Ԝ@s�>;���ֲFɊ��_��e�ȄAZ�4�Oih���L���aX�e	[�����s���U/ie�}J- dP"��|0d�3E�_z�#�Q��N�a�M\C ��u=�W��jg�F8�S	���Q�~y�n[�@?1ט�+�Q�`����B0�4����ml!�@�1���%i����ZlO��aH��_�������o5��{��V�S�h�z���h�.���j�E�:���]Q���--[ ��
�!�����ˣ0�`���j#Hu~$U����D�]�5�k���6�C=��q�����ީ����A��&�r�C��#m^&7j g�S�Ryz6<pG��L���Ki�@���E7\���J��T{ _I��.�	�
�_��gbC~3����[�2��%d�>R�4�i���������@*�f�>b��f�u3XJ�<vR�d*j��++*�~����,3		Q���Nd>�C��jpm�N��sb<�%ʚ�é>l���cv��U�$^-1�2 ���8 ~Hbrf��\�q0�����;6��{��t�ʃ�M��X��`�EYb};&D�������;10�X��+�����ȸ����K�b���.�U��"�B�n�]9Z�	;,4����*��L�I�u�K>���ג�k��T���4����oy����K��4�a�k0.S�C�1����ӫg
�d�g�@ZE���������~z �-�ljQ;���D���6�2�Q�D������b�9���d#!Mr�ɳ.Ɓ!�ўޗ�BXU^q�a�.=����ݡ��&�tLr�����yI��d/�?-��{��u�g|�r�^g�4x�\ǹ�0�H#?���S��o�27�ͯֻ�}`փ���ڄ+��Q�Q�M���;�S���8��V���M���Sxt�KU��Cq;�(��+�i�g�?�8�D�0j�R�͂���]������2�L~4!3eon�|�9:�����|�NU\�h���1�˃I�e̮t���#���}���M���*/a.�&�T0 �k���0�������r p6~;�-���N{Z�^���^P��J~.�Ny3�̧o�S�ߪ�P1�"KE���u��	�ǂ�����H�|򥁘�C`F8�P���߬�b�e�]p	*�k�?�x�r�6ه8	9P���"Y�����d+����o��>����a��O ��(�`���� �T�)�]�"��S��4;��c��MC���j�a����
���\;�p����H�y����+��:cZ��+Uy��ݎ��|V	��,���<�=׫��o�X3	oP���C$5����L� ���'!<O�K�s�>���7��4�~�PP�����8wl��,���f2s����OR5��wJi9K�O�cH�\����媍q�]&��5l��e�~�󽷚�^��@�a��f{g+�n�`�|�w�w��^����n�Z\�[�Q�T{dB3����	L x*�
�o}Q�]�3�'T���&�� VdWYWf)u�mĳj������L8�j�Ն-)��gh`��ƾ�3�
���
V���B���E��$����������5���G��Z��/��-��2�gI�+w�`p�D�/��r�1�\bҴ:�?`��\��O�ڽ��v\�w=
��������G�$dp$�e���}������S���w��5F���1⹸&���y�勥�������/�,=��R��W�}�;l9�0��r�g�9:#�8��r]jwV\u]��OǶh�Re�4��N֊숱ěͪР�2�3�];p��w�2�W��_74 �t�?�!��QEH�Q�!�ޓ���xa�1\��,%h�γ�:��!tȤ�(^Mrǧ+ ��r[�����xzQ7j��q���Ʀ�f"�Fs�D~1�p�VW�������՜�+&[��[��LN��4 ��db-��iL��0�K�*RO4�!�FsJ"��r��M�`�F�i�.C�������c�5+ʼ{a�_I,-��^�����+?���D��8�*�� d"�߳���w�*l�snV}v�#�y����d�X�]j9^��j�Y���a|�Y���~����Ox��B��J�{,���ث+�f�L9S��� u�u;�}���d_
�,���k�fi�a}B|A&b����i�{71m��q͂��s�)���u��h�UR-��!�ǟ����"����r��d:�fVW(Q](���T9ED��]h���h�������"5�'��+ћsvֹ��N��� �`^�����iV�ǯ��{�>�0��SZ�싌�H�I��j�EC�����/��懆�M�>�A2�r8 ����c����եQ���3������]X�C��Ƃn*0qlUW�M-a�=�f_��%Z_=�I�,䔔
jI�g��u���y����N�>�Cr������F&)lK�	9Z�|��ؓ9q����w�a��5VXw����ׄ��6����F��e��{g�l�+:�(��<R���E:ݾ�^Q�}�si-���j;r4\��l>?7-�"�)I�Y�����t�m9ڎ��,Ρ0 K��[�f=�>�BH>S:/g�W��.����wn�_cj��F��l&?it�3)��;^~�L�ه�"��1!Ùj��$��7��:w�6:�A
A��B�\z
��ؠAk4'��j�բ������W��N{����yQ��7f5��4�R�I���W�ma�TNW�3ڱ�W�ϭμ M��{�C�+,ɣ���b<=�g��Cj��g���:�����IL=a��Ô<�c��Lϳ̖Q臵쳪��MzU1-��q�N������g|;�T`�Tz��$GȒ(43>m���S�ߚCN���H!���Z;pt��~U�r�*�sjqi�v"\�!f�x1���`�/�rJT��&C��S�'���<x�x�3+Z%-lƚs��q�k�6${�=��e�U��V���'D��J��f-^����௘���*�y����3s^��ahX�cF�y������p�M�~� ��F�W�%:TV��{�]$��)�k´�2�_����>�}��N����d:��
 $�9Z뮚�F��$�����^�\A�
�2!��ރ]�B�1:�&L�zsL��\�k}g5s2Yg3X �,uj4-�xXK�����Or���=��qUO��j{���Bل+��\;yyZ/�&S�%�L6�h78,�uϟa��4��y����KOY�����2m8�;��7�ZϬ3h�%&DZ)B��e�����/���u����x0N ׫�9�[��=1C���+o %��X ,
vEۂ�7;���*�Td4D����:>5ޞ�*Mj���"��}@���Y��|��G�ۆ�&�9�����o,ʟF3P>���p�b�0hp�ے��qs���ğ��Gj�W�����FG~n �&�-`%�8����j�ީa#A�C�Ѧ��i��+e��qA.��>��8�#���&�ʆ�3��`�O���L�� HEЩc������!��vo��c?Z����"~��r^�9gq�:�464�6O1c��w�vD���2	P�v���οa]˦��'���c��xJ!��綞�˫
�ga��懎E�=j�W��}W�
Q�%��wyyH-�\^�h+�.ig+B���C�Vu����2���Գ���͙�A�z�%OV���tmѝ���Ѥ}�z�V�%���;�n�;�oj ��k��6erxF�C�f�ӗ�bv]˺@�t}��תE�8�p/ $)��>8�p��{�&�v.L-ЧD�g�J����z���2�q��B�A^�b?��k�e�(���ѡL,�cP"3˚����WWVe�Z|'�`j4Y�lL�XJ�>#rT$��Um�I�^=��;�\]f �+��¡����"}�a`�D��0�T���0ra���s:�8��ϟ�_�j�(g�- 3��,X��o��]��ia�@CW�&������n?a{80 d6�J�ap��1Inw5��2��]~y�1
X�U~C� �T��m�~��������ZL�6����&?6��<.E�I���B�O/�h�k����iU�J�?!2j�|����aTX�\��juLX���"��0�2�ꫢ��'�}Lx.�Ac�H�E�W꽱�z�"5��NL��,��$ew�T���!�\m �q�P���9��J$����X"�(f�B�i�br!t�1><�}�v68m�xq3��;�h�z]�����[S�灍:�N ����Z��20Kx��QA�J^<d�<Q�;�ma)�T�:~6ƫ�{��8䡊U3Ӵl��P�ǖ���H6�] 	e\�/�'�YtnG��,��V<a�5F��W�)��}��ԋ9�j���!N�!Q����G�a��2�N$�\O���ӄ2T�m�0m�.P���RN�]�2��zB��{�2zp.�Yb�/��j�B��bB���:�_��%�9��qx�m�y�7�v���tz�9����Ќӿ.MWyf�Gjc7�������a��a�մR��׻�4�7�ĉv�ʚI�r�3�@�_��w�� �O�բ�	�nT���鸣��u�A��#��x��N#ٌ#�xmӡ2m�QK�= ^ �Ȼ!t�6��K9�e�)�F0z�����yIe��1T��i�Z���ϊ|<9Ƀ�����W]��ʒ����X������Ƨ�uD�j�N�#]��y��j[�~v�囍B{-��[��&�oR��z�߁�X����ri���!]+���Px�
C��qT��+�Ex �.��I��W�~��?�4����[����Ǡ��%�2�g�<��<�+��-i�H�d9��>hD�v���
`d�[���qU���1��XzDB,�-�L����ט�Jߍh]�ϯ60��K@w!;�+՚DG]�P �\��02�'���/&E\�9���<����T�Q8Nl=M��j�t�S1,1Yc&��Lć03����:�RSE�ڻ">XA���G�Lth%��=��#�0�����Í������a/b�8��WGxŰH�dZ��:�8#j����d��@F��;6�[כV��gd<(>�K�b�m�D��к���5%U5s�#OuQGb�itP��Y��/n��~�����&�/�:6&"�S�C�N�XIV�s�����ѫ�V��8|#��~��InŪ����0�7dȎ��?���Ɯt��q�~A��t�|�J�ޔ4��0Wb�y�ѝ�2t6��&���\F�~"��k��(F*�����@��%��aa{.��ǿ�k��<�>w�B��[�U[��mjؿ�L��mr���q8������{�d��N l��`�*�<���p��J�4%ٯ9�<4�8� (c�|a`Pr�S��6��]]�
pr2K'��K����C7�wӭ0E!�O������z��|d����F���3St*���'��td�c��j�e$�6�P(s7��):M�>3�-�yA�e��zEa.mM�}lj��TJ�09�z�v�T}�p���L(FG	�UJ���/:6L�^�9���n&56A��F�`�ވ�m�V�ȧ���~:ҩ�������5s��r���t[-B�Zs�R�۳�c�wѡ�[�< ��=v�C!>6����]���z,�����Υb�3@��
��^�*)�	H;�eO(�%����T���W�H>���20�Z����6�Z�qTr��x�teJ)7��v�c�r��c�N�a�?�JWE���̴p��r�8�Y��5Ȫ8/˗�ί�g�Eܡ�m���*�qk��27mB �>�ly�"םk��6�J��h7�Sb4���ޭ�s, �
l; �Vۇ���Mڎ��<�RM��{S�#�dX��\��I�6�E�o0�!��`�Z7@��Z��)��N����Ue�<�6�+��Ҟ/��(��c|.��N��±>������b�>@�o`د��`%�t�e��IiPh��!����	�,i�B�N�te�L���C�b\byH��!��r,Y�K�ݍ�/�)�z��p�"Z91��)q�áj9K�bҕ�^�.}É��Vi)%�J��P�Z�M$M�֩���f~���D�G���,.�Ba��
#��p�9o����K��
l_8�@u��4����}�xIW�J�=2yU��/>�P5�K���3�L�PYV�&�0k��<��)� X�TrTn� �C���L���$�� �}&ж-cU����& �w%;�z�-������X�����D(Q;�vn~;��f5�8��P��m�����F0�*,���{INB T��5Ҷ.Lx�����l4�)�4��f�%�00HB=�c!��Q��xb�����Z���4��) �8���=:bf�er���:\.	l�xt&o�;��܃��ypz�9@G�0�D��K�h�N�7x�m��g5��I����A.l��u��X�dV&�J��0��8�г�Á]}�B�T ��/��e|v\N��l�&��G����M�
�?Y���t������0���9�[ ��N�c��k�u�m�l�|�!�`2�njTS%����̊��9,Y�	����������o�,r�+��o�;���B+��5�*�>���7b��f��jZ]W�=$J#���Y.>Ḣ^�fT�^��,��`󟐳G���D[��2F)�n�3�]�D|�(b��c%�]!:X�I�ē0��J�R���d0$M!�ְ�I�����rM���e)�i��{?=pR2In|�O��+�o�_����d9d�}��c�ѕ���=��<��a�q�
:pgJ�ʤ}|ٞ��WQO'6b�6-q"��N�3Ba������X[�R�+=3�{��bι|ƪ��+D0e���$A��b�z�� Q�(��\�~����c=
jWw���u���r������{�2�u!vH�c]J�``�û��r[Mm�m�s���$B���h��\�D'�k3�������Uդ��c1W�y�䎨�	3��-L��& WҳÙ��u�khZ��6�\BY_H�|G.�*nm�`y܇]��ekfy�e������jZ/,=�;�x��d�0<׃����O� '���L4��Q�ݝ��v�H�a�I�R����d�\��.�&�b׍2�`�Ϗ�B*�;��s�QOj��X[R��BnrX���1;cp���Z�ܸ�d��E��+��0������5���q	�#��T���*���>IdV��.I����=9Ñ��vi���e
'R�r?Z�k��\��{u���;0�rՒ?�c����'���2���w���>�W��ہd�8ݧ��v�r��	Қ�}�D�ݽm�,|@�2�dCGO��u��^"�b�n2j�Q� ��yw��u�g��� �������]lu�z�ȋ���X0k\� k&�AʳQ(�(�v��)�$���-k��mcJ�5������6�����$g*�6���,w�]Rۋ����i�,����+�!N�v^������s��xjv�;�y��j`��o���{���:H�������:��5��9�v�7�`SV�o2I�3�t�)gg�fq��|��t�	��B�]v?��Ɲzq����"'�EY:�?��66iSE�(�\���o�ےq�%M#CV/&I�X.�Q��7��$}c�S�M�p����P��yr���!�[���#8'�1�ԃW%�q��s���AgJ��U�d��F\,�N�����)�(d���%_
�ui�t�7�:|�t#�v����:�ƛ}���>�
j L��%�rJ�#U�hD�kb{�9���#"�DOMif|ho���&K��ܿ|�f���I��%�q��t���G2Ӑ�5��Y#z���\W�Pd܍�a�)Ыi�ʚ��_��W��R��Ϩm#�8�2;���x�1J��5G��6{���)�vD�3�;e�w�m蓟:Q�#����dH���|Q�Io).�a\��	(�+D� �Q��!?cϐj��\UV�S�����@\�q%I��<u�)߽�~�8�o�]����rw+�����L�C`���DHzO[x�O`����rz~/ʂ��H�ڌmf�c��	�$�~b���e� p:�<kHVLzW��w���苚�x�5��͔����A���#l1�h��W�Hl3D�D6B�w��æ�n�'Ti�9��yB܏����)��\�j��`��q���vR2���L7��]0����*�'z���9��X�MN�SJ��6\�z�9����{����1 
�c��h 3 ��~��R��iC2UxX���`y�=e���8=3y>]�$vt��<W֘��^�KT�,^LhUٽ�lM�q�8t�l�,93.��*�O�HVԇ��zz�Z�<�z��/���b�P+֝�t/`ƹ��*�ː��`��n?�n� �~l����{�c�Z�הr��Ey�/�I|{Y�pOf��x�˯t>��a�Z�ʿ<�Fuk~<��|�#D�՜����L5�X��t_v�#4��9$�b����=�RF�tp��/�G{��WO�E7^&�U�E(�	K�ѣF ��6�$&^�-���[��a8e�ƒ*&J���2��V����I��C!��4f\�UX�u5K	��ӡ����)�)�)�y��nj�����P�PL��$\���7^��D�� ���{�r��0i�]���'��c��4�o�[ D�v�jT��1V��%�%uэAQ$�P�mJ0��4��W��¡�,���w�,) ����<w���'�s�>-q���t��^�L�}U��1؇� dz�<���;��<HP�XBA����E�	5Կ\�R,1���

���D
-�~�d�qE`8bG���}����[�C����t�1"Jʄ�Կ�Et�h�i��x(���
zm����.��>#�ge�3K�!��-0�}��d�j���&�ߑ�zN�b$�7�ף��
/�7˷��xQ@'�ݮ�.7<�˶-iU)�W�,A zB2����W�������g5#|��:�[��
��gr�#f���b�c�?�I���ynvKh`�W���1�}��}��<6α�\ڧ���Sw�Ԛ�Z�ց�\V'lx����t�"a^�	�B�;���h6���ϻ,<�K�U�:_k�,a
�0v�"O�Q�������
�5�{���]e�	^��Ap� �qT����Gn0�b�% \��w�n��b�nr���YQe����@Ԙ�7��$� Z����QSˊ��S�x���/����J(�P��(�{Z��>�K��N^&�*N�f�e� 	�0��nL���S�ֵz����FQp�܁;���X���Đ$+��M3��*M�� q�l=\�,�QjQ ��~pDs���}Ǩ��[��0E��)W������Zf�W��:�}"e���+i�ސ��lJ��Ur���10�?�T`w����o?���B���t=EJk�A�4F�%w�hО��G�-^������o�|Kj@��l�ya�*��}��3@��MD�O���pO����m���>f����PU�0��;Y����B�2���þ�V�)�5�^S5"�DW�����ϐ�G�8e�Yzp���%��+�F�"�z���'�rd����*3�/8��'��,��`{Jm����Ay~����0h���k8F��u��P��x��#h�U��{}
C�t~B�C��������
���'�.nj�%�DBZ��"���,�o�'&�8�F��AXX0Zu�*���CX�A����Қ�z=���t��i�@Bť��P�=��9Go���i3��^�F��;��3�d�UGZ+*�5�F��q�h-d5�����P�%/炨��j�f�8/x����z2��b���	M?�{��7�	*�C5�@�hB���<��Π�Ā :��;��c��Q~�8�lg�R�)E������J�6�ҵ��WB�=�*ҡ��_ɱ�xh�$ω%9��*_�VE�D�ޒ"Xk�ŕg��9S�.�����YP έ��ko�(e�����@��s�夒���>�@�ʠVz*|� �����X��a���
=N�����]��ŀh��,s��q����%�<��v7v��n�P�rG�����`�zZM��~�f�E���N|�!q�?��#�^&o��uQ�K"�B�g|D|�`�I��1�̊�NL=��[
�S? 4��Eż�1>��e��9rm�µ���i�6n�w��
�.�ϱ�\2y�J����Y��c7��|~ e�]n�<����k��&!V|���,�u�ԛ�U+�)�����Ύj������;�K�Xzɯߜd�o%��+&"\�.�˘pT�@�)�U��y��ͽN��G��÷�o��RR����7�"q��zCE�3����PY����ܰY�}��Ǻv��#9���\�#� W0�z�I_`�}���y��c.5?�C#Z�<�T|��X1�nT�#�x���O�hJ7G�nYz??�f����M�]_���j��(F:w
d���c��#5&*lY�I�ft�	�r��E���� �"�h���~d_BP����p:��K�-n�Q���eK1�<p8A�h²����T��az4726�ڙ�O.X��F�� �0�T]/�K1����l�ʉ�T����ВJ���K��9ue?�YΆ�^/����E)߭��5X������" hý0�܋uc����R�%�m�:I9��;��O��gؖ(7��1{}�^��e��F��K�i�Z��� Juw��XU�;��u]:Dx�����1�>tZ&9�EBk���]���}��z�N+�5Yy�V���ʹ��iJ�1-�Dsxzk��uN�Ms8�ɘu`� �o�H��A<5r�0?]�TNא�u�\�)���0���.����)���\����^�ا�`�_][A=�`	��Y(:Ǯ]ڡM�Vu�Y��ۛ��;�YԴrq!��^³�a�<����t��g)��g�=�!bL-��gTSz�����uH���Y�r�)����!�g��}�r9
��0��D^8"�}1Z�q�1?�W������-|�ʎ���垅a��Y�H�a���Wnc�	=�u���*��96 �ȎJD�����BLtf|�%�]*:F��o�\*y�"<)�Ч#�N_tc�s�@pA9���_�L��9�e$6{����%e����}2琘�
�ёȂ=|N�K�;�@"ڕv��Z���0�$�o�~P�kb����ޑ���QPݞi��q��d��{ޙ%��%+��Ҕ�M'f�4��=��#�f�oh�H���ԁQ�ۑ�qWrH�j^ߪ�IB@I�u�
JE�*3�	��]W� �b.�dUd�_�ZQA"�C��;�~S�,ɓ  �y"aʇm+�lړ �=3IM�k��ơ���y�u��9
�B�E�0S�RGN�x���G�q��b�r?b�.�d"35��C݂����ݣ�A��fQ���Sk��I�+;���i��\`�2kp}�²�p<9!�f&q���N�4�}i2�)y����O8@g��RK:Z�+�@,v�±�w��9�Zov��}D��$��'��4a��K�,���%�q�l�A`�F��<������uӆ�W�݂�7���1R�|D���HO��ь9� {�R��#�����[��|#Zh�!r�)�fA��|;?��]v���G��y �iK�\�)Dc�����M�x;=}�����Pu�ߜ+݉�C��U�a��n�%P�Yw�|�]�ӡ
my��`�ޢk�Mp�8�3 Ai��|dF 0�#'�����D;m�P]�� �!ebW��W�#-~r	m�p��2���
����'Δ~��
���+�zE2�F�h��>8YO������u�S���l��J%܊gF"~�We�tS'��a#�	�ང��(�Dd��{̭>X�X�.X{��U�����q���-�2�l�j�{�r��G�L�4�L�'>���I�cp�h1�K�65���Ac�^HК�Z�&ZG-eW���,N;ۂ(��FDܟ(/���_��k;۬�����AY±8����XJh"��ԿP�������F�^c�ҿ���� �Rޠ�v���%�_��6&;=����+'�8�P��z5n�"�)��&��~��x�0D���QK���8˙ɑ���,pA�C$sp29#�`�BŴ�XV��^S�������<�?���h�07��:O�b|�T;O=��x�z9�1f�i�i=p��t������J��Z=`h�+/Ah+6Ę�]��Hί�������4��5�#��ɵ����
=ƤN?Ї�<�ԎOh�j�Dۚ���ٛ#��	��l�ۻ��h.��è�u� F�N��;��Y�ç��Q��^8 ���]���`|�*?ȃ5�u��L�
_M�i�o�?/����[e�FҚH�D���\�Ӌ]@��t�|:Cq)�ϒ �K�B����`����:
�����E
-ʉ�ϫ�x-��+S�k��2t��e��g���ްȌV��c��q��Ѭ%���/Ll�]�"@�"lN��|���cg�=|*=f|o_��W_�c���k���&0�Y�Z�vIc������,���33.���Ő7�@E��y6���9�@Z[��	��1��;X�{v�Aw7"s9��ߋ�E�ˈ]�����F��LV�N%��)j>��Uk������,���1�w�m�MP��4�S�y���J�����M".�a8�.��K&0��������}p
�Kua�WE(BN���5��wr���~��$1��4ӄ,�߾~d؉��e䗂9
6
~�v�H���<�r̍��=���e�!��e�����0+#%� PNT��2��"�����813���������b�W�E	z*�?�qk2�꒓�*vb���Iˉ���m�8�Q�o�J�]�,�ܥ��
��'�n6}8:'�
��P_��	;Ey7�K��������Ok�ǄP%�v00��+7&&9B��rowJ�ހ>[���y?�`"<�F���ʏ�w�U��tsz��'��+�����H)��|4��y��x�'�^�e�G�˦P�t�A=��m�L��qB-%�5	K��
g-Z�f
l�q�w�{�J����� �O%�2�Q��]�S�ډ��R���dT�!!�$B�`�h�i�u��Ȁ�#�������eQy�(�ͯ`�1(�Ɨ���f�x�*��>�)�_�U{���'��r�#�����/_`�{ɔi�i>�_WF�%�Cs�����O�k��,�Y1�_J�����CXi�oX�85t@���#D��9$L4�����'%I{��]�rشa�Ŭ�oV$r�x���`'8N�*rY(��v����y��;���	�,}O¿z�d����'/yj�Q�_�Q������H҆��R�77X�
��>���T���/�I}��C1�E��ţ���@�y�F(��V�5�v �r���1������[v'aP�,�����S�bK��j���]��LU��1j���[r�ߐ�q�}vW���UY�ǜ�3�\�I2��:�#�ʀr�t���G�ą5���y�A��,�W��"?k(v�yhγ�e�AR�s�E���#��3�V�S\�e!^��0���hGh]�w�c1N����N��#�|Yjm�c��ia�<sf�����B`��፜F��A�w»������JR!l=�/I����4kI/���E�,OXS䐕�����P��s�Oz�4�s��n7xI���'4�ke��+{�k�z옅_Q�3�j��.o���g�]����N���q�a��2�,O�S�0�%0�E0�<�Fb+�0�R�Iō��	�`�;��)`����S�6��%d�'1Z���h�x������)���>A��Ƨ�稢��8s�oUUi'o���T��,M$k�O���B���T�^1l��M�V4=�o���|�nR��X����B�^�R8�H��d1Sx���X���E�#���nI���#��v/�w{1�A���[C��qI����`����W�#��-9�jRr������e�s�Q��N�y�K(-��B��f�e����M�_ێ.�8`z]`J���<n�nB�總4ՓCj�JH�ٿ��[�M#�SJ��,��+9U�i����>�H��#��{4�i�`��+2��{-�
�gL�A�XoGe�B֗���8����0�g���%!�2(_uB1J�A0�,0��?�<<d]n��lߡJ�,3s��%��B�$�yr�[�" �D���91�u���4aa�C��>�� ��hC�!��8˪�ΚKH4TR�C���/�I7�u0V�{H27�h�X�]��Ϥ���H~ 	�e�
/̩��P������Ss��<n���R7Om�-�1��ls�w�?5'�}�ߋ�I/�v�i��A�?��&�shM�<���X�B<<8�����h������ޤ"�I�l�-�g�v���rj���w'M�g�`��4�o:�jb�	��]�ﳠ]�L�݌�+G�K��p�ѳ���$��KMq���u�s���:*l����4ς*9�f����Q�`6a}����;ap�v��S \�XE�ta+f+(�u��PK$�x��u5P�0T,�䇦Ĵ�"�6�&�,�Q���Ǧ���YO�/�@�8,$�q����;k����=�U��E�OL�єA.V`��Lw7�Yy)d��4'jx.8w��c���[��;Df�BC��Y��e�ڊܪW�3|߼�D�{A!����C���d�Z�o�50�	ף�s�Ip%(Q��{���
@a���lz-+���q��H\��.�_v8
���6oru����/�"���7޾���	�N !}z�)��F�A֍�bo������=x-�'8֘`�d3TÁ�*f�mP�>���+	�ǔf���F�����9比Z߱C`���<�㧫~7@`(|s�����̱����������Z��������8�M6���S+p�;ė��?Q�|�	��>v�H1�y�$W��g�����3�+e;>�b��Rv���>8��=��J�o��)xHM�a�T����.��Dw:�@�J���p����Uϕ�c�P?Ċ� �#a�h���H���\��Ô�x��H�%��v��?̯��E���s�:�5e�N��!��N��=�2�a�0ţ`s�L=\��^C)� �[�p�?	��$9W�Z��'�WJ7Wl2�S5�u�d�t/��ˠ�b1ɼ4�%/�5���J���v{�|-t������]�8"ު1�״{�qeե�?�����kmS��M��i��(�w,`�Ъ-��a]�0�~�*�0?6A��_���[����E톖SFtG;@�����f����ԗ}HQ��Y"6͒r�!M0&����YKa\�.��S�K�J"
��?H���0}���`蘎�(�d��n���
��:<�Q;�Rh|����@ ��s�Q�y���3�^��W�b��Y�j;�A�؇�UJD))��S/>(38[k��c+����%�H�z�C����AJ�3/X`����.{Ar}ƳpF\Kϫ�3zBo�]
ˠ]S#��"�4c0"
�SBr��ŕ��!`���dw����u��&/�|g
y��J7�R�\��-v���i�]������5� &-z��\�rO*�V�ԯ�Ǚ(3mS��\�{���3��yV��^�nN��
l�C�zG�B}� d�)��ڭ\��L0��	��n�Z�,T�c��C1�e �v��A$�V�����L;��miw~�.��%�r|�-%f��������3A:�Q��b�0�F0M��j�Sr�F�����C�3���NAdRr�ci˵f�Z�ǂ�ġz�E}�,/S�'���D�L�Lm4K��?Q�9��Jg�n�E�U�6��f�%��#��W�4[���_��i�)<�b�{����+�x��	�x����ۛ?��3����0f��<�	M�I �����W�%�䔻3��b?�d��5M�\��7�����*t��d&��A��z~���'���T�M���Zf��c�2H6!G��=�4��v����S��+��<DV�r�y۾����Aaمig�h�P���z�OF��=:Ӈ�ÒK~�%pS���l3�^���6q�o��"���C��	h�(��#����9��Ȩ��J"U�|ڍ�w=��|\��sC��\@�SZ׆S��:�K��N��b�u0*���k��?��S���LL�_��Z*�Kc��z�:���,x�=�N�~�mXlm��W锋m~6Dq<t�.=`]�X��=*Ȁ�Hi<\��p��
��ȇ?ک��f9��t�[��)�(;� 2NWC�����/�J#P<�b�^<��oTИT�k/.+iU�^ȹ�2�?lX�y��/N}M����(��S����<��� ����wi=u=�g7pDa�e$�����Ƙ���J�̑�_0Q�{0]�elE��HX<�nR�Ű�!���i�q5NzF���{@9��72<�����,��K��\:_<!��&�Ƨ���;:�bcs-D�\���j�n��)����eͧ8�mQH�xb�5?eLݷQ��n�����)�v�Z4
9K�u�>y�g�'�9�0�m�ʁ(�������fʇɋ�l�}���>0yc��~^wc���Q�!��w��2���05j��w��YF����3��9���qPSƳ'rwA3���3�w`C1��ZA�H`3��*����4D2/�v��[	1tI`M{�_Fk�{	�]@��[�rn�W���T�����E�����8�p<��wy�р��J(�rӹ#-w-y��'����*	�
�A�zt�Ex;m%]�3P�u;��m��L�i7�3T��"�x��4/g|&�k\���r׿����ņp��9gB$�x!�S�'f�M�8�sX=�N�Z�X5���zC�TQh� �5�>j��
W�redD��<&��;�QB^�X�tJ��o~�{m�h�t���$L�`�)�b��Ղԯ?�k]�~�nq���BO;�}���Ht[4�89j,�o��Ԍ/K�de)Ǣ��4辌�%ʆOs�>
4�CCS�d����v=^a=P��"
VL�:��}�A�y9Cx�4�u�����0�X������&̓`�0g
��<"���|$�|����u�N�5�&րl����AK���#(^��v��X[����
�>�P\���显n����	-��t��Hsqw!�����k^�j��g�`�0�Bv�r�y5ǔ�"��*X�6�\���+OL���PUT87��!���< ����O]v7.�A� 56hC��~�V����0���4�ze-�޷��h;�Q�Ջ��Z����������L���{9��U�⺊7̻�:�@�U��mEȭS�M7�T3|���"�t#� [g&���L�	hc���6jR' �	�W����p����ⷠ���+O6�3����/Mư�&t�I�IXΑv:f��-�T2NMqI�s��e���f�&_����g�#��į߷ $G�s��s?[���`Tx��e��q�X�=X��\}>�m�2r�L�WI>��,�
��q`�]���O��ڄD�ݪ��<�G,�m���UAp�ܨ����� ��@u��(g��ѻ����)����!���i�߮V�����W��"_������7��I	�.��"�e]�IX��ЯQӎz}7Z�r����wNO?���M|GRDZ����/���1l�G�w���`�FVd�B��z����tA�YY�ı[I\	 ڴI}����+�5q����Le��Y�mfQ#i��6���1+�%�!j�N8�"#<���we9s�P:ۨ8����ew�Қ�I:�-�a�I��O7���7�^p��*�ߠ*�-�F�W������B�'a����T�o��'Iؒav:ZJ����#q���8�v8��PL��V�*YS�p��|p��Z�ꖤ0ܐ9��3Z�B5�����.ek�HU[j�me�/�F��X�~���_J5���؀��~�;���]}wN �'� �	�I�_�Q�!�θ���	�����)dLG;KmA���)�`bkM����8��(ν��4@��x�=����z�s�r����k����їo��K��*�ᢣ�t�����<uoJ����`�[�M·�V�U���h�_�	�I��Iå$^j���BQq�Lta\x$�L
٩�p��y+�co�*_\�LSs<}N}��fy�A�5Ϝs;��[4��ƥ%E�_/Oa��^��WzYN��FEQ���f}7��}"H>}��'�;���]巊���ґ.��q;>���CB�#���l�Iy��Xq|�Ы�7~��yY�v�����R��@EQ���0��(�H���Ȉ���Q~5	Ke� ��Y�����v�q�(���6e5��P~���� ����������T�V���,s*dӝu��fW�W�ʹX�E��|�4����aa�����%*�7�ذm����)4�w
�߁8�p���̀/���ʽU!���n-`!U���5�9)V[��v#��m�Mp�]��5X2��7�.�aÔ���գy��T�O{���/��W� �i�b�"���fo�"�AL�3����h"�����X/��������d&ʞm���_BR�G�)>;�.:��`��a��\ʂf�Wm��z�!�����F˷_lVJ̺���3�<��������[���1R�����0�|
AC�Ų���hvlȃ]�"���1���{�fD+����E���Bq��rH�#��3���u����"���ѿB� QW��Y��FV�x���O��o4�	���	5a+ީ���X�n�!;���~��N�:���%K$Q��Y���mb-5��|2��*����N��B ���B&\V��#gV))t'���P2Dn)i�#�Pz�c��B�6��ld�	JUx�3�U�[0
���zH��~f���A`rD#
^hu�4l�A�(;BEXg|�H3�4��<E��[CUUK���>32B޳l[G�4/���yk��e/g:$R���)���
��3�K��NI❒��w�7�l��s�Y	V���y�+�\RzW;	�0|��ەT�ߦ �S�����a�`Sh+���j$T5]�8ְߵ9�� �*�O$I��qd���43�Tp?�����]h���~��ȴQ���#$oZŨ��*;=*M�J��E��@�%V/��̃#8Ɠ�a��x�Ռ�3��ڰ@�ځ�is	�������ꮒ���M��(:�3rH��{�F�\��z�k���jE�U�
Ϣ��ٙf�DZךʽ�(/��E��gg�̬�YBh�֛��Uّ��z�?mi��o/�Y��K�'�\�ǅ��J:��ܠU�t']� .]+"s�K���Z��Wd|�Y�E���-ϖ$Rb^�^�<}5�w���F�����7�&:��u=�<=��V�kq0�!W�F���?ߏ,d����,Z=���p@�>k��-B��D���7�X�����ƀ����̇��*#����A�}�L�]`:�������"9�;g��+����5	��XC5EQx	�1�_j́\�xi�l7�ȓ[�*~�Hj�����y�[`�C��NO%�'��i���_NZ}l.3{�n1�a�'��X�baۇ;�O�z	�&�_���]{u�n	��n���gDK����D��p�W�>��� ��LEu@�9����WT�VyS/��>���"��F$�雁:�B/B�Ѐ�;�Z��-�O҈��m���ܺ�1�u�:u��$�#w�K�l*a����A E=��JǍ�U�G�K�^��H��A�ze)��b'NlT���ud�n���s�4���0�~�hʥ9zoz?i{Bm_j�%�����1��	ih��pz=�d�r���ڇ6��S���˱�[U|�l�ܞ"@������g��l�"� y���0n ��K�W��?DM��sr�0��`f��n��z�r��\�8?ـ��Y���и�ay��f�(<�;��Uxw�k�6 㹡���Z��=Ν��u�\�&�+�Rc�
�i"0�U�Y�e�9�aE�͟xv��7�����2�X��}�(�j�������ڸ��~N��1�g���ߏB �l������uDǛgg���#�7��!Пt٪�SH"�H���M�xf�F����h�m~C'0+����,qn�[�7.�i��(�0S��bʰ 	�=K�������P�cǳJp���=��>A+�=���B�@����÷	2����sN7P��ٟ,��0�����M�m���,<�J�~}>#r}�9��kA(?�A<�?�Z ���u���lĉ@),Se�4��Z�S�.� Z�M�fH�fa�~̐s��w�|Θ����Ơ���B���0}D}��	�N# M��dw*�E��}�E����5���R������߬p��b��9�s�1�N\�Ʉ!q�렭Z4�/��A�g��߮�x?Jқ�8��7���O������ɿ������
tL[��5�E�%���<E��vL����E�E22��o��#�dC.�pY(S�������>U�k	�O��q%L�TEĘ��a�ꌵ�b�W�.~�,����qi�q� z�E;=o���.A��Zc��F���D�vJ�M=�3�8~d��Yѱ�0)��B5dI�Z�����" ���f9��JlFM��R�[b��
��g�]4oY),5���9~����q��D���l��,
���/*��E�X{QE���f��/a����n�)�fu��&�q��8�y�Ntx2C���1˟��n�
�B/A�3)�Piמ"�%C���ee_z?�>|tж�N�tqh��<�|x�\d�VH~�@�(�L9L3��R��;p���*���}�a�>�e4�Ȉ�؜�'$�0��a>�	u��m��g�ݽ��)�������	{>���X;���U��A9���;;����g[�*R V;��ypٌv@��*�:����*��מ�� �f�e����ȹ+�Y�jV�t!���ܱ#�0.ɏkb��>�c�u�$[Х���A�'M%��k�K�}�ܠ��V�(N@� ��7�z�Gp�b�=Ge�b������f�ӷ?ދs��iǎ�5S�`+�O^a��/�O���#�rS�U}j����a�v�?��v'񽈅�)q�C����I�H�� �����wNp�<��$8���ŧ'������l!�5����A�t����deUt�2�w�v�����䢫���+0kB�)�߾ϥ��)�j�ֽ7��T\h3mn��L� %��VcO9�����~ȗ�/K��6��L�V_���_��mq:��N�`����%����$���^������h�s��^�k����O2��4�#���'+7���S�%LE��	=����9GtF*�N�K)h$�w�& P���p�E��}ۉV��K�����k����˼/���L�q�=*����g��e�A9�~��&t [���dfv�X����Ɵg@ �o�������vF����� G�rH��|7W��bf^����Ek�&�1�,V+�����DÀ6ǜl͛I��~Ғ���g�W{�U?o5��=�1	��?*�%k��(�a�I��pI�dDӗl�v��#8����i�p~�}�h������vŉT�/*ø����e��R����C����F�q@K�3�n�4�w$�6�����L�|/ĬL�����5}��9�ۮ���b�H�i�;H:�&�c�������-��k3T�!KH'P�p����URR��M�
ئ�OOs���Z���d|���в܍��
�vHF,��
�+�T���gh[�h�ƢѤX�4���GH��p�?d�ܯ�L���3�lSvN4�����`�z
^�C��'�ذ7�0��0�F��4Z����a�$�К�h�5�&�.�9�=Eª�q��?��c,2�Yj���_�u_�d��9�3ͱ�I�<�-�a��Z/j1}����3����0��T�@�1��%|ۛg� Rˊ�� �X˜T�u�c)��ܤr�����$�=қq�̡Ɇ:�E���6�a�v0�
��j��U�礛R��e%�Z���]��p�\Q� ے���.��qз�f��s�>q�;I����öp����"��X �yP����tʵ���el��W�ueY�_eK+t-���(Z�������┭�v��Y��\��]ə�͹�F6>����X��2�@������L�Fs،.�ӈ`�Ά裙E���c�QWVC]S�*wO�٧�x
%)�s�&�w���DǅQ���|�{���()�>�[
*�S�`΍!ć_�z�]˹�kB���0� �0~�߃�]x�e-���Ps�/!f����%t�6K7���Ps-b�!�=���h�[��"R'�����ז�6Rb�g�Q�-J�h#[��fG�{��c��3�V�� �4���������rW��ҚD��^]�i�L�4	�@x�X��,�����+D��
�6��X"Wb2N�B��_��mj:����˖�Y��[�����s�1>�b��J����.$DdF�?��?���,[41�šPm7�'F|a���֫(��]���M�J�t�nC`3�(H:*=�pS��H�;�OAr��Eo��*�����gL��"[��޽�����z�i�dyi+Ky���f�?O��
�u���6����۠�]��Fӝ���I�����)u:��l�
��g-M��E�T[���Lo��a�鴽`ߑvS?��I��7nA]9�/�6�#_�j�YZK̄ ZY&�C�����?�)"�/A�M��ƢxH{;'���D���	�[uvIؠU*�I|*T?�!�9?au�(��/��O���T��-ؚs���G�o�OeV��*I1�&�u����P�l,ֲ#��J�2� X~BYK#�;!���Z�_���{��R��/�*�E�'��ZzSnO��W�eO)�_j����l�˭�����*yh��?6��
�͗'���T��w��s�=�~��]F+�+$��k)O��5���ן�.N�AW���(���^i�];k�δ�7�%�]"e�a>(��fe� 3�!�����N-@�Zj~��U�=�R{�@p�I��B�[�3K�
�]�N�d�.Za�_�����I�B?�����z-��h5�0]�/g�P�����C����m=��v1�y�m����������l�!S� �.���Ƹ"M�;�]�H,�J���ڊK���:�_:t�[�g��r��!ab&v�fBkW����#���r��:I���!.	���p�>�;NqF���?��v�q1jL'����#BZx�}5G����Z ���h$�C��6��:`�WS�4�O�8��!0�;[�|gf:���*����Y/3�(����+��=TXX������ۋ�C23
�3��@3O/�}1	?��,@�,Vo��ңEy��I�w�M8�0OA>�Z^cH�k�u�ye�Xj��X���%���1��w����T9�R��D>�9�=W6�Z��Ԟd��T_��׷J��D{^��Q	�o:Q��02�-�B��щ"��q��u8�4P�sº,���
���RP,��|�U��W�q)KP�Ҕ�m�� ��A����N���w0Ǉ��[4�IR��0��c}X�޷���1������a�Lm�J��*��K�e���@�oE��
iG<�������߭I�z��`fz��%{���f���ҎnO��<gj
�%T��΃W�p8+e\���M��#p���,9���mJ�F�������-|E�-���ݕ�C�p��O*��b�Tz�ԥ�D���2��i�S�ȫ&U�%�ҹ	�5���L`G���;�/�01.͐L"�9PJ��N�q���W�N>� T�^��I���� ���+X�9, �@��l�o��݆&p�P���w�O9���� _�6�ff��*�^L��=��jM>�I�g�2����.��ύ�:�3%7J�8Z�.@F��x�=��%���t��F1�Wm"E�b��U3���l�S�%�ѽ+�mȨ�!���;�Q�}��wK�KͰU��n�D��"�h`>��
~eA̒�0m,*Ӌ_�j�A�7�!�&����/v���=�
��
'�v2��yj8rA�]Z������`f���Nw&�F �%�:g���R�T�7�:D�ὠI�{��^��xTB�T|
�3�&��1�c�/�zP#ƨ�;�;�W_7� 	�S�UqLx�`9���z���k2]��>Eq���UWw�O���Y�&ϕ~���@���M$��i�b�Bt&?�<�vb՞0,d�߄�'|�t���_
xId;aN��'�~�~����_����l�Ňz�`J+�1Lهy!�ۥ��&n�j	����o��)�q7j��ͧ3W�%��|?���D�פ�N���E�Z?:"j0�����  ��%\��/U����C�Hcv!J�y��	��N���o��HM���Iq�)=ᢙ��|2���e�MtMm:S5�C[�g��Ӌ�!ZF���:�~oq�lz�-FB��-�8 %U�gJ%[�=%)��.���?#=��e��}��1�pq�f4|��6��:�z��d�eT"�Hqfm�I~��������2ˮ�� Id�/V ۍ��g7��7zؗ��9p릵]2zO���0U�e[#� h�;�>�TR��%���� i����C�Ɏ����6hh5�>�k����z��(O��$4���D����S�;�x�w��A��U��Y���F���~�*���"5C�b.�q���3T��}��!/��z��(*�Yt��MQ��%h��q߮V��'F�r]H9��է׻����8Kr��V��	�L~۝@������l&�!��t�9z9��9e�M���y�}�ґռ���V"����[F��,��~}S|n4E�q�81�HژC*��#E�	��QΆ��d&�@��J4&d^�i��Jt�uq����v#oeӮ������m��æ5_8j%.�(ߤiX��ۯவ��k�X�K$I�#��	��X��׎-����m��)���p7���]��dZ8D��^�-��ȓh��ϟuP��}��m��^x�8	%�J'd��Ai:�v�
}S鷕x��=�jdt�F� G-a�F��+7伖ta!I<s±Mgb��_)�u��8O�.��mb�x(OwK���eu,U)���ǆ��L���Y�� 6;u~#VQ���v����qUA�0�k�H�X��Q�U�~%���M��1BY傁R�97���cl��������n��6��+����"h��X��9fQ�9ˬ*��NJ�m�D3�S�>4�O^dgqq,�sRON�T[�B�@���g�ئ�V-�9�={��rFj04�@��[�܁�3%}3�c§����j�P c�\�W`5���<����Z������9��B���nh��p�d.�}65 W�h����E��>��鹮�������'��]�d��D��O�i
G�߹�HQu�����A!8*�5�a�r+IlS;��.�c����a^��p��%ãr!4�h��C�]LL-SY�#�>��4���	T��8R��o����ǧ�7�� ��	�de|9c=u+<�f_h.8���9;
��䤗�i�8Gky1�}�Fv�=@M�/��C�������Cɇ<�'�k�.*�YF�*�>� T�}������Tb�1a!��#��3}'`j9���d�~Ma ��=fT��ݝG���Ǐ]K�e��@^���w))*	��w3�\�ʀa���&F�o����o����W���)����p����߅�-�%�n���<e@s$"`~���g7�U�U�bcO��n�N��V�/��
�>ɋ�������頋���8�@��;������?\>�3���@Ɠ��3��FF�6\�S�ʇ�	ZNWG�Հ�g��&C�[�WQN���u��5��KF��~��y��������O���e�b��@��m=Ryz�������܇^�ʄ���'Qve��$ݢ��A/'�~���%����0����6�&&���S�q��<�c	�t�'���%$ &��3B~�d9���A)��aם&)�u�ep=�z�(��J��FlP0�<׍����U��E��}M���.����^�vz���+�kcx���Ig��bј��֙�\���-�x��z���F��1&���$E�Vԃ���NFAC�^��蹲-��Ti6U���b��������8��v��a�hw���&�(��l��FY>Y�G����Y����QPWԢԵ��-
�H�	�	hίn�R}O@���$sq��A�`�'c�i)݉Tӫ��FRy�Lrw�j��O����E%'�0Y˯�L�����zg)�V����w����/�����'W�ov0�fU�"�i�>����7��f �.�ў��!�=C�"B$e�DK�q���bd>Q��������/Z���L�$
�ך�R��ۙa,��%Rr'�p��C�h�؂Y�����1�I�++�byp����}ѓC�<�ί�s�|�)�c�'!���uױ\0[C��,3��9��9��[�?GRb�7t���j`q_4�E��@��o#�%˟jE����E�8�QI;�j���x�F7���a���kI3 L�����Jǘ���Ȁ�x�XF���w��� �N����#���r��⅊S`$y ���}^��4�Vx���e�FU�xβ��Gfj�p�55E$G��_�V�![Q:鮰��ը���1��A�֎⽬����#���Fӥ^6H��'� ��|b�h�hU 3��w+O2���~�"9i2H�O�P>��M�`n��h�ī��'t'�)ԆÛL�N��X��%;Խ��r{�T��JEĠ���+\م�"���=3�	:�-瞧��e�����k̹XPZ-�)�]P���<p1�΂��T�	�/��α��I���r�G�V�����޽b��FC3Gmv�ÅrD�PR�d�����P�	������vϐ������� ���1$�ؼ�{.)F�ܴ��F�n9y��ys�k��R!��K5�X��\���6e��jG�]�[���E��Fǜ��V��g��폇�_�@ �+#���� ���N��(�/��E ����VM,�%��f�kru�����
��m�GyM�6�����+�C�k{>=nT_^�z|�y�[9qF��a�=J��Al�f��tHM�_�E�CdD���^/�͟*EFA���4]f�x6b��Ӡ鵚u.�R4ȏ�q	$���&�j���+|S�K���p�'8趼��0��iL�������z��F�s��K�m�"��I�1���Ö�)��@/^�'|�\MU�x2S0��!�u�BL�>��b'�Mv��]Ƙ�����8E�F�}����.6��㡭==:��;�$���Ld򴦖�d~�9ç�T���:���H�oZ�4�V�Z*�h<\?��[�8G��Of�(����#h�MP����HT��Y�Ґ��ۂj�H��dݛ ��Ud6\FYUam�(�/�')-fD�%�ZVyy|%ek��O$]��#�3��
������m2=�F���PC�1�[,�>�տ��������D�Mi���oT�6�|V�pٛ�D^�*��_�u��qq~���``��ɋ��#$D��2��-`�r��y�1��o��5���]�I���z����E?�t�"�T0����9�7w8����X?��mr�U6� b8�A���'T֍K��f 0����\s��[�ҜW%��I����b�a�w�2��~�f�_�u��~��Z�V!�+��k�m��MNQe'�����n[�kk�+�r5M��;ս�����h��!pr��Ԏu`��.Et��1����-�L�;�8�f~�S��	]�������>�8�d�D��M��j0�]^�tu`fQȺa0eu4��VW}�h\�[
!6{bD��PrL��#�׾腞p�ҋ;D9�j�+������%&>`Yݼs�ag�M@@� �S� Ve��+j���{W>�r<cN�"���[l���m`\��Q�~��)l�l-(���!B���_6,���@��=��X&�#�8	���\J�B/(��.�Ǉ,u�mBarU�����bQA���oi��",�YO��<�KE�6� �|��M�b�,+/,v�j$�ˆH2@��o�RѺL/��}˲�$�--��{c?�֣�|C���Z�o'o�;t&0c�IB��v�|��鷲lÑ�H��f=$3M~,<�LIN"Z�ȃ�-ƙ���-�f��:�� ����2^8\�o�}aE\՗t����*�} �F��v�A�>�}�(�t@�|YQ4liBc��P���i���x�5n�f�.��m����u��D1�y�Y�񮄖+����wV#�I^ɵ{1�v!�_ �i-�#�c�!%7�Ѹ�L��m뼞K]�Yo�k�$�' ��L��~�D��;�^k���,-�k�B��X9]`�CtQT�Y>�c0��S���y��:'�fT��{:]�%�l�u%Ξg���a8~�^�NR:�������b����P;��}KC|Oi*	 i`߿#�c#���C
g������ہ8O6l�b���J�c;�uk�W�@�t�m6���<&��Ƀ�oBx5/a�s@jB�Q�D�����k{�����`><�̉�5�?�(D`�^-&+�T�$��(aPV\1x��~�uy�B�g0�Qag������)GϚ]��o�
K�?���8ğ՞�`�ju�m`�)�I	Xiq���gp�4�!�!��<g�����nm@CUo������5��X�+ۛ#)��!�:��b��ہ��l
�JOq6�1��M��E���w�j��sQY%b<N�ܸXL���?�il�*���#%�Z~'V�)E��=�C'� �Mi�D-�yC��)j�N��zɟHs�����̽�tڭ�t����
x���E�yq�kq�aE��MY��lB�Ȣ3��:7R�&��I�e�"��Ï5~����I-43��p��o���^;�9��T9)����fނ��~��|֠lZu��3�Eh/���15�pO�$��gn�4���B���/!YA����xP���XL#,���n�п��x1��,�zL�u�uaQ�D�pg2n��ц�ԟe�\Rp�����g n�Ck�_�\��!�!xs��]��c�?�/j]�!qߍO3�_&�%�q���gAf@��St~�:j�Kr��`3
_�Q��WZK�
��z�����$�b�դ3��3�U��{��0a�Q�Z�Rjdĵ�0�|�e`07�Ee�Ɗ77���y.� iS�}ݳ�K�D-@�Z=�s8�>��u��[������dg��"U��@i FX��ް����и}�(�Rq������$Lt�NVf���b�E���Q�:�����i����2 %ye���}gH���se�����+|I[9����15�(#����~H���5��N~��k�DK��dZfP��;C�2$!x��������*��C��u�s	�{1�V�E��K>�\�\�J�*�4YΧ��o�j�`]����\ ��Dɽ:Ǿ��u�:����h`w$8�X�,E���w'vFiH����U�M�mI+�?q�Ģ�<�S>��L���B@��c9~��`r��j��1!��y}�Ҿ�` >����~}�o?�zL���4���LL��2���q�6k�o�h�A^�T ��FP�ӫ�~\���5DX6j)��g8Z�w;O��v{��R��g���$��raƒ��iQ���]��D� g׺�?�B�����Ds�ۡB�[����H���^0��^�C�q�ɹ�kf���������"<�� �j��$��_P�O���d�M�aG<ֱIR�V��֤V.�� kF[4<�*>�:��鎦���~d	/�0�s��/� �I����ޣ&�e�G�1�W���pޤ�J�:A�]Q�y�>��=�Q��N����d��
ۂ���yԼ��p���� ��j�, �Ѹ�!��Ä�`x�c/ϝ	:��q��� �+���|���<(UI-�>�td¢{g�N�L`�����]�|���Џ$G�t<nr��ϴ�O��!e��lwB5�8y�.�������Y�̋�Oՙ
?�h��RT<���jۆ3�dyu�|2j�)3��R}1�� ߦ�����y�%�v������?{S�&#5,���ݯ�-��P`���CĒ�*x�P��PN���A_B}�y>���%��_��.�r9���� w�d(x}�f�mh�?QE��C5o��=>��N�M�46��#���.��}Q��x�R��b�t�[k�������	���9��U�ml�ֱ-1�P0l�?�K�^-0�*���q?Y�-	�JbW�Sıv�愈��8�#��S��\2���;=�2+ޙ^kH",Y���+�-���y�d�Մ��g׈��oV���`���
RB`"�5K(9� �M�q�`
a8��yV��%��GCT���yy(�"l�j[c�0˞�v�ƹ��gS�SV�;`�ah@��MI�k|U��=���pQކ�;����n0�.�:��y?������'\O� P^�V�!��I��?���OJ|��Y䪕"Eo���{�X��w�����~�Z!�+K}��"�<�B���m�ls�A�WX$솯��ZS�S+��kN�=9��@� C�B}�ˈ'V���!�;�n�T	 R����� �1�bIr�L��s�H���� ��ќV??�p"6wQ)	�����1Jx����-����Q��SDm����t2�ִ�Jw�ۯ`4�"s���ӫ���������X+(^ �Su�2�Y�};�ҷn<'���z�q%[�����F�kAt��1���ʕl�Llq�2̽YW7ҹQc���c���p�g#�1� �=q��\�*�(��(;xrT�¬MQ��X{Κ:��x�i�;�$?�ߩ�2:���!��F<_��Z�u*C�mB����9.�KE�qo<�ly���P�eq/y�����me�����OЈ��KR�Nz.�6)����/���#��Kw��x�t7�jm砍9+�Է�#��T����-*u�W"���{=|fr%�ɪ'��!ҩdWjHn��g.���.N���5�������d�1W�}o��'g(��������N�llF@k|wQ�,|㓎ڟ�� ��ڜ�\ђ�\+�<�c�%�b�f�e=���ۊ��/��(���JLG����;B0�gZ���E�o{b�)"_�cځT���S��~��ΝFh����;�+*y���t���1��H�ϡj�Υ���^���%P^8Q���%�<Ǫ3X|�z������k����Ib_�/����<���2n��N���o+N�{|�	�{�)21��:�����w�bŊk�l�&ѿe� F"2�b/���ˢ�d����Z�ܟ_�n��akP�h�U�"��v+9}%�.ؚ:z=QK�@JY�s�h�z����|��5�K(1ým2&�3!���T��8�N��p$���e�z�cH���G�H�� .��}�x�������Я0���1;eIB4��O�%��Qt%���r2��%�Q_o���E�DF�����Z]�+E{�Zx�9\5��.K���JT [ϟf��&�8�'�&�Z����bl���U1f���]ǥ�r����p&
�b>����~C���'�:Ln����`�my�2�E�KCv�WV��m`���5�FJ+��sk�G�,�Ϝ�kݒE��-�$vb��a����_0����?�y����:�[]���&��o]�Ӑ�/H����r l���SB� ��m6�ya�\�e-~��$��7S��$�����%��[y��e�Æ�����
�!��՛D��΢*IM֍ ��
 ���g��nv��[����>�&�30��V I�������<����	��▪>T��tUs{��BA�ԎA�&c/HF��	��{?6f�c� �|��X�w?���f �I����)M�\���F��s�7���:�Ȼc��?)�
\�f�Y�5]��ɴ@6�f�d�z��~g����
�P��т�[K��'�d�3V����`"r�ٰog�����>��j�GиݰQ�����[�A��C�Ǝ5����,��z@G��R{ZѳI�_�`._�WR�	�m�����/�&�1j�!�֍N+Q�8u&]8�{L�.���s�ˇ�.0`��0S�q(9��� �6�ꉚ#IV�-���>�b:$|cY����g��9�-�4�{����B;�Ora�b���)b��N���bO�&S�堉��=;�J]��D�Io�L���/�݆r������̸��U��#,|��ZY����\) ��B�#��إ����O/��9��S�5�z��t��Ļ�v�ι� J�*x���	F���</,@������+��.&=4�r BI^�7b����n��9�F���0�i�D"{bx�����3�e�m]�(��;�������=	��%�	 ���ɐ�֖D����Ę�MV�l��P�v��v41z|yq���ց���L��М;�_�F����6��#���_L��􇨖!��d � ,O��7վ��s���v\S�?�<84��ւ82�Bw+���#�
f-�,�̚H_,��\Әd�z*��8?��xg	�G��Rw�҆S��މyKZ����:��m_��.`��*��:�K}NS�HK����m�|9��~ի�6����6�Va��B�1V8�ɢ_�OyoQ�*,l��A���bBv���G�+�8MI����<���c��@t��7G��w����[m�=ijUZ��R�Q;̇7�����^8�Y��QUоI�ɌUK4e���UA��	��A~I�"�l��{ysu#ȅ$�Yę�^+)���*��~M\88lW���$�N��KG�+������cv�G�����!ڮ =+��o�B�\~%'�E��V�M��Y?�mݍg]�"|O��L�K�e���������D�e\ͤG�Z�U����.P��zc``��E���� �ڑ�c�4��_Z����Y�3N+�\�,���Z�Ӑ8�0r"<¥��W���%�.��:@����vw�[xo��5�*27dC���QB_x���R��˰�v1�t�C�f�5݉`��e�%L�vK���@^SsQиKA�X�(��I�v|.nӌ'�_�Q��*���L�TIyF�f'�յq'�������X6.�'2��8Uξ��l��!�	�rd�{f�&���p[�R�Y�h�0:;������;�L*�v���+хV�f%pL�[z}�!�)���{���h���ϟ@��:��銩̣*"�rWZ��y��C������uQS�� �tV��.G�Iު���7���V��iU�;7{�!0_���D
e��L���	�.�I�j��𐭷{�y�=�l�֐���`vI�5���	L��D���W�X���W�뿵����M��R�r��.(M��3r4�|.���]�Q�^��2�Bh�������d���X�F��C���١�8���qb���xS^�x�ܺ�"&EEFIֻ<͛%��cF��!���CX'���}�߿�䴢p>@Ȟ�j��=U[��Z_"�S�\b'c�t�_���׎���0�.l���Y8�9�� B2_XN���������V_�#�~ZϴE�k�HΫq�@��RyZ,sV�0���0�?�i�#:� ��&�-{a�ہ*�v�Ǫ�Zh-�����,$юH6KA�s`f�<2�k�������׵�P7+/���� �'nWn�I��PمTO�-#f	g�\�%~ �j��Ѷ�L�w	�Z�Z���V!����D��3]�<�y}�����m�h�("yMU�n^ ד������A�y��2��4������^(ڲ�{2=����f���9W�K?�Fx��d����<~D��\�I(1���_������zLҭ����+R��[S�Qvf���8@�wT�
s�QA, }�YՐ��Ȃ�a�qp��T�g�:�I��ɼ�@��� ����Ё�p�}L���?��GSb�:aF)`��|� �!�����#!����Ooʑ����{����[-���Xd�)���:,�b)�8�@�Ԑ��2Ml�^���U����2X���09WM�S|��Q-oT�,�}��{��1�ӭ�0��m#�;�uD�TU��+�S]�#w{�����OB<}�k{��P�6���ԉ��Ǳn/�WC�&SW�m����\�!�}I['#(	&�&
��[�jV���w]�e������ħ[�1�e`D�m�2�����p�9�	��j�����0��%5<�~-����	�!�R��ˉ�vv�`�?����E5�ֱ���{)om�UU��U6��,��]p��U!�BS3ԦW׌7)a���3_��c17&-���4�j���"�Wn�p�U�Y0@��ܙ�T4ܘ�:�`�pc�� (RV����ǽm�����"1.;�%�hf|{����r�(��\@�}�řR��h��2�Q�;�e��.FB��6a�kk��^c]���CT�ᅄ���k茅nX�x�ԍg�7^B�r��S���D�����lSub��J�6����
1��L�
�qlӮ�$C�Ѩb�*ܞ�$Q��i��`6͑:�(�.���h�cW���=����1�w*qg�zp7���	�8��ߘD�?�J4�(�:��_o+|[�BZ������{��_���j�z�>��lԠ�rL��Ea)���hg���#�#K$���ۙݷ>\�-ê�H��4�D�f_�v{kF�����`�*�8�e'ێh]H�<FWA��dn0Sfm�[s1��wO�6�l��ZݚCѸ�2DUlt}�Xje$+6{[�屪#�Tg��.̇bP���yڞ���~��]G�\���0^)���)�z����!ΐS?@oN=��_v0Ȋ�"<�NL�2#��!��7�m{��)��x�{���@=h7�G�b�q��n$�H��0�����o��Q���TB^m~�����]��P�#���V�g�Cl��2v����\�V�w@➧,]����`���ϳ��v�C}��n2����*���X7*�M�	.����r�}j�64MB:�^� n��c5 M���!���"�n�{Q�-���-M�@4`���
�!������v��X�b�'��χ]�x..h�.�SE^'�l�+���3��<�'x���]��ţ���,����^�r��A��u�v�"��}�Zff{4}gx }n�>#�!�֙P��w�a��W��\P�'���x��\2<�F��p�����i��D�_���O(�x8��9!{�LU�&*@�'op�V��^�Af��i�%q_��ܒ�2<�y�Ju���Ju�M�)���N��4"h%B�LfQ�=�R��� uD��`�鎤ڋ��>��r�9�A�Dw� �H�R�N<�������&W�;��x�w����0q�QQ-����Q�З�{�jq1����w��vw��	�*4��ե,���f7x��޵��3��x������-4�N�,ڮq%H����Fv&fߴ�w���(�c�w�7\g��E�X���ls��g�s�6����~�^ǿ�Ǘ̝]���&�}��Β�Azk�"a�A�����qvG`(���:�`{ēB]�P�?˕I�(IغcE�Q\8K��/�:X�.6*�2�S����_Y��>a��y��	��b�U�#�����ji���56<��ն4�~��J�A��6�Y"��k����ke*��_�V.���{͓,�;��<h��n��~��z��wv���C�X`p���!�[L�4�u.�d~
��1��.hڝX�0�Db�!�؃��~1C	���V�6el��{�]��w3��~����Ҩ���l1|�J}�����S��wV?�X�A�J㴝�<�)Ҽ-�������h�Bןm�&���/݋[��fI�^��j{���:���/�KU��o�M]���B]��f&����F���.�`�i�Pv:=�3���Y�����"�g%\^�G��Xi�>]DO�*AU9F�Z���QG���(F�W�'c5�/2��SJ,�;��Z3TV��|��/��p��i���E9ڄ���^Y���d���^��\gy^�4`L���-Y�j�G���@�;U��%�������
��M�%d0����9�<IؗS��8�Y I��P֖��vEί��5`�I�VcU���Mu�I�/I���u|�B�܈݆��S�@�����1p�P㌌��UL��\�u!�o�Yp���w3��h�?2�4Ą�p��/�#	�J]۴9}�l����`�p�Q�YA�����R~��vK<5J���]�[-��`/9�<��O����Q 4�Y��������\&!�p����o�#��9y_�c��8�1N�uԀ�>P$��j�TVa|�%��;v� �9��&�ƾ�Z���٩��_�N:_�"]x-�j�r&��,�{�9t���q�w�r��iJ2���D�곀�����G�[�t7U�4*��D�� �UJ�o�ݍ-C��&��=���t��^%C@I�2�_mY��އ�$�B��԰�vt����d����&��f)B"M�q>��.�.��[3µ�@�h"��7)��hR�~�f;;�#�6�L�Ô`Ф�-�a�W�M��_�z,��6~�Q���P�� �	W��JP��'Y�[�dOi����;�0�� )���ތ��b�~���KV�-�|]��a/�U�8\�6��?���O/���)m,�A��{O��)���A���%Csm��Pa��0d�ͨs�����h˒�S+s)��Bw���|���B�G��Y���Jw�K�������1W����g�H�U�`�D "%�x�.7�����XIx$�Y�Q���9Y������F��h��v���񐜘�0��Lc�(ZK(?ii��&�������\�>� *q�U�m&���PT�>����@_оPx�T`@�����K������tփ{1���s9�U��l��m$�aG#����a;��p����QQ�3c.�d ��&)��V�C��L#���� p��Rmo]j����17�.y
Z�<��j]�Y�
�Hg��ss��T�qq����X�+H�\�{���*���<34"S�� ԟ�)��.�5�;���.��c�V����x	�e/�t�M������%���K�e3 J-�N4[K	:pD֒,9�i^x:Fsy�%���f��=�\X�M=(|b^QW���&t]���#�B��^]5��>�@��w}"W����]�C�G�Ke��?��8������������ؖڬR�'{ɞ�,��Pt���T��.k&0j��i�Ç~[��C��K��F?�7�^y��A���G�Y�t~��P���7�U��Q-�RM��G�Yv�ǯ����r�5զ]Cl&P��g42�s;�+~�jrf��R:{���M�ϖ�&�	���T�(�w��E�����ϗ�:��څ�CCg����f�
>��VgM�;�	>@R��||��|%�D�v���
�L����yj۷C�~1~��!�ꞕ�`�\L,�b\ W��L.Ww�ҮD'b�q
��=�0��Rx���TIV��@������*�?������ɓ��e�aF���so��e&��,��D�ػǗA*�W"��x��gN�9��M0M|���Ճ������s����}��Q�X��w��--+�^wa�W0onK��)qi�j���kO ��z�\㕪;oQ��/�D�Rm���d�W��ž_�A#�!�>�n[:�pH�^��!�G����o�X5�sD�Z�tՂ�
�a�A���,�nP���W$4s���56A���7�:a΁�r�rY�w b��J��V���S
�:'T��������ѹxW)'����J8ؒ�T��q)+�Xe�����?�3�8��g+o�7�b��zP���Ҙ�����,|�"W�!�0�'��Ν�����~��%�����������ؽ)̛v�g����wP��4��T
�)��(9!j�wVL���/�t��C�g�k���3؈�_;�@ �'�p}h��24�d.7�h�(dĀa:r6[�h�<z2d����C�? jV- �ru��U�E�|k�.?�n[�9������#; �=˂3��=b��*�2G(�[�2��,8��X�wN ��3�h���鞋�!�6!��r���Z�V�݃,e臎�XU�Ze���C
C�]���F�|��s���*ĕV��ڸ��}�pM�����س�0yx�F�\�`4���F3�ܷ
r_�J� �m�-��A6�I�jHܥqRU��T_����ގ��n��L�n�X��8j�7Ү۽�L{���(��1���4���BN>��?l�U��@u�C�J�5+zm�%+��mKK�+>�����Bm{���:ӛ�Sy�$��t��������/:|^M��������p�y�mK�ʼ�dq+�I���cY��h�AT�6/���Ӕݾ� g�VZ��m]B�I ��;��sHo��v��њ0��ܕf����Rr�*!_?���23\�&��G�������rD3p�	�U#8"�|��-���"��C�vx��p��B�Gf1h�����\W��L����dtM�'xk�'�����2~�V�ߚ�~.��b�FQht�V��G��/�p�T��/ɨY4@��ó��E��ݠ���0��K��f�L��D�K��u�g��N�8�X�,��|�����E�S��w���C�v���)���J�(+z	�`K9�������'%IC��F��{���<7����[��jobm?3��eca��5`�zy�����o���0�S<7�ǃ��W9��`�ɹIx�H��v}�J9�yf��Џ���KTt������W�Z)m���[�I}�5���J�Q�F���m�}�O<5}�ٻK���U���}	�^ړᦥ����E�Sdg2�u�Z��i�v��-�250'�{�LF�l#��r�^�(�r���G��V���/o8�p�OKpl�s��=]r4g������є:�hI)�_&/�`#@Iݏ)�R���Cb8� �3\�VZ�R4� �H��sC�1�q�iw������N�Ү=)//T0��;�6FFw˂V�����i �b�t�������ވs@8�\_��;EO����%6� �	h��iƊ�n���l�DLxz����g�<X�-"���i��W�����6���t$��A�鐲�C) آ2A�p��Ӛ�9[��I*U��KL�v�,m��le��x� ]gj�
B�~z%k���0����-;�xrY~�G��l�(K7����K<p�����B�L�B:}k�V��=��Nr8-ŵ���cN-ag���<�B����3saX �ș��v�Z�
�*�]n��wʘ�ϳ���"�L18n��u�훎O��:�:_��^=�+$��(b�yW�Yd����E]~5�:�cҽr�9mF?�H ��r�'�����l�w�w�<�:��uSH���o�ۅ*�YX�4�0l\���	�
�A�+3����
3��|�/o�x[�<�$��" ����'�i7�'�޹���`O��4��qq��j*�[
��ze�>����TȀA�GD0S"* Iy�
�1�:��FSb�1H�Ŝ�npv��r�� �#X7+5ݨ�n[��Ĭݦ��=/n�Ķ�3?X>>� ���d�q����-�l�^Y��w����+"�5H���C_r��9��("�E����}��|+Qh�Yg`k���x��Ғ
Fe���\�!U�n�T{���lu^�l����_~ �zZNj�Bm�9i/������9�D�|��Ƚ��R8O�`y��VF�<����LY��X��cd�U�l���!�D�cP�+F��,�t�eiW�2��	 X	�ѷ������o�sK��N��Sݔ�՗U�a�~�!�傝zH31�M�����{Ҁ�.lA��8���k�SZ%<=�����%%�Ǵq@��u=�%���r2ke2�6un0�f(-����q���b#��)�F.`]lƕ��i�X�	�>�Ұ�R��6<K�_���L�5E��	 w�^�/�"��TL��	�˦�������B�`��u�Y���uL�Mz��v� �¿�
Z��ە ����|d���+�޹)�eSE�ȇ ������:�-;�0<�J>�Rܯ��7�N�y�����I�>IA���i�����HP/s�R��&��Qҽ��Ov^��L����*OkX��ɖ�C5�&Q�1���S���\��K�'&Iݶ�h��H׷���\'k<?��5���/���\�sȣr�e���=��`�IR�)�9県��뎙=��G+]ϵ�'�[�^v,È�B�iĈ2D��(!i}���ۃ~��G�q�n��k@<��,��8or���{�<tK�5��Y�SuV�,�'7�{]Zn��Bv��&�*�hA�k��
����)�З�ڇ˅!�2~E�C��t|��%��QR1����>Є4�|t ��d�)N�)�\��1)�b�,��פo���l�F�0�^�U���n�,Fx��w+^lq��C�!�Mϛ^lcC��k�7t�C�ؖs�[C�/�6xj����A�:�����|0�!����!�w?+�+�Ò굲��ms��:��֮B� �^�0�bMA��C{��������~�d�I�_*.�i�N����	|���0E��j%��b�lg�:����}�����c4#.IAֶ��2��c_�D���S�9�Y<5�{jl �cU["pM�<Kޑ�ޘR�E��Û{�8Ī����40+&6�Ŷ�D�%���A%��;��R���{���6�W��qȦ!�cQpٿ���s��S�F1�8��V)�9�
a��D��ɛ�K:��XV �'IE/��[�؆#��#)�
0Z�%�=�8F�9 W^��?tT������r����j*�Q7�3�1��H�@�Y��:[�EI.�&����T"V,e��T�� KV\xĻ��0�(�dI@ox��aD�|"�����H���{qx�n��A]'���N��A�����fʹ�wX6řz~�x���%
�y��6&��G4vC����G�m�*�ش�����+)�le���P,�}B�]�Ń`��b�����P����Z�����]�)h��O����\��=�j�y�G�9OeQf�<=h����Ύ	@Y@�Bڞ����6����X�GXo�B�|�B�yQt~K<7 5�T��P��# �?�y�S`J�Y��P5�/�
Y�n�ڗ�4�:���,�o�M;�X�5�N��i�͚"j� [V��cM�X7�3=��1�ZQ@L���� ĢlKwP�F��ڣWd����B?0��n����"�?�::<�x�-F�<*4=�rR[��H_ӧ|��BC�v���� A��<�b�����ڂE� ��,9�n�eg¯���`P�ؐ��2e��d7/��aG'R���� i����]�&R㺚��)�r���O6G
�+l�1�1�g�gT�Ьf�MY7%��&����^+�&<IlĬ����)�iO��(�>�|���q�&��i����	s�(d{�0y�V�𭙟�$}N5o���=o�я�N5���j���'��B%~pC`s�*���Ӷ��Ԙ5����҄I�H�����J�PV�(���c���1�Ç.�꣨}����S��kd���1���4�g=ǻ`������~>�T�U5�L���±��wE���T0cJU7f%1O5'~�q��@Ԯ�^��ʁ9�\����> %g��f#ê�c!Bi+��MT-js������DsMcCU�Jr�����q�y�.c����d�w�z���yuQꮅ
����m&���������Y|����w�����"*:�����Е����ە���?��MO�����># �t��=Hr����؈�	$J�74!���Û89�5Pp�O�3�l�R^�l�����P���h�!A�� \aް��2T���,�����ʷI�2�_D-����k��+�5��೑Z;�E��y�r�&��ú�Ks������zi�N�@��ύ6���X�XأtLG4�ၫ�kcwgz'�.c���ǌ�.\z��w1�6�Q�O!J�C毠���T�����:!���$�;o�8����EJ/�x�P>��'/l��Z:td��3(����c^v����֩�F-ThpGQY���y��81vS�7j��|���h�A���4.믰D\E��lBt2O�2��픝=��P]��q��#�Ѳ�G����4��-�}j�x��U�|1p�, �.�o�aHG��a�=u{�%���<7���>�`�|ּ�$�ݼ�+���݃��>�~��������^i��� D5���ǧ�������J��+|��ZĿ��y��/Wr�p?���#J�����z���f�+G�����Ͽ�.y+�V���2��?�t�F��!*�xxӺYtunDNN��ѓ\9	�OƑR�HJS&@�)��m;��*F��s������y�S�w�f��cr�;n��s��F�£�B5p��a������~�*�}I�8�_mn���y�T{T���X2?��N��~�7�v�A��P��Dp)�\�ɐe�� ��kX���b;�#���3_��$�������e=}�E�Q|Ų_�H:,Z�;�"�Յ��֟zr�m��}�L?��a���gF�T��4ڟ�����t�D�8,S�6Fo#�kWn8C&]L��C\� �V`�|O�/Ǚ�_(mP�p[��Y%T:�b�r��V}��L!}�pݗ	WS�`�K�5!������K�&�`	0tO��E�8�ʶND,4|� -T8��QM��epA�l��?é5�ц%�Tj�ڛ{��$tux��b�|`����8-�����NE�R�og��f�g��W��B�D��OR8��ļ��<���`�8��0��0J��d5��6��7ߚ�_��������)f�����̒��i��KPkJ�!z�ȧ�@E�"�-���Ƴ��a�o���ir,�	�z��d��Ph��#��"0���o�-	 �C?���뵸+NH�Nz k��H�0�A�| �A���z�׻5�7w)�#�ū��6q�^)��$t͛�SM�bJ������C����W���ZK��^��d-#�K�=w��uj����y2��P���ذ�^� �}�s�k��y�F���9�,�uĮ`�T�ZQ�TD�΋Di�yF�fhKie��*q��;�T{~�Ѷ��1�*.@Q��&���pٳ�٧�~�qiVU���(�A0JD{�8��Xš�L�])�����:u^?������e�G���u<���8�.��[��@��]�0���/&�Q	�i��C 	��ApӾ���V\��(P��C���ie�n�ڝ��[��,�T�X���Ā�M�F\����d-X�aѢ��#��o��޼�xK�	^�;��9�^�ܥ۞�k��  �A�u#F�>�Y�]�S�H�%��6�5u���(ڿ,퟇dZ7��r���w�I�Y5�F�A���n����x��G�[쵸K�'��VFTD�N˱���:��Q�A�WWdW����<���f��lBm�l>�6D��R%׍�h��z�)%ɢp��(m&ޔ�����?)ve�[W
�h�� �j]A�^>��I@��G��'���e�����+����fHcZ�H��Hy�0Ïq���#"5d?�@�� ��*�^�ډG�c��P�~��Z��u��u�*H�Ϻ``����$�ָ������j�0�Od9�25��|-|Jf,��ߏ���[ۣ����Ԑ���.�\�e9�1���P�4j9]��8j�nrP�dhyuY��G�8l�Q|�Ri���ty��,�U��M�G���])��h}n�&R��M����Q���l^TXP�Ll�2_J����9ICS榿��@���F&v��mb�ľ�X�,����
-�ڷOn��C,�����N��J�b^�]� '��
0���Y�O�ܲ*zb\�(؍�Fm�����0�mI��hhY@"4xM�g"Y�dE/[���lw�G3�'= n,�	ܬ������c�-������^A㼈/KT�t.NA���g�Lɰf��z�����2����6��X6Г�&��]����݉u���+�`�r��(Uq����S�rd���u�ɶ*L�LUӶ���������u���_ă��=�ٛ";?��*�G��N�	(��f_�;~ ���IY���M41���5/+͵�v�N��c	:�P��3����ׅ�j���-R�pt���*q\2."����� �H �:M15��+�i���\ø�~����]�z� ����S�f' 
�;��}n��i&�����戜Ջ�Arr�����)�u��2)��S�N��U��J�cŇ��bQ"JW�4�^xS(�X�Ra�݀G�ô�հ�,%+�O# �ޘ�/�[~w�ӊd_n��ٴј�۷4>�s�s�(=����:1���3o/��WU+.��x�?��ɍ=��X8����yA���U��(,?H��_�K%�O �wdh5�F;Վ���_�@��q��{�q��>�ȩRe�,�&��j�|iz�2��]B��YP��&�t�Fm�~t�J�'��S�i�R�x�E��yl;�n��g�H�X�p�G*ʺ�+�oW�q��F��
w���Qb�r�$�0]s�;�١O��A��$���݌9���[&{�m�|���Apc����V(�p�Y~�m�(}�{�\*B����3#��@�6�|�"O�>�.�m��}�����.����-3���~35���>�K0��hH;��$���D�eK�L|'��O��ԗ����o���P�����_�� �\2C��H��L�#���X�GфZ����yv�/9��#��;�󦏏�6ym	��p���)��*Y+�;���[T�Z�Y g�����7�z��{o
��(��ꂡ�������i��ZN���#��W*�ɾ��j28�"o�6i������u�9;e�*������F$`�oˬ��)<On
�1O4O(Gd��M�\'���ƈ\���\ȵ�l���Yl�if�O��������@�i�Zq��Ӄl�&p�ʚ�[��lö) �2�4	 6�IQ%vlA��[ű�.S�)����4�3M��`���J�F�0 �����	�=iN�T��wByU����(�;Z�䍅��2w�2��%Az,+���&dz��.ǵN9.�w���w��&p�ܑj5Jo�^Zm��l�x��Y{5I�r����bq���#h��I*������7Ƥ�VNQn����3��>����L|�+�`sA����>����2�&�v���.qS�L0���7��Z�/%�@ךfZZ/|;���4��+ܷ��� 2Aj?v���@w�p�Bs֠N�Ռ0���AJ���_ž���w{&��I�GE��Ǖ?i���o��/ɤԍ�U�(�W�*�Y�����A�2j |?{h|�
#���A6��R��Q�\�	hYskW$F����f䳐�����_v���Y�K�ÄrN�v`����O~8Xij`؉1���K��]HD"!�'3�k~��K��5���d���� 
Z�K�̨/x�^��f �Li芰�l�3�˒T  ��Lk9�<�[�ҎW��s�fc�"B�D8+d�����馏Xi��	������b���V����zڛT����]
^;�8<5��۞� �?�Y��Ĉ8���хO	��҇�N�%��Ǌ�ǁ��0@H�74�#�Z����7
�h{��hX}�3-f+}�k��@/��x<:���zt�8*���_¬~�\��ʤ�b�k��UQ���H�@I7@���U�\�&����Ma�!�Qo��j���9-҇���-����>_�
�^t���?�MK� ����:��*C����b�s׋�O��.����65��|�Ƞ?�D5a���t�5|� ��*ѭÊTR�UU�����N竪?��u���y��Y��^Na*@�;(ј��ܫ�c�lḬ��Ii]�6�v'�=��{d\LOM�I���V����N���?��J�͚���O���ꤔ��\�Hn��aD���7V��O�&�wA����~��)_~��qn{��7������6�E͇@����i� Z��!������2�f!��SNz�6�6F�jJ&]�*N����䃵n�hvV�rHU����ܬu @`����)yT�«L�f7�����Dhp���k^��\'��4�9����L�+9
�B�)E6S��a����vtif**�\�x��]ۨA������%2�>f�-E����U',>^��i�}~4�ga�H�1��%H�?n��®t[�/Eu���$��Fx��_{-�E�<�~���Uo�-2V(�0�J�%$�)�ﰝ�+�j`'�p��Z�M��,u\�$6��I������
�I Z���c���$�]E���!�Au�@����_�|3�<+�;�6D��еL6a. Gc>M���rQ�l�Tgf~�4ش�h�3�qA�:s�ʚxV^e��/,�A9��>Gl�v.��
t�%������˟x���@UFCq�_���,n\�e�չ�Dh0���W�#��	=����� 7�HA��]I�.�J{a��ü����s!�4Z���UH�;2��G���l�W�{�q�����M���P!�XM]��jX��F4��<�UR�/F��_��OY{��L��@�T��l�������S���7�O�x8���ߔp���c�z1����E���m�!��C�:ON1��O�s3����#�(E�qmWۓ��`\���.?��ly����<O�z#ҏE	�Ț�WaNˑ&�9y�*��X�_�e�H����(��)��M��a}_�YLcﾳ��͗��oϧ�_4��T�q�4��ũ48�,� POG��d��=mo�i0�9��fj��.���J����$� Ԭ Ї�#���:�6�H�N��u�M\��!CH����)Ï�ʾ"��A��/�Ԋ�O�P�E�1� Fm����[�����ƃG��>��Q)�u��������@l�؅t����"/d��9R~s�(P*� ��,�� �:j�R �q�r6�����2�ɨT(Χ�6���iY�'�2���(��x�h��`�5M�� רVf�gj=e���n�1ג��zjM�IZ��]Ws���.˛B��u紏w3�4����g��	�ֱ��9�F	$=o��a���A�;�0�;U���T�\oʹ�1ۘx���樓WMp$tȦ����7����ߕ�}��(���8̻�����Z)Ԯ#�>�Ș���Fb�/<|f��xVs�N��c+�]<K|M�W�pwMbF��mנk+��_�j���P�����*GW��A�s�sw�(!d0D8�?���ږ5|ƌ�X�ϝ8\��Nh�}z�\��xz�Fΰ��A������)ś��RA[[�ϯMϋs��6��&������s�;���A��V�_���(��K,ӟ9:Dj%�]��B(�q��G�u�f�ڋQ�]��v����o�j�ģ��>2f��m$�n�e���S3Z)
�G�[4R��=X�@7��ꕍ�����_	z�%�U��wJ0S��x�5m����y�x �G9�mn��%B�5�'�����EԱYY�|����wQ_�ǡ�PB���#⓰Ym|�}p_�~0�0(f���BJ�,�)c��Q����Oj��H�E$�mĀ��~ˁ��)>��� �$o��UYGb�6��q���5sݏ9��+�{@�-������a�q2w }��%N��#F�'�enѤ��lJ�e��J�����92υ��vD��oJiB�W�s�U.�y����1�-�ʾ�/~HG�� ���Ű�3v��}����.�7�+cQ��C��_��C��Xd7Y�b{�(𾩹	�G�gy�I�����U)qkK�K��e�6����ڒwQj������[۹B|�p" gi�G�]�܅'����C`��t,:�B��6���Ei�fb��
�t/q���Ҽ"3�癕���5L$(44�n�S��t-Ԥ��+�Z�Gw��`DlNA	�X�~�~�yƴ� #��9���C�K6�	e�/�K�{�7!G,�r�k�6�ޙ~����H����r�G�qn��?O��ݫ�4+�^TD��r(��,���%x쥒>E����;
��[k��;����ܡ�r��Cz����蔹W>��٫�a\���5�j܍8HU�n��nU4��I�IX����yJUt���g�{z+�uв��zۮ��ɤw��R�=';��6���&� ���dOB�c����\�oM%	QT���c��C)2K���Rm�CS��;�3����%Y�HM_�a����*":$����$��0�`���"�V]q���V m�m�g�^�6�sA�#��f�oI��u_�v�9W�]	���B6w,)�R�f��LЕtȞ���EC�_�o^��ͭ�}���"�Y�VB���tDɾ�x�Y�U-��B�6�l&�X��4-�#�_%ϐ��e��ܫ��B��Nq&#���*2pv\U�y�;���ŗ��Wi��*R{sU�*O�(>�;-s����5��E�����c��l�ݔG�fH��Z��!]���+;կ"��jc3�Ͼׂ�ZJ{���{|�g��$�����x���~P�����5U���u��v��4-������E$a5��MQ*�k�!�҉Ԏ=�r�`X܍�]s񄂖3>���r'$���@�Ijq������6��R����� �����{!�����'u5B�a$! �#�a����X	��$��y@����Q���˕�/�H�^26� 
��=�Tw��m+�B��Q7�)��ʹj�V��%(����U#(SZ5Ki��P)aZ�M
q�;�����.uwq�rf�?]Ԃh`��7�Ӛ.zO���B�I7U�m�����Ƹ�_��T���Ġ� eL��?��P���]}r�p1���w<~��ɀ��\О�(�⻒�tP�\�z4�ك�L������#�P��3�JTj�K08��+��@续�h&��PV$�MӶvT�2s}�-�c�w<l�.I'�5B���_\rJ��!�:>�^�{`��=��[�����EHԖ��w���7d�l���b~�`�;�̭UYP���"<&�g���'�ł3�==�f!�1�����7��oŔ'c�ŃJy����F�2�%�����^%�K�3i���i!sѰ�e��H�L���T1���2���Z�c�Kn�A������C�^#�X2�����v᪨�eυo[�H���� C��?R��swc�wn���- ��t�l"�Se0U�K�x������P��{���׮Rc���+"`!&uW�O��P���$fY"���R�ȿ�\�]�EK� T�8���\W����9t1�nG�։L���y�� ڂ�{bGo���Wٌ�Z��u�\s�>��j�t(]�U�"��E�6���b��&��{c{
YXHF����篭բ����'R1J�@�`f�(� I���&S� {����_έ�@�M��iW�e�O-�\��d_����<J����5���j}ia�h�ا�����sF�M/hF�� ��_0Y"i�M�)�Z��o�K xL�J�P�a a�n𙽷���D��K�4ك�A��DB���ſ�o���'u�}v����̧�q�Dn;e�p�A$T�N�N�y������DLe�6���>�Ni��zZl7�8))�D�Y��Ѣo��-_L�#Uv�DL���/6y���+@��T����Q�tl���I��-�) �/%}ocƮ�a��h'��"�`㽣�'f)�ʶ�1a�TBޜW�%���4^��~���Ұ�a��4�1�9�=]$&ݿ�R�Oϋޏ�ȏ}S���\�s_r��n�ٞ�Uۮi.ԕ�_���?a�?0�9����^����s�0��>T� X.���ũ �td�^��;1PǓ*��$�s����D�	`2e1�!Ako���wI��v����?ԁ�)B����0�n9��d�v����B�A&��򢒧=�Sx�,����}z����_<+;��c����j�:~�_.e����0v�:����W�G�r�=/1<'p�E��Z�A�����p,-[�O�G�L�� �de/���{r"�g�����3Uc�2���]%��(�9�V_"�k&Accx�=���̰X�D5f/�{�-��	Kw��;�,pD̟�ux�CN%b$�!���(����6�r�(�7����XL+4�͑�P���<*�P(X�Qr:�q	$��-�"��S�Vm
@*P���k7B,U��
MФ�O��n�N���Ù�@�����z�.�W��v uJ�
t�M�LVF�2ϜߴM7� �ּo1����o�"��M���nzo% ����f1����:U#��#�r7m��XF{�S��4j��1&*ǉ��Gv���22�}�r� q4H2����d����H�%Er��0�۩��|qCsc���v�\!{_���$��Z|�u�&��V�@��u7��=��Q܏� ƍ0&�]|����$5�i�w�}'dF)�e��>�!��ø�b�q��>���Q���*�	��h�P�_�xʗ��N�2#�L.�Ͽ#������6���X�"�[_0�7����,u-��W���K�sYd��n��{��������_�DU�<�KY�d��E].�<y�2��塲~7�<�U�؝���9o���:}� ����?���W!I���x����݈���l{���p3�|�/x e�7�!��5e�|��E�xޕ&k�`K�xxlT��Z0�#7��
_�y�?��� v�|3����P�N�#�`�m5JW]�$ly$��1<��q D�zo�c�/��;v�N��Tܣ��]�|�܎�M�C���������q��{Vk�W��C�ɓ(?ϒ�
p3f(�����6
��:�:Ⱥ��ocL� � b���h�G��Z�iB�����%'�U:q��F�	є���S$w��/^)ƛ�5L}��q¼�sG�$��t�x��ܫB��
��*����`��D�%�N��/S3�w_a	ʏo��ȧa��Q�d�I��v��{�#y�&C�E�8|�E ��3)�Җد'6�촫�74���cu.j��˘���\x�N�^c
J*�gD5����*����6 �V�T�%�ȇ�g���*U�"?�E�ӣ�F�RB����\�v'YK��LIR)�_<AݭD�L`�z:� ���>�Ȼ���n~FĊ��#ٴ���P ����;�M[yQ��\j������ߕ�!&4"	�B���<�y'����wI<QhB
��"�Ǉ�!�E�_���[���hXfm�(έ�Q;o��,��b~S2�﵂p��50֜]�EG�o�`ْ�h�J/|.��&k�t��c�	�?.��N�ط���X8v<S?:����1c�{׽3���L���d���V4�@�E�I�K�Y�|�>�aN���[$�}K��$~l��86I�.�K|�R��ts��V��3�狼�24=p��@M6^�qzb��@�6�������P:�f1y�?T�0�L�BvUb���x�mT$�-�H#����ja9a/�\(���Q@p-���F+\V�$��,1��<��}|�Ѣ�V�]�+q0(D��O�(�H
Rv�Q1!��nnZƏѾ��lӹ� ;��%�����:��|��S�U!>�+RHUsSSw�Z �pf[������U�މ].��(XP2kZtByj�x�02�~((�s�,��/�Y��1N�Ѥp�z"H�\#0�;X���#��B6VH��`��W-���ÿ$"��$Q*��|!��ti]���$�#���ˤG Q�zx��'x�:���8��`)��D�"#w��8���L#�}Z�1٥���ޙ�4󻠂��3��1�'@"b�����8o*�4༓��
r�>%BI�Zy]S�{5��vG��ꋶ}cc<�Wa#2Q3�:
��{�Lg8؞82�|(��_h������R�V�0�N�����䎇�9/w�[�|^���1Y������L���d=H�BH�-w8���ֿ��Q�����lKᨤ���K�Dzh�MQ���^�O>A1I��H���BW}Z�ص�i�[Z u 嚋�@��(Lޡ�}O�R4~'����#��&����#�O�\�����5�4�+L���R��\������1T�YGY�c[*�1)��x�"��0Ř�(m�5]6M�$�#���g���m�a��ԑ�}�A�f�O������˥����o�E����0s(���v�F�D|�o�n�MjF׃1�QOǑ�*P
t�)�Z�1��%cQ�7��54Zy�F�ص�E�Bq�?�H����H �u��\u���`D&�R������^M¿9`�@�PuE�s�r�n|��������I�[����h�8a7��%��=�B���`��3�."¨��<���K��,�W�ǤǗ�����qwH�@�Xs�|�9k�#�m��.С@���a0V>@1�t�P:}�4�^�ދ+�3�Vg�ߜ�:�����)�h�6�~Ա�^
���YZ�eu@���-�r��N��D+R���	l�"���� (��ė�޼�0f�Ȱ6v�p�a2�����pq���S�Т7*�&>���b��PKn!����-B����CL6�jm����0��+u�i�Q���ᖾ)9���J!ۓ�A�Pҋ5~A+XSq�-�ꓽ�B;aw��N�^��ߏ>YD������c]�D���/���}�0����G9� <�昞M�^���N�Z���S�jV[Z��w`s]?~����(è^�b]�y����U�o8l]W��U)[h{*�8F6�H7��!��#=�WZ��}x����$5(��"bW��T�n���4�$�����|5L @�6�|�!�,�%�]R���k$j��;R��9�!�e�� ��ȡ)7áV�ƇZ���Q��nuH�O��-}��F�KR��a5�3t��$��L��''�$YLD5oB���}s�薂�����𮴧�u3�6k/�Q@S����0����-)�ư��u-�]\ 1dci^ˍ%���P�K(�o����ժ.K����\c�K}=�me��wp��y;�	���Z0e�>;�r)Ϳ�t��8*#�QI��s��*���Is)�����'�W�k�S�փ���O̣�����t����'Up!�82�:�l��)�1������g_Їl��Y��%B�:����4$�l����ˏ%%��G6���w�"nу�
k�uQ2��̟ڳ���֯��:���w9�84�x�Wlq/���2Ѯ��G2h���)�}b��p˱%�3o����������,5��}�=��ƀw��pk{W��G�]Јy�K$�<�-��sַ�&��&�ous�+j{ ��W�z}'��3w��4���1�k��?�|?��S�P1����V]|bwu�e��3J��<��Y�<��������u�A-Q[]��X���Y�@� ����Q�Y���_4�n������������Ӎ�c�D�������3I����	���M�P0C4��b�$v�����Ü��G�u��(�%Z��E�ABu��A��j�{ue��y�A*��J���9�Ϸ듴��D�|V^�W���w�	#$��i�[�; ;D�?�9��|lG W����ö�ˢ��9T2SH��+w�X��O��6A�>�{���K ���1�[Rd¦kX���QJ���-{�Y|^��IV�Q{���+�$�(��ztK <�ڿBM7:�*��4O�kl&��V��X��\ʅ��٘h�@��#4�-����;�v�*/B�y�� ���8KE%`�4����x�'R�i��m��˯����Q��E���%���JAe�`I���oIA��*�8ʟ�L�qrJ.��;��א���^��Kq<3}d�C�yjW�Pa$������BF��B���M�E9J�}=ob�BT��\sL��� J%\a2"U�j�#�GR5�Lw��N���}@�:�c�nF۹ŁNb�i0I�U�5*T�+�u�Q���Iwa���<��!i5>䦒NSqj��
0��Z�QϾ9��xy�=���>zN�B��p�v�Ӟ���w!���&��b�e�٢���(�e��v���T����;�){m2�
�+��ԇi��h9����p����ܮ��wLSΣ��NgL>�TEb޵�!T���j���m��5��7XR�� R�+��9�cx^�$�Е�� r����;�Ι^�����QP�aF���]�}6��: Q���=�fJ�Rq���;S����*Ȅ�vݣ��	�c�U���jSKNW���m�>�q̙�V��*M>��h ^�m��U��;Z�8�%6G���J"��~�1\$��_�¹��0���H{Ջ��֗귧ۢ��5���.����=u�����l=:�c�|q6 a(ڽ�t�S��m�F��5�oҫ{��^z��u��ݤ,	��۠�Ȑ��~j�m$����o�ָ%����b����6����&�f*�]������3|ґ}�Uއ��<і�s}e:�=�V��2��+��j�i���3�CD���S�3M�7{�����*�I�����8�N<�h�t*vɇX�k
�3��
�)o��ܨ(�N��8�a�X��}���J�4�jP���LA��	�h�ށ
ҡ�J6EcB�R1����3O��D��<�a>6��p18(2$]��=f�x=��
G�%�wx��MԜ�5�,B	|���պ����i@��t��W�׳Y���/���|�*U�P �����"R V����	"��"�۞�Ӗ`��۔*vx�_C��`oj=Йt>�	�Ak�����ի�]뒿��-Pm�~=�k��}����S��J~�ӏ��;8gT�M��{PQ��t�?�Qdo�)���^6�* hYM�� ���}���0hf.WV��u�G� J�\��6�H.O|oN���+����1B߅���-Dl��a��+ݱ�
�'.	οs�
�Z�!s�Ư "�Wy�VO^j����%�P�Z�h�K��e��#c�8]^p������4�$��o
[8�*[���vP���F�V[8�ԏ�tl{f{�y�x�i��D��_	q��5 ��_�W�T�����8+�W 
纺���|9ֻ��N*��%?�n����O��0Xp>��0_��߉>(�P��3���fa	_o���or`8�$�T��0t�e�A����eޏ�n�b� ��Մ%�h�g�/d�(t�n�g�<��1f���̄n�G�Ugqd�;K�7/�V�$���hv��*Q<4��poK0[�ا-�!�V�tv�:�E�����ܙ����#�`c�\Jd��D�ZfLד@���U�zT
�?ԉc'7����h�CA"ʣԚ��_�T{�9�j�}Ө�s�����Fv�� �e�$8
�X�D��7\X�b�C�F��w����
��(K��R�����9��6�As��.|d8�Z�E�.�;�7�Q��a�{���=�&��,Y��>�q\�I��͇���9���� �Ӗ�W��p��>�Y�,��Y��qm"??��%�!��;�[��o��DY衋�����dÝ>�s#Iz:i X�&�����S�'j�W��]���JNBʙ6y���ʀ�q g1j�@��i�U^X·?���Tl��?��@��+U�H���2�pُ�-���Q�����st�i�����N�b�����D�Ȍ�;=�xb�a!Y%���ыAQ�#�r9컣v��Nc�h�_���s/��t��L��E���.''g��+���(l�MJ���4v8U,r���K�g���G�&/1C�oY����n��M�݆H�w m=*�hL���'�Ғ D�3q]A*�'�U�?��l W�p�� ��6�c6��e�"!|��@���in�r��	*�K2��c~{]ލ�V�H˘#��r��KI�b��$��g�owG�APџ{n����S�E��l$��("2w]f������-dB�-Ա{�0�Q�dA-�%�����i�3i��j_̜�C_�)@�U�K+C
y���4bs�l�7cW�'^,�l��ZG8���@�ʊ���{�ު���ٞ<�ѝ�ˑ�%з5�>r<֠)�mjN�]���s��s�d���K�X��۴`�Hb6�Q��^��t�o" ��c���<?�ڪ=I3�׿׶:� 2Z�3&���}r��h��q"2[W���LU�AFv�D��Yf�C$�ټX��Z�Un��w%�U�zJ2�կ��Q7A��s��O�_?d	��AP��K4
��f�
Q�`GX���o���:�"�Ź{ax����>J����6l:�%ckI�Bl��Yİ�U���zҝ�׏�8�>S��xն>�,�/<�BOx�pV�Y�[�"�0���w���;�1�'N�K���~6��Snԓ%	���Z��١��W�m%T��p`oM�o�����?������^����T��D[L�&�<x��țLT���A���l������+8����78�9���~70�6fjV�K���ŝ�o�<���ɗ.{S��;V:`�Ӄu�kj-����^��,���4��:��Mj�ho��&h�R70ަp��^$x=�R�L�N>��ی�k�������Y��#H%�5�q1#�5q��B�m�{ݢ[�i/~1;f�1U�+ `B-J�M ��#h���-�����I�j�/�b�h|
aMo�x01#�e�)����q��v_j�(��e�O)e�GK�D���yc^rR�_�q2����9��	7�u�U���������& D�^N���4*���ҍ�������ۏ�������U�������E�S!=���_��z�S����Z\���n%~�gG'?��b�<��d;ޮ �>O��E �����驼�z֭q��Co��!���f�B��X�B�p!*���Pֹ�0��l��F����n�zs����زTU��._Æ!�v�Td�� l~Y��9��m����J�y�?����lj�D����C �I|a����.�m��� �ug�([$�k?��R�k��9^
d��yp�~�;A�M����fDv,�q�����_a�W��<da�:�J�����6En�]](+w�ӧA����܄��x�;Z�G��@�����M^�U��|�D��_CV��^�8���a�Iq� 9��Cx��~�5���0���������O%�P&���O!��2ۣzB��[f��֜��#,ι\��+�*Lh������~��,~��_^v-�	�eR�]�r�w�2O�T繼�#g9�,��|@1����N�s4���ϒhơ����@)�(^�̀�t4�����dp|߿[�ۘ���O�/~-OבK�����Ձ!ܪ��Vg�C�^D2m� ��"*�Fr4��q����s��K\(���^=k�,=z�* U>�h&���V΅EA�'9�(o+�{?Ζ�����ӭ��q�{���!�]�MU:'y~���+�_�(��3k���t��PKY[u%<_���:�A�8�=P����),&N�3�	C��E׺O/���ʯd� ��q���&����F*�^�%�����cr������S�N�����	�_]� �S��@>9�}�s�v��Ե�)�L�%�}�\��au���J�6���n@�O��ĥ�̹n.�ʎ�]�#qQ�L����q�5-��Mϯ�4��Ũ40C<���e���S����^M��N	���`��Wn�[(^
�8����`��R;����2�9]$��n���ñuv�.�aʴ�a�;�^b������%함�0�E�f<ks���������˫ٺ$�����n��)��]�5�f�ҋhx����d՘�'n���9��Fy��[�և{���xP�d�q������?F�yQ��*]��T���֥u��*dn�m^V2a�f��T�ϒEx�Q7�e~h�U�xޅ}�m��8s��<���1y}-��%Z�457:��-�t�^�i)�&lD����� ��_Q}�Xt��!l"T��r#�քb�"���'α5̈́�Eb��������]rO��P�A\S��*�K��Q�����Yҽ��~L��s���ܔ�ҁ��BY�SH�0�~1C��v����������/�v��B��^���]u�Ϳg��/���1���5��%cH?�J0�4ț��b9INn�ϛRd�^������H_��67�g�C�̰��X·���1��F�P���u��x/������Щ���G`gT��
̙�[|g���Z�(QY_֯�m��A/})Ȫ#&"��]\�poo�=Z��Q�%��4~��
`�C��T{��=M���Y�VR6��d�E��T0l�A<E+,n�!��0����˶c�1�ߠ0�q:��G%<@�g;f��^u�{������sq���C]h��΢�~01�� t�`�
^��ҁ9y�CZ_�x�,�z��?�+��OE/�M�y���!�*��	L�Μ�RϘ׊�X7���D d.��qVp��X5�'׭�����A[/0���LIx
lfg���{qL.Y58������3�A��ޕ�w���&�BO6�(��c����U���֞Gi�"ן
��Yt�ݏ�X�
c���b�RT{Ў)yc�\���;�$$��Rr���yz�1��w0���b�l�M�}�����@$�z�C�7ɏ����pp�*��^�y��H���{4v�mx�֧���q��w	���]�������?��:�K��g�6e���!L޸�&W� Y{b�^S�����B��b�b��7��A��ǡp�-Zɮq��C/8���'����IxQd��^�� �1-5*F?�6�|�,��ؽ q�g/��Κ��EW�N���)I!�
,�J�S%C-5"�������d�� ��FH�ٟ�������Ϡ�V+��LmI����| ZTQ��]�����g٦xJ�"tͲ�2�_{>� 3��6�3��#%fR[@K���7�jw����Ի�'�X4��L�VtOޮ{�:�*��A����"\H
8)�s �G.Ԉ�qwRջZ��[o��Z�~�,��C��ɘ�I�vXf}�}A1#`e��E�Ў~��3�ōyú��("����p����_2nJ*������@�1�ۘ����⹷��o],����=�5�k5�N��{�݋�k����3:OHёəI���d�L����g��Ӈt�ǈ���G8��f��c>>�R3P�ج"%�ˋ1(ֆS=�.�de��}��g�-��&��AF�$"~X��|iAa:��*a�30z��?UH)����Oأ�Àహf�q��f�l�E��|��	��YC-b�CN����8'½.3�;��{�x4C�B -A�]�ۓ+6QpI��2��O�+�3���ʮ��@��|��9�m�ܹ���#vOc�7o��t��S�I�U�;M�ƥ���7���Boh��:nj�r�@˃���}ZlͶ� Q-�C�s�"��1C�-f[�R�6e�-i3���/��i`���W�Vc�oVr�wcXilX�C)!D+_���;�C՗y���]�L�~:GSU
�Ɩ2�A? 	Q��N�P���v���u�l���{� ��=����T�D+����ۥ�G�[�Wo��ժGum��؜��[����o!�20ż�7ےш��-H�3�𹯩�U�9O[|t�kʴ���0f�ԙ��]�J�lZN�X�awT�S��� �?PX�:ṓ!��W�*)��"vɭ?DO]�!���/1��1Tq�NV1OIܳ��n�������5��T*jo'c�L{΀|R��!&]�����`��E�J���&5^OL'�a1���\� aqly����K���	�l=���֧<�����.�����DQ%+*#W�I�����v��2�UX�2G�F�+�	p)�0�l�6�A��E�i��V���5ާ.?��E�q����HgR<�{��a���m����N�AiF���S=r�h!>��z'�������MJ|g�ַR�����dd(os��]���-��)�߀�]P�`!��D7"w�ˁ�vD��MVH�G���Ց�ኵ�k���y�w�ç�l��<JX>��2�:�Tz��\|�d�z��"!�x����m���#>���R�-���53��W��N[�m$'2	o�9�?�\������,'���3*�}��kx*�-P`½83���jT�Iw�cW��6!��/�d�yމEn�:|����d���R�r��Qf��G|�^�4`fj<M^��r�o��hb;�6���0��Nv,�:�����J#s�jZ3�(s˫�n럓��Y��in8&��H�:�k��(Ճ6gS�O����8�+�|�a�L31*6�2�끈
�U�-7yI$����V��&���f�G�g�������W��9Z�����+�RXP�B#龜͓c�0݄�q���d��&��7A%C�ć�l��^.�|���!(׳��`:��(n:�z���0��b0B{\�Q@v��4[~�n�����ܾ.��*Ȍ����N*h��pT#�Ș�ߚ��l�I�!�*�0Ӣ�!�I��F���@��2|I�q4W�X ǘ��e|D���� �*�*$u䥗͙}^B�G�*��qVIE��G�]��}�� ��Ajk�c�ҋ�I�`4�
�����-�x��?
V0��/O���D`����\��p�:���%+��,w��w�nE+C#g{v�#y�d���Hq#���hGɇ9��܀.w9A��!�@ړ:f��v��>½8!4��. �Tup>2�E�˭�l��!�"�lg�J��Z��Eu��]A>��)5_�
�p����BM��(2�I�a�g��(���@ˍ�k���Zbs�������ʍ��ļ�!�녁�����+xM��OºT��!�<c�f�b�,�p��{?+�tL�����s#<�)���l��|o(�Je���T��ۍ�($�����m�R�H����w��]W��� o��������U����>�(�8޽ǰ��|��OAnI����a��U�o��H�e�̬>aΞ~�Y}��H�"%p?$�#�9�cx0m(��c�+��W�?Nm}A&5VYe���� �l�d��+7�c�ْT���؞�ж�]&׏D�����gg(y�ذZ�7M���{h��Go��aLm'N��]��Y|���5��ʃI�<q��t�ꌖ�|���p%ԦM*t	��Z���/쵒U)gh\���ظN�0��-M͊�b% C����rn�2l-��}�w�͊�ל�<���a��"���D��7�K����A�E��`��0���V`}�Ц�\ˁ��t�W�Pkj
��n��mQ���((��F�^"�2�
�����}��H$�2@�aɯ߈�D`��E��|Y:JT���u+�Mp��#�(g&Q�u�vQ������?x���E_��d���7���l�*"[���6#��c[�� p_@��fo�&ek��ӑv8����8��;'��l(ױ�ƛ.7ܹY�+[����� ��ݝWQ�\і%M),}�	h8�����Һ�7V���Y�1ê%�b�#Ɉ;:p��L8��oߐh�����)��ɣ�3�u��bY��-��6q3T|>�(��N1�^�F\���Čc�;^�hLWµ����2<U��!`� �R����V�x�5�k�B3 �ˠv������!k��"SO�?��J ��v|�R^����}e�FȄ�d/�?�,��� 7H��#z��>����I��H%o%��`qST6�m��b��Z]�ĪF���1��������ա9*������Q�D�9N�3<��Bك���gJ1Z�`2�V<π�L��	���=�7��=zx뇿�b�9&��I���s!zt����N��fK����K� uw�6I
�����ԕ@
3���[�Ǥ�1�,]�F-|	յ���	�A/Sd��-}P�x!36C�e��d�DOa�]��*>@��R@q"����3���f����L�M�~W0�Z���B!�����@����a�̤doS��S��Е�v���'���GI i��7z:�d�W�x��ZI�(.�ۦq��B���nHˇ��[rr�m��:!�R�R��� =�"k��Wu�	��~t�A����5|x�>L�EY�2
���V�������+�&X��JB�Ů�lO��aݟ3����s���8��e�?�"=�}]��n���~��
]�3��*��=�]���:����6�<��лI���[�F��Y�� 6��wRC+���s��`����-�V�׺��U+���'���������+!�rYrG:R�����c�� �
����D�oO�N�k���
���
���AKs"h$��R�ÿ���;&���;K�bR�Q4���cŊ1}h�Ѹ������ �@|G�,���%�>�O���%����@yWo&��=����1=	�����$c^�����W��U�+ߊ�̇��z"U;�K�����mx�Ϭ��V��j��8@��
��O���OՕ�H$��b��h=�ku�)M�v���nSUU�V#�.
X�!&��}�Z�M�=���˫\?��(~F*n�����o�rHls�����?�d�L�M�|�6�۩}��\
�����fQ0fdM������������>�}00���,�a~ԫ0���+�L0�8�˅���?��`�ܳ�6�d�\KιxG��&!�^�Rg��"����I�o�~ۮn�o�\E�(�Ѿ9!r�,�� q@�a������W�h��-!F�,�C'��v�谽��/G��pr�߂$��$�7z�E�]-'W#���*gx9�e�P_��.*�r�Rd����_�g�7媯U�$�Y�������։�;�1���Vl��~�<�"eȺDys�je{Ђ����Z9��mm�:����GӾ��]�������-��&n��Vj2�/��T Z���8��شC�A^~���43fQy�+]�9�)�+�N����q7.��l
�V�@���r�x����U������;��^'�t.?|yW�*��������{���	th�~<x���
�%#��8l�+`���#q��� �	r�!������2�c�z��� ��a�	T�:�A&۫|<�	��P{���n]�y���}/�=ϲ�>QO9�#�x��	e����Jp�Ǧ0aAl��a>BP#��5BV%ב�ɆtL�J�k �t�:�"��s*�p缋��^��&'�[��Ϙ�Z�p���[��]x�`7�*�U��)
�ߙe���I���ڭ7����� n���`�	u�{�&�ʾ+�����P���L���>��K��5��8ʣN�V��d��sY��F�%Rq�٦������@�8���lpl�ɥG�l�t�ǇO�f�:�z?נ¬�u�i�v����4^'7��6(����e������!<��st�!�KZ�K���t�N�8�Ҳ9\cD�"��ث�C��W��V�7��?vfT�ad��=�I���i�%	7A�l��S��c��h�֖���,�	��r�<�'Pw���CM-�X�i���'�=~���I�_�D�7�H9�dv{Ē�|AgIq�� �����`�ȴ=�)!�'3A�= 8�hVϖr9��M�� � �f�stl�c6�#]�Z��V@�S�9�֐�\��hB�֌����� �_@׺��:V�^�ō7i��8�*R9�Qg�c �9�����K�a�)f-�����6�K�qyYV��c8d��M��5���u�e)�B�ٺ[�(i�i&�gQ�&M�/�]j�Lq�S*�Q�֏L����Co����7�k]I��}�Pvv ��{w7�ǉ?R��50�ud���Qٙ�-v����֩����!��ݡ�O� �qR	��T�O���;uA���_�E\�|�FN%��]=&hr��`�F���eX?BX���Ⱥ�c`�#9+k[S�iuS*���]�b�2�Qp����+Y�+/�@�/���ܰYjj'&��O��n��RO�yfk�7W?�ob����A�~;z���΍�->����|�����O'#�n{�r�Șl
(�n1	�-N�:��j�d�P-�ӄ�j#�/D4����
JI���U�,����#��´c^��{A2�\�ɻj��^��<<��Y�g��9x\�޽tm#�)���Z�c�*㔲z�Q�����i��ha�|�=4B+dd�G��R+���T��f'z&y�v��C�;YH����6F\��+X%�l:���]ˑ3���W�j=�XT�;}=���윗B��5%��jv+��tQ�X�.e�hX(��7Tk?%�8|��3�S��b����-�+:Ϥ����j^���������F�����y+X���-#�;w�<����<�I�FN@5'~�d<2�4��P-4�=N�q��F
��.�$��/�O����G��8�E���5gl�C�e�#ȫ��x�h��Yh���b�D��{u^���w��[��mJ��g\�0�-A��NC�����.i�z��H��v�j�z=!���Һa�n̈́�"�p���:o*փ{Ac䩪(�,qy{S�M"�&��!�1�=<'֡t〖ݰ^���m��YRo4*���ij6c9J`Z����ꅷ��6s��|+
|jUyc���7��ne4�3����@
hXt�9G����B/d	�+��B�.��o��r֒�����͌(Q����s؀�a����򓻍o����V4��<v�v��s�a���c�.v?�=�Kg�Qy9�Ň�<�.T|��H��˺�R�\j����h7mB ��>����9%���*4�)u"3
Jv�]g����@���,y���{�P#�yI��p5{e�/��&�
k�C�<�Y���62E�/u��\mz.	�vۘ<H�scGRcN�$��7"/8 ���#�����jk�q�f5ݨ�'�s���Ͼ�X�Y>$c�+��BO�ɷ�f�ܯ?�}�����8G[���ĈZ��F�����)T�I�~��1�nY3P��ť��U��:�z����`�ɴ�����L��<؟���� ��l�(Rq�R ˁ�I-\�q������(0xw��S�	��ޅ�G63N����S��p�:±<j�1�ꏒɱ�0D����q�Ù���A�ߕ`[���z���&�޵�I�<-$����`�	����5]_��R'MF�����G
����l9�U���ٔ�R�1�8�Y������+�Q�{~t����C��"܈I���kvti�BV�auyO*%�K�LC�m�n�d�^%��Y�};�x����U�_��
���N�[ǜzo��x ?�0�É��$���t��6�u�4��;,^VL�!�mO�����na��J�<xԭQf<���0d����A\D���MhI�n+sCVL>Ԯ���[2B��&6�?�|V���jXu~���=$Z�/�js+���Z�A;���V��7 ��6Y�J?����gNjx�J��H��}�io�-Fl�X�|U�(Ů4;*l>�һN��U��L}>y��;�/�1�8��M�ɬ5����[�֡
��o�Gh��ϩ����ήG��]FY����4��0sbip��$W�lݗ| ��n�pc�/!<�;V�#��7~��r�G|^@�����v�߀\2�x��Gl�Z�_~F}���AӥX�ha��T��t�ٞ��*�0�H+3�Q]iD�lm�!�Yz	����̓K���Ꮘ�N�6h�x�s�*���-Z�g��IN�Wo]v�1z��&��۰a�s#[�;i%{��<�����R3��0dL��
�'D�pbO���c?M(-�)-�[y�S�;�z2�yQ���AA�P�	�T%�\�`����k�<�d �����6q��Ĩ�`<����m/�lA�����[72#F��d�]0=����c���u�<oFW��'������K�4����5��1PV���3�<�v�N�7aDiϞg?�9���}�3*����D@/��ceoT�9twBh��<A*�ϳ�L����Ȇ�3��xʺ>��x6B����{)�ݫ
�Xv��f�I�_���,����hˇ[���l�����x����,�F��%���0���D���V
#��Yc�|ui�����j;	R�(ZD�u�RDpJ�|팋���Gg
e9�����٥���ɇD1�k{�y��A�h�Hd�iu�.j7����b7�'P�:҉�E3�����
��}����霺
�_Ҡ�K7�Ő�*��5K��:��>3�	t?C���5Tr^��w\v*gaa��k���a��[�i�	��*N#���S�9.��_T���D����o�砩Y_�~��ط��f�6�=<�Nf��g��@���<I��={�d8`zX7fh
�:��$��B���b���/`�{y_�b�8kvɍ�Z��?÷ 
]2��)V2��D��R��T�Οq�!�1�� ,��ǸSS��F�O���E��4�����Й^��m�@���:w�(D唟�LT>gp'�V��>����7�V��
P-���*��ع��@���xj�5�!�OE��$𥛁(H$�CPU�FT��l���O/��b���ū�Q 8�$��+��E��{q)���Uc�ļK�����/cٶ�K��o"_M������͞�w"���y�.�l�C���9��غN=�32 ��Y��R��I��ASI5���E���O\V<�M����2�&�.ȴ��� �ե4���N�W�'��(4% ��Vۖ(�'�=l��`�������,��Dë����'��~D^�`�ET�ٸ)��#/'�NL9T���.׾>}`M�ߊ}���S���Fcu���ǌ�샍��u�L\z�m7-2��"&wTJt=�]�M��޹Rh�����j��˯�@+�hu�j�z�̷���Q���$1�Qq)�J$b+L������A�2����g���x0}�M�"|��^h3�R.'&{
{��1��94��;�7�I����9A_5��a�X�W�!�:k�w6�&��T2�tS�A=5al��R�����O��d�v�R����x�i�a�Bל����G�?�!E�����<4m�b:E�+�,��x�G�Gգ��0&!�	-��"�~����Dm�6�'ޠ} >���s�{���DMr�����j�W�{\�r^Ǆ�i5��`��Ω���S�UJ�02"*?�_�=��%U%E��5(��ᘰ;֣��*!�:�àa���x�I�1�����r诶:j�r/�I{�@H(�N:ٹ�����T�n��+���c8�es��S�eǒy����&j7����' ��� ��p��m3B�܉���3 ex�ٔR)��5�S�&�ì����D���˨�^�Mr��sZ����vȈ�!�}m�������|��/��;��MJ��o|qY$���.q��NCW���8���[�)8=O��[�*�,�`M���>�U}���?���.�HsK�������nW�|���a
��r�W;�q�|"ߴ��*�/N^f���F��݋�;�'�_��я�Xï;WUܔ�����a%ƖѴ?�٠o��4;Gq�P~%rL��{T]���W+Z?񪓤=
�&ژ��DΕ
����ir-�r�G�_�Qr��j5d���e��
Ɛ.���,W�}��|��ALbĐk���j���w�k����Sb݌.��Fw)��ow�vV��	Z�˛B�@�U�=���*����v�C|K�+��<�9Z�����	����x�g=�4�P2��Fe5�VAY�g6��|O���x�ȢYw�χ�
*i�5�Oi���ԤwLOu��w�Q�=�~��~N_f'���	�Y�n����������V�N�dB9�^Er����ݸh�~H����o2��xo�0�Q
�$\�E�Ơ���h]��rl�F�%��-�3�$���"���D�{�����6��!���6�4v��߇;���A�`�m��ߗ�V�:ؿ���{MĢT����s߀�9q<wn��#��/B?�-���\�6���c�r��P��-jO���'q�BgY�9D��v�n�Ÿ��N��3�3<9�]��^!��ݶ��6^T��(��|6��ѧ��)eB%�Ҩ��QRK0�\��ԵI1�\D���ll��̷��6���J�q���<r݋y�(�`pd��i.��0O����6��F�x�ƀ݃��E�H� �4G⬖Ը��,R�RY�8>�A�48n'�IJ4G���G�yC�⑒ZK�s=*�V�~pj�Z;t��4�p����BAJA���һ��-傗5*�2��yJ�̟R�CI˔�d_c��B���	�RՇ#j�l>0�`�VZ���ؠ��"Z>��KG!�/VWR4'IQI�Ű�����*�����Z|�i�v"{��ѩ�5Yw�w�k6�"�b=D+�ٿ5�����Hy�t�����;��#�Js�ςs�^���O�Sk�Cߤ F�^2Rd��=�TL�� RN8�<\���w#�_T�c����n@�X�<�o��p��~�����,S�Оn� [�P�(1�"{����N3��,"Y��+g�y���?����/~�"���� %=��[��GB���c��R2�Lo�M�m]G��mֽ�е��`�Co�C]�0���_�C��L����n�<'	NC��9t<%:����T�}գ�oNv���g���xV^���a�љ�0ڑ(�#���?�f��.���џh`���a�K��54�j	��2Ƈ�Y�r��n޻�����|l�5}��[dO�!.ǌUs�T�*�{� A�Y|#��Ig�|ruP�Iƪ�D>�s�v)a����^4�~toS~�H�Wpiّl�BR�cy�x�n��I�N]p9%�]��p2_��ro���ʟ3S�g-)�CCZ�授�*y?�u�~�^G3��X*#��?WF��W��pRm,k"K�r��>GV2��v���b~����c���g.���0P%��N_\�+�~���:��k$X�����T#�,��Ī����;���uęY��(�Ky�`M�c��r"'�,��U�|x����v�LjP��f)I� �f��;�#Y]�� � �	�;SW������-�W�P��3d>�p���͵�����+;�z�~�1X��V�iCӍ��q��Zڝo�#W���;݃k#^r/�����vء}F��RO�[�O�d.�+(n�;iuc��xrf0�(X{�F2�X\���>����|6�G�����%(�q��b���`'9j���1�;:3=�vY�9��;zBw�*�n^���n�Wo���P|&{��D�*�j�0�n�gg�Mke����(�w�'�����e��@V�����Q!?�4���1��ml�s��?�I��$��̖����`%�E�����/�g'G���ϑg�T�%0�{ L?W�	�BpÔ�n*&���9y�)�ǟ�/B5\׾m�<jF��w��=|ccؙP z0��B�Q�ne�uu��넲�aP��F8���0��1�����'��8�"I\JT��dRl>٥�_�1(�qu��oo10��@m��^�|Ŀ��Z����b�Ψ��6���#�;A׾���&1�"�R��AtՄsJ���g�F�0���\*
���G�@�cH���on�r#)7�ٮ��h��x�����>,u�?�%.Б�q�O�k�H�-�/��l���l���{���\��ь)���:q��O4��DvQ��̏�A�����N��ҍ5�o�ب�5UP	5�`V*�i�m��Q+�6��b�w�"Rg7�o}��}_�E���7~GT�q��ge�hܸ����M��.4��$с@����DK�����9=�T%pQƖ� �E,#�1-5�D���i-9yb�����W+�
�GHm�>u�+s�xO�hcr^���22i��i���ʆ���c6u2Lӂ�^<QaŅ-�(ȫ,;��iw/�he��L_�MH_O�\F�z!r���� }�5g?���$(4�w���o
���-�dBPY]l�t�k�@"�{���EW,Tޔ�8oMɖ[�ŇX#q�ʢ��E��Kf&O�f;r̿�jk7�2 mh��v�Gf����>��w�����y�)g��a�m���Z]�ų20(u���H]0���Y�d[U ���Dd�'�bՅ�cq�B�@��'�є���O���E�
p�&Gޙ�A�'��Sf,�l�|\DΗ!Aށ&�՞w)�k�d��I�7�)��c�z]��fV<�Mr
0p|����@�� ��{�~&��0BLm���i�ᾱ,=�;����X����P�ZJ��2����;i��Lo���d�6�4[���P��G?�8��^A���f!h�������ܶ!�n�>� =��g��������5� �Y��4�|�-���q�o������M�֖~?/�HDK�uȦ���x`t��������Ŝc]�o���������Ly�m��l�Ȕ�B�Q1	<���AL� $*��.�g'D�h�ed��΢3!�� f�(���w���(:�htz1�"���ny������2������\�y�W�c���C���fX �������:�oq^�S١�b�����P���D�� 9��*�6�L���H�b�HMۻ�whZ�!��m2�,��dDU���L�g�
�z�B�P.w�cP>T,�C�]'�����C�H������*��a9d�����U�F؆hg�����E�R��A;��{;?��������&F7B�g[%�jhe��a,��:�;FI�j�G��dr�îp�3�	Lϔ�8+�`ZA-j;�?Z���|��i_�:�a���$Mte��S
�ȶ�s�0dJv�D�Yb��2
��������x�4�+�4~�N,t@	�A�~�~���2�U\y*�,���$�!a�v)�HX�%��جl���,���*(ۓ]�z���q*�:|��I5"�d,�	�KUP6FX��ar�ܱDlVuЌ�9��Xq\�ꍘ��^<ҵUH�������E2����9,�K_/�@��X	�S�"��7����A��\��񛒼�-����7w��s[��N��m��ْ��:�g��G�������T�@jZ.���ڿ.����&Njz���P�aI����D���>%��-�R,�.����Fi�E�\>X�J a�2@Ȭ�p]�Ry�c�[
���]:=�������h'�o��?�����v��)}\�A6/Q��S�s� � x�O�B)�:'�,�YX��R�VA���"l��XPv]�*Ҏђp��؟�xJ(Γī"�Ӭ�a�R貞y���ArMug~��>
���$!�?�		��d�{�<�N����DG3�rxm��Ǘu�����S^FYZGq�Y���'���6qD:��pU���d�D�d@c�Y���?e��4l�㺻CAk��> �������qE�9)E����� �b5���,O2*I/S����K&ߪ�o+n���.�a���8��Z9���G@(�T+�,�$z��p7��v*+��O��A��X0�m�g���ǚ�RG1�ʥ���΅s g������p�ug���E�G*k���Ssu����)���u:(����
��#��CT���񽌗vv�v0�b��p��S��/��זF������V=�Q���@z{j^{ٹ�;Tԥ4�w����]y�D�
P!���Z��ޗ�g�����*�8ۤa�;4M���p��i3�E��DU�,�:�Z��<
뿹��@����&u��5Q��(�=�z?_����&����ye����Ȁ�z���n�4o�P�;�ZI� ��,vā�#�o��'.3�E�S�J�{�d_:;L,�wR���X����͞��E�]'Og	4�*M�@r&%GN󀂁Ju:�(� u�s���ݙa&���W&�flCB-�e�|?%�,j��w΃����6C�y&X,g��S���k�:�y�
���Wv �
��8�y���R6DI��S����T,z��9���"��:�h�����:M��,�������� f�gjT�{sT�`��c�Gn�'ӊ 0k�s�Q
��*iG�����	=�7�D`�|׿О�S��U�H�$�|�,D�v]T��Y�e�&�R����إ�Vv���E�d��1t����.8�^b��cK}��?������EC���=���y4G������, Ӕ|��y� ��&����p�o������H�c_#Y���:�J x��.]�#��!��-60k�ZiG�^�d�r��Ə��>���V
�19q�a���que�z�D�-'��*ɓ2��z�jb���H�=�܄��G���8�?3v��R�o�*�d����Q�h/m�oF��0l]��rd�c���ܶ�dcew�̼��i�C���3��E��╙Z�G%���~2ق.�����G���j|o?7��*�4r�^��Fd&�\�I�]�u�k5>��T���袶�ӥu�af�\jv�\�cֹCp}K��I���������}t���؛3dU;]�6�Q��ɿ)��}iOYF �����h�0�M�'�}Q\�Rj�#�1��`����=rm��A9xgAk5ZZڄ|~PJ 8��c�MR�I��+���HV�ᇡ}��τ�}�'5Ǟg �kIo?S�OH��jF��]�@f�xu��W-�ti5�����Աu��I��J��T���P����q�o�n����f6b6�2H{�?8Y���Ҁ�?Y^�ON��#����Z<́��1S~��x.��5�hF�O�R5I�;����ƾ	����D]$ޜ�k�b���x]��CѵAi�֘�6�Y04��y'��g�i�U�;āb��M�i���4�-��v�	u�
Ta�8_������r2�
��`� J���C��`ϛ�붌Ť�q�:�"�d(J5I�([�/q���f�WU�?g,��_c��O�C�.ὓ�3�ҿ<X9~���x!��2��-иЦ/��ܝ�lc&⟷-��uC:�ù�Yо�
꺄ɣ�_��o���j�q�j��i��C��L�[��1�z���[��Љ��c\��]���"
�HR8�񩗉W��I�E�=�� 0Z�S@8z��W����g��6b����A��wۃ!���n�ﾎV.P[,Iw�U��w��Tti���V8�L�[�LVx�KVi�_�S����D	;�T)��\� �Wpg9�ZZ�Ӣ��,zzp�'�?���1��_	pc o�]�l�jT�y׫�"a#%E/�dPr�,��	�3<1�'ƶA<��|-�����5hD5�����e��HT��o���2�{�b�'"	wĜ/u�v!-���_�t$[7 ��I�E0��	l�QZ�?v����	 �����s��b�
�v�h��g�(1/;�[��Ad1?0,���0��w�K���Q��Ҁ��-z{|\_�uB�H@�1P*v+�r�jW	P��̊1^��}��>��O�E�h6�V?bV|���ҽ��M3U�#X���B��L]M��$XE��m'
�b�d�g1/ )�+5
��kӭ���B1q_����.�|��2A�U�f�+m�G@{ATɷLdN�@�<�F\�Z�A��Ȉ�����}k��K%�7%W�\��8��)3F�[��+'�vV�.��V�g�*�7���T��df��8׾p7�Xu����$ծO�(%�#WT��Y�0�l���j���];���(�a�b�\;C��"��O5�����k��(��3��eC�g3�~��'�`@I�%�����ʪ�;ܸ����"���F�;C��Ŕ�2���5�2Љ�������!� �K�]g"/��Tn��Sf�|4�sDށo�C!���\��w9�?M���t���SQ��Lv;�����?`4xK4�H����ͺ#��Po��6�E&��Qx�sI!p�ڏ@���V.A��GD�w��!�r2`E4��$����lkJ��l�QR�����(�K�����j��VX�'�YW�������@������R�=��%Ku�}��������ď�@i�L��W�}]�ּ{�8�q��\��IsH�5E
A���joŐ9���5�s��ܑ-О">�c��}9N�� ��+�پ��Vn7��*���m1��P�9;q�B^�/�A�e���A}���2��%��Ȫ/�k��6[��ҧj�4��w�+���{�yA�}G�a(�&�k�+�̑@oDܐJ��@DOJ��J���~���%��y�f8�;n�f�<,Qĉ�_�)�6�M���j���G��i��$M>-EP�q^�D�M�K��:��}ם���;3�v }�>��5d����� G���1�*=8�O{~t���?���q�TVk�6�E+�OK/��c1Ƕ�aj6�P�?mr\2��p�9�Մz�.\N��#�E#`)��v�4s����v�(���Ⱥw?�{;މ�t�Y]�|� �ݴH>���	�s #=���w�
ǌO��ھ���9/����(SͅHlH�E!B�Գb�t�3�����_8��=�|���_��wh��ذ~d��=y����W�nc��B�j��^�J\���)�y2�����^�Wl��2\��]d������ؐq0���!x�=u���i�I�j�9:a��[toJw�<�b����H�n�#�C� p�u�@�t�}��M"��q}@��Y�vzҝ@�)"�w��ҟ�w��sm��{�S��Y��F�h�/��(}�&���u���翠 4ZX� �ϙ���>�(�3�z
����"��j	o�4p���)�BOf %k��^�������W�'ܜk��d\'I�|yv��G;�:W��\. q���Y�/F��d?�B	f�z��Jn@��=OF'�i��i�X�E��+���[�����9&�%��b�����ظ0S�=����˙��<��F8�x��0�Km��,��h�
�}!k�zB��u=],������f�*�Jhs��5u��7e���
�h<?\��_'>�݇}P�ʚ�s�0��Ձ9��m)*Q�2k�9Nk���=B4�3f�pU���(�O��1�gy ���"�!ʔ����-N����g_�����
3����U|�vZ��Iȣ���fBL��k�(�'�m	r�FP��£�?��Ά[=��'��ilL�7B��5\
(p����	�s��#ݬUp�O+K	*F�3<	Z�o�]#̡�Zw��,<���A=N�Η=��B��Q��=<�R�9Ԣy��!\a��U|��OD�z��ЀtF S��"9��o�YN-�-�N\��Ha?���\��#s���h'�J$�#2U�JXQ�u��oN�a�Q����6p�U�r�
�Y}�-
�
�$E����(C���g�J��x��
��=���U�GR�����(A֐�b���3J
Y��ʋ��K�$K������N�}����׬S��:�����S:F8"?��S^��1�k���e��_T(�O��Eߦ��o���9/L�^�H���No�E�M�����S+��A=����j�7!�S)����������qF-���K�J`
����'~��Al��>�3ΓF�a4vB�`y�t�OJ����c�C��A.�e([dWk5
'�+�U�禩�kB�X���b1t�#��!�f�X?�J��Ұ��� �����\��`�U�td�`9�s�����������C��ؤ��J֯O�mBE�6@�q�A�̠�QJ�'���;��P�wp��S��Z
׽{��u����b�`��@�N��^�qF�x.f���u�h��|��a;;�9�,X�э�X�����cu����}�=�lN9����>S0yԘ�G�nv�w2�(t� �)�{Z$���W�m�6�W����D���Lnw�uh��c (��G]@'�o��u^Z�0Q2P'���T6��]vc/Q��EF���{mc�m��ڪ6�A_6܌�P� �2�q����A�#Nd��5��k�~W��n��0�ճ�*<1�bzy=2�:_$�ˀv�CV�xK�s�Y�K|AN�ԭb-b�NB�6����6��"�/T>'a�I�8
��#&K�A���)���	}N���������$�"R��QEDj:}�_z������dQ�4�_��Ҁ@�F�b�_��2q�E�eM�}`[5�ȷ�	�]�����zR��2s*Up�}2Pj�u_�D^���!T=~o�7�'hDC�p��5?=���|*���r�����J3�K �ZB�����(��Ӧ\;�#��qhS��?cĒm��Y�Sp��WD�qJ`�~<
��B$�'��AC²G���������;jk?GÀfvtTw; ;	��t��;-qV�U�.mj�//����x��)��jy<�{�]��JrП��$
��Uq-�5�g/1�I!"�A���D`$l�Jr���O��%��>&d�f�n������G$��G=^�x���k��:�`�)`hsD>"{f�����k�T4^�d����ў�uFj�}��:��d*kr������&���y�����܉u�\lC��I�S�����u��ʸ�w�kЫ��k�{�0h�.��6�M����3��l�����T���WW���}�-�߾ԧ���<�Pk����0~M�%Lr�vk[`%�H��^��g�ŀS�%�Č�g5���|5q����>�4q�q��36���YE��.pS�ɫDZU(�,e�7!A������K�h(�k���˼�'��O�gʃXF����������PU�����aw�-�2��d4K�1�.�?_HR�L~�U���r�����zu1�69�b��5z`HW��2ٲ�ȸ$�X���W��])q�w�'5�c�'C�`I��H�'�h9zT-+��=�{�
�O�1�|VH�2f�0�������T	C=���AѹV[&�C��-r>��̋�1�<�zIw�q#t�e�Y��)J4]��.���~�B��]B��q��{$�[��r�A|yF"����z��:�����vj�)�|���
�S�&�����Ay���Zի[g��
jI 1뻙��ڦ8Z�qd�(��<` ��E`�7��ի([!7l��:���9P(��)"��	vwE/�`o-��E����k�)���l��?��i3%�:�VP�x3ƭz"�AM�����[W�QN�?Q̐��F^��?;��|�xE�d�<��r��4b���搚#��ӿ��*��@����[��E�~��&\�̎nX��L��}��)��_����q�ߔ����4�Q-0�	H	8R�.��L )[��\��� �@g�Rj�D��l�6�,��������%ޡ3g$(<S�֣S�jZ�.]L�#n��	�}�$
�����M�z�w��>�����+����@+����������~��� �Ռɉ���M�qT�Ϲ�Z�K�e���x�݀�K��'���j��܈��4P�-�>%s�8�.t����jXv��=e�=f�F��u�L���y�jS��Yk�Z^��$���d z��P���d�����?3����Gz���,�x;�H��K��Sf`��٤B ] uL���Z���d%�K^��7�ԲJ�2�8���\�^�b�.1�7� �������PR㨘5)�M��5c��� 8�^͇|����KK�$�7���O|��t����a�,&b]� �L�&��o��:%�>�`71� @�2��ш����z�M��e6_0���{<
£�=��y�S��٫WF�4�C{"�{�����wg�@d\�k� ��h���"��G� ���x��T'�@�(&��S�õe���d7msu��� �b�z�K��mX�W@�l����h>��MR� ��'�.ٓ����p�Ηh�:亐 iB�P@f��*��sD(�%*�i�okO:]����:-�o:�i1�A���?���Z�]j��ŋ9�+%�0&�u{�y?�;�|w�ޕ��u%��#�g����ɍ/A���_�(�vh)�.E�.�r4M��Ҕ�vT',�P��Hߘ �Q�"�&NM,�ib�&kl���Z�r�N��)�������2��q3b�U���V�`ʏfn5.xRM��D�R�΂���o��6�n�;��r�( ���n�?�U,�����0x3��V�"�g��3��e})c���k��X�6�w��2"�)2�*\�l���F��^��׮/�3��HG�6�����u�dK9�wّS%;E;�h�-BRb��ѫ�	�gk��d��"�57	���#�����mz����X��#k�:y��T����GZL%˯�t4b��>� ��ɠg�\!e���k�.��g��7���v/�T>D�<%r�b���Q�\�O���,6���#��`��o�i���a�R�e`�UǽuRz�}%z�w<:��7��=C�F�z�G�xw�ԫl��
�"�*A��w��]|���Eat�O���?|*��	�)���
���[��ga�C�9n��y&zNT![�]�F:�@'׌t�V�7�}�0W ��+驉��<��N�
cQ��>-�:��hd�f�Z������0��Җ�)|g�K~���ld�g���.�]A���2U7���ߝ)��8��_�>�@��9Hfk���j+DV�����\P��N�_������m�c�ns��dd��$I^����CL<�+�f�Ǿ{.oB�2�db��R_C�����ʲ�e�`���\�����ix�[�6��[q��)�K\�
*�O��HV�W� 2�؞I ���]{�{]�~�Gbc�y��ؖ$��_7T��}��{�t�o�6���)pL�|��<4�re��4�u�@����三p�uM�8n�u�b�-�7b��0����S���c檖M�А��B.���<Jp1����:�1�ؾ�P���Ǔ�:F��~�N��Ք1��/��>v���l�]��7i،�,]`M���lǊ6{�.�L�� (���0ܥ.;��':�NLc@G	���5����w�X>�u�e�s�#�R�{$��!�יGs�o��#������]st�Je�����mO�b�U�_3�� t2\>�,��c�VXl�/�Rႃ4
9wI ��3���AЁS�#fJ\q,�bN@f��y�'�l9L�A����v���`���B�&�����J\�]!����4?r�>"�=/8��a���!��M��PR���Υ�F$py�<0�\D�aY/N�f������`5�P��-�"r��^�0H[���.��=ޛ���PX;Q)-x��)���I�^������0f<cz�O�g�����he��^���D��dP��-ח�[��O��l���Ī�q�闇�-��R��_vR�6��v��mk������b	E����Du���wf�n~��~ћ�2�ޥ�]��&��R�Yd~��#��e�R+�g+�0��(�his&]XU����@�.����3Zj�6h�#����S'I�	���`~g��>��,�g��h��6����:�ԧ̺�_d3u�kC){.��Ff�+�F|yk<4A2���<�O� �������S8�VZ=S�,!��YZp��%��SG���G敛(V����g�m|��g�:����f��"b7�G3��i���l�I�'?�`5'��im��oݑ�%b{]�7#������[0��C��G�O�	���c�}�S���G��Nz.@������'n>��e� K�e2���p��̺�W�y#��w�9� 
�L1�,�|H��o�z����89&��	'���1|�rއ�v3�Sx'�m ��$���E��I���Z¢/nm�9J!��vp�KϠ���P�Z�n�y*L��\d SX�7} :��f2?��$��
K��|�'�do7;ۿ2ܠ�2ʪZ��?x��
D�p����Ղ�H6H�]��݊�7�f{��Z�V��n�}{�/�rk��Y\�� �hq?��,3��� ���.6:;��1qӄH4O���_k2�!L$�#����:���ԛ��Z�Zy�M6.��d���pߜ�" ޭ��6�;d)��Jum>䬆ޱgG�����M�\�D4���׫p����f���ք��U}	=8�brN3XR�X����C��XN��\��ɫ���Cc]����`@�����'���+���A73wƢ���/�FX��12�6�X/3���tW*� u*����V�4y��}-XEV�tC���/vy��t��St��
i���P�pom��R����$�R�c`��t'������J��A�K����Pܺ^����}
�g&E��*(�0��X=��d�wJ��h�ŀ?bK�S��]�+��!�lh�E���g�~�~c���#֪\����U^>\������.�O.w��I�BCT���N��R0�[�jl�B�+H��.7/���>ɪ���{��4�g=|���S��0(�\9H�?�1��3~�N��B��~��܊U��������_�U��x"9�Ӕ�%M�S�w@w����k�tӶ��
1�^�g��O�#�ׂJVx�>�Iy���T[����v"a�_�t�-�)�ol�P�V��%ZZ~���"��{�J����1������C����d��l FfX0�J6�7\�.������`1?P>K���@F�r���@B*f�$�nR�&�1�s���幇��V���?������k$�͊N�>�{�!��G
��([���dv�v�en9��듊i^���
���T��por�sW�6e�6������?A���/u�u:�X�
&�q�:�9�0�'�,"q���2A>��M��(�����͙�{!7k�gy�_[�F0 �
o���"Sּ��Z�ơ���d`h��3E�*ꔋ�G&6 Kk��e�k�m�YS��w�^�a��2m�,���u��gj�o��xn�s��+x�����<`���;k��C���ܙ��~͑Ѥ�%&��p-��Cgmݒ�����8.ҳ�ꭏ��f sS~'&E|�n�Wߴ�	vJs���Lg�3o7��H��p�^֋�\F������3� �k{ʁ�?i���ӃvǄ�.��DD�;^J��A�6%����3��d�� ��+'�H�a��t�~����D\3 o~`���43W�#Y_����Cmݚ=�r��ʀ��x�k���m���. �sY/�CE�}��|�����j��-���0��i2u�JF86ue�x��|�z����� ����q @C.U��-�y�����E|X�wjPe��!L�26X�&��KW�O�O�� u+�{���F�&Q=��b	�����	?���dڞ�����ॴ�C�������v�i�D�H�[`�Mq+��y@
�N��Y+�OF�F����h�,.�/��Lc�����?�{�G����B�-*��/�����	\�`���3Cj0ԩU��u��Y��.梜�d&еUT轀PeK�]���`��Ÿw� �<�BO7��i2�V����U�j(�/��E�Su����-|e#����շ٬j��A;J�E��貁���N}�#e�lm��(�ـ"�j(1I��O��>�B���v�&��)k��n�EhPTy�i=g�����X'5�	��p���۶;��Ҷ0���b����݂�q7�M��KB7�Wr��I�j�D;��`s�_�A�Uv9�eo*޹@�9n	�+�������W �Fx)��4����T���b�������wf�/�����&�G�k�^k�VF�i��E��.�8AH�.����b��D�<�j���P��0t����Z\��b��4+�jjy64�w��a�F��+ң����kx{TiH2o�[� �2p��mR6n��F/�R=�e�>:B7�!��=���wF�~�3K��q�mQ��a��+_��(-�*�����XZw��//�#1��(�@3�,~���E�Y�Y�����4�$�KQ��L|DfQ�́=FW�1�%����*�p�
�� ����{3���+��.O�,�C�$\�i�Gm��O���C�E^�l��)��>g��x�w��p.���1Q��?���$�q�rA�4N�y\�	�����SV���ޗ�z�[&-(���A,wfwS��P���ɟL���a���h�S*}x�Dģ��_�!R+<0QGM����Qk	S��.��Ϛ0�W����By��ʭW��u�ƶ��>A�2����i_���� ?�f�(��������U��K�x�����������o:��N���e&H���2X���|��]���WY��#
R�5��˩����C�TqAL}EL���㰴���%�D�����~Z��G�0���B�it�����`g��Z; P6c����+�,�QЩ&c���!�2(;P'hoZ���B����	&��{�({Jdүȓ�w����Ҁ��9�����x��zU^�m^+�['Fs�{H4C����l���Us��T� *B���{�^vB5�ܴy)�?|WB�U�[��ۀ�����8�,+�G<x��d�k`z➲+m<p2>��jp�Qe�V�ػ#f4}���?&8P���!�ڠUG�L�9�OcQ�΅�� T��/2�p+Q�R����L���E���)^����뽸|}�Aøb�	�g���e=��K����n�ė�������"���.���
f��S�x�s��=.�(�*T�P��F�q'�	��Ӷ�l=tt3�R7uY�=^��UO��v��V-��e���$�9�H�i�X���C�Ҟ�����+t�z�cͣ�{����h��Y�3����QA�4�o+�>X��m�!¶v6M)�j���}[�tP
� \������{�_�n_�[�]Î_�SБ392נQg}�Ν�ER�͏�{٬{b�>4B�x��X�=P�'�2�� ���Q%�p���C�~ӵl�\��eyY�y��|� f����x�_��S8#�Xҏ&c'�t���r~|����Bw��Γ3Cl7�}5Y����[��S����CH��B�t���X�=�H]��>�hv7N<�)�jH���y��A�hÌ�$��G������Jj`��w�tL���KD��-�by���?	�	Z�r���O |A{�uW|���(�E�z�Q�i���)�\4HTVMe������`UP&#ވ��f���,���p��#�*�$0�A,a���,���%�P�T6#�E/<��Wy�tq��%-���4v|9H��vS/7G$g��R+�?��C���8�|��0)ݰ�fi}x�&����r
�E2lJ�~�� Z�b����^�����XC�L��v3�rf]����19��?��w����-L�V ��b6�Q�����'�*YQY5e��������F����"n�
uz�t�,������D暤�/02qo�| �����f�,�ڸM��.T�Q(�	��_�LE0�y�.c*� h*:�Yi:	G2�`1e�;t�������6ڽj��Ҷ,ʑ1�+�RB�nվ~�~j�.�0޺����y�y�=ze�}�x8-A�Y�l�y��6zw�G�CK����C�h���P%!HXu;p/u$���;]��Z@W��A���+�35؍�#�Ȅh�����D&�٥�X��W���ʈY�GNoy��<�d`��Q��f5&�aj#m�0�����4�G�s����HB�d���3���Lǽ�&�T���=���S�yB�К�܄�eI9fB��'�P��3�.�`)<�j�~���è�;����C��;�G�7��a���D�lM���p��:4X��0�F7ة���?�k��W��e�ϻ�ASSi����S�eb��b���M�[O��f��Ug�YM��l�@�$��[v7:g��%x���37���c�:aC��bfL�otW[C��W>��__����Sș� �J�4{�_�v��͞�������VR�������!��8V]]
Z>/-H�Mma���s�N�������ݛ��xE���W��v�f�t�i�9M�ȗ��)O��4�Wl�w��t�Fn��Od^���А֢�x:���K�i�cG��0n��9����tL���U)߷�f�^��9�k����϶�N��¼��N0.��Ʒ����P�]/8���֝:�t�[�3���mw,xg<7�އ���D͝���Q>��]R�8�����%U�u�j�k�{�W'o�y�U[��.��Ŋ�SNg����_�ӳ����im�w���L�b`�z0���Z�&eB_�6�i��xI�ՂM��ǯ:Ru���.-I��N�Ŏ���Ҫ��R��.Û�E�����{��M�x�5���w)�@�D����+���ZuV�鶛�;g'}FpNV��sfy���X`��Z��k/�:4�?�8�{��S0���f��N�D��X
0q)���w]��8��g2Mi
U��g��2J]X��;��oK��x3����ܼ�U��?��,�bX��<�b�(%���!���Z`�:��tݛ7�0��#��ٰ�{]��D��j�_
��)u�m���	��O# h�n�����8�k*�ΪF{Șמ�AdY��I6��?
E�ࠪ��l�d1s_���#LiW��K���L���㕏�]��q��'z8p��G�U�̵�>#�+>�9:��Wy�ݼ̨�4L��}MA�tDp������:*_i��it�:�06��m,�[�����z��d���LZ����[�gS��Ώ<��D��ub�w�Y��*�\�:��^�MRR�ⓛ�5�b�8fa��tHy
5x
�ݓ����=LB��BT��=������س�o�i�Ie�8��ٟ\Tqv��:$����#�ڃ���F�
~'uz�Z�q��S�sdG�]���y$�JE�$��������"fL#`,�L�J��]�C�ds�TP��9�#�)tzbpmR{�@��[������7�=~�⎅nQ@��ͱ3
��Uג����:ь���z#m"we)��fr��kҾn�O���U!D�r�u5Y0o�#��	k��2�4y����ͤ8 A�EF�z#�֋~�8Dψ9u����q8����VHջ9��O9�\?�q��F��L��<r�%�_�������3}X�k��o��T�@�r�������������<U�����Yq�άڈ����CwsFS���x���~.�n�s���?�Bp��xP��W0�7t�O�|�� �H7��?F����%�IK��IR�#@�V4/H%�oqp���x��,���a���]ΌH�$�21�+0��+�^ �Z�Z'�޶͸�1�7�u���"�p��8B(���g��J��c[�E��':�3�	�qz�ĎpS��~�V�*�b�r�d�r��s�܍LU���/^��A>��r�O1��������t�1cv"5ǂVu��s(t� /	��[�,�X6��M;��`5�{�ɬl/N�94w>�1�6G�XA�gهy�Y{?�(��p��^�.�B����l���$��0�"0�������G�-��P���DwӾ�h8�����P1f*>kn+k������ufOvD<�$;񈕯Ե�C:oE(CAZ��d�"�>��Ϲ\�O�I�@2��F2;)߮��(F�Ak">i�ŁjR���&���p�-�=V�C֡.q�R,16eG�M>���Y�?�2��Y�;޹��'*<u޿�-R8-
X�m�����|`�%!���&5ҡ`�T��ՠ������P}�{�&!��rb��6����~@�Xw6�]���<����������=�ɓp�Lg}��>Qd�o���t�%!�� OЏ:��|oc�0�����d_ԡ�������M�n�.�\:�O}��֡X\�(��g(z�(��d&�4uf���)҉o�UA��J*xM?�8�B(R��^�S��#@]]�zm�D���<���G離Ϳ�+ۑ�W���4���`;g�37����c��7M��\�\]BM�eKXhlk�&򵌛�V���E�)u�2��ς���u��`QN��E`�,y����/p;\ru�� �Pz�b��Dj��0pI���#�M��9C;�}��=;�p��EO�P�l�w��6X��L'�+���@������7	mx�M��ƚ����8��y�:��I4<JXȰ�!� � �U�����h�i���GT��S�p�8f.�/ER��b�l&�^���������aL	�{�c��2�,�RS������GR$�xT	b�3C�8&P�(��Eu�ca� ���;guDEW��q�{܎������?-oS���#��H���E�k�W��J�����^��OԯP�n)W]�u5�%o�v�SW"�a��#����"��G+��k�q'/�F���Nz�K��]o��U
�<M �lB�$��)jn:��]�T�X���J��kSB����B�(������$���7����/<�2q:c�D��_xH;�	@y��U�h2~4�5�ՆJj��'oSO_!�	V�M�7?AC�1G���;�!�L�bo�4�/!�D�Oi��|0�tzZbB$���|�RE��5e���9n�/A�3y��X��wYI�(�Og�f��N�N�#m��6c�GD%uR�~����R�����H���r�:����x#.���+9���-���_ lMY�Y�S��C�S�ɉ��!�"�}�^]�����^�q���`-r�K�}ۈ�@��X?�.�p1�R"��2��k��XZ�˽�D�Օ,Ai������zR���w�<T^�c*����p�m�,�+�Ԃ�{�+��]�"|,R�{�t�9�x�RV�p��TwB�x�8�d���;����T�ஊ�����^`@~� q6^0�*��V<��1�U*u��ɕ~I�5%,��;&��ѹ�ژ+�����G�q;(<%^q��@���_�$}�i���:+<�Z3¢p�W�tt�Z���Ts�� #/�~ɰѵl��b9|��噐�;k� �pc����|y�?�Q��֬�"'SD��e��
(r�3�dtO]T����܀ϔ{2�S���j I|��7���in �ԡ�W���zt�M�aQ���Er��4��`F�D���O��2;��*�>wNg�� Ed�M�j�
�����D���,N�������+Y��	Jz���Ϙ
�3۶њ�*F�+R���A�4F��ˇ&<�nUX��a����=�F�N-<����89�G��f���P�8�%U���-����Բ�<Fڛtz![ND_��V?�wksJ��k����P4~&�}�'(�;gr�(�O���ԗ�޴"v�_s>�/J=�n���%�d����'YF�Lj(U�|9��8_��bE���x�R��^�D�(6v�.�85�\.�w/�)�:+A;����d��aLЭr�˗݂&ճ�mmb��9�nv��H\;�G
�Q�J�A�f)~�l�/Λ���]s�G�þ��������5�K��Go�ԃ�$�ľ鶛�9�C��ubc�3�t�6s�@i��,�����(�G�pd�zUnӦ����Ӗa%zQr�T�Y�E�0�e~�{�nll�QI���E��r����z����s���lR&Rnb�Y��*��`@��x����ͷN��l�M¢�xEh# ���^E�	�#1�[`�7�syIe/���X�¿.�CK�F�L ��\@.�b�xJs��M�=b��b��8��S
+AR��(K��=-r[��n��*��=R�=U�ː:A֬��1;-����0�f�u��K����V��3�َ.ͽ���>�*���2)�=(T�ǋ��$�₍�4�"�M��9J��@q.�t73/ɝ�*|h���s��7@7�Z��p"�qrd�6(�c�[����A*?��z��k�!`�������Ț�.���|���y{p��1[79��ybȲ11U:��b�����ς����k�5)�������F ͞C�_r�o3�Ĳ*md'H	�w��7VV�yZr(�K�u�؋$!@���Z���i)�*�(�.�8D�&I�]��<W}�n?�%�ّIo{���Oy�FE���3C�.�� 1�.�y�f8���P�>렐V<����{+�� �X8Τ$L,�fj1'U����o��M����_}?�e�e��b���p4^��������@||�|^�2`>�FjÊV7����DQ6$_T=�vM9@J�%��0��!�Ґ�GD2͆�CM���>M�`K���Y�*U� ���S���[���k�!P^�j���������*���`l�~��~(5��#�S/bf�{t䗏(�	�c/ײP��9�zRV1����_�2XYֺP�'��*��d&�l����' 7�6^���y�^�{���Z�c�tR�D�A5���[����d+V��i�_v�H9�oi�=R)�M7rL'x�o_!�+A��Vm0e;_��$=�s&�\,��@�P��9��I�Σ3��p�+I��Cq�aw�K	��	bRF#�w1�t�;���Qi�����`X��zdhg(%&~>/����5ۀ%�mߧ�XO��X7)��x���ǯ����Yڽ���>�P����8(T�dT�sVh�2���\!���2�.��&�ySW�He-I�W+1ddx��K��k��B��RMɩC+\��TؒXƊ�D�'���uԂ�Y�aJ�}�����.�Ę��d�?Ux�Z
y��m���<s~���!r�ǀޒ����H��y4�W� tv����k ��܉����������]jG���J�"�ep��#D�.����)r?��
foc���E	�e-4s����0Zƚ,��R&�!��O���uN�o�<��$O+���؃�~�|{'{��2��3�������~>�[s݄2|�����NjቝחG/�~�#�BEbn|*3wB�&Xʔ�8�Fn��
���3d��|H��d��q��M���3���ڥ�����|���v���:M�tn�������p����WH�g�7a�Puv=Mm�Uc��q2�vUc>���X�����H��	��U��y�q�۫�'�Wy�����_�Qց�/L�=�HV2�+�s����zyq��ENMtp*XX�U	ϷE�����)m�4p��P�&p�e]�yԢ\֥p���.���9vXƄ0G��0&������1k:R��qC��덢3,|����zO�
�Dj�:� ����1���?���E7���~���<�/��*24�4Uv��"y���3"��n�ORR��0N�sC%!�fTmAø�;5��Zr����K���_���Q5���&d�58!��������ҳ�J�� 4�VF������ӱ��s7��34Ӂ&f�y�pK���	�V=L��2�	F����9_L�F#���IC��ؗ�?u�Q�/Pa��:f�@tnvD�8*q�8��4�R��6��B���*�4��)��(�&��;Qc,	�Y��S�saS"[���o��)��sM���}O�� �s����w΁ �֏�/7Q߃/�M#:S�A_�3��Q��
@���b�p��e���v.�$���I�/]Q+C�>���>��I��*�������$<a�r�;IӣsKC|���.���lX�ߏ�ϧY��n�k^i*�I/
52'����R�r�6l����.�vn.=�b�E�g�ukn�B��-L��y��YRn��sT�V٫���W:��%�޻E���y����4�Rv�2���i\I�nd+u���]Vpo{)�H&W�
`F�ϋ3�g~W��.zu��<��X����aK�!l��߁Q�5��j Tۍ �Đ�B\�2~MM|g�,I�Pv[1��aI#`0��K`���m��@L�2OQ�j�ꢔn�U^�6`�޲|Z��u'F����H� ��C������
���"�e�*�Y�f�r��� �U����=��YQٕk�%�{�J�_$��MG׮-�l}$�<1��s�P+��j���N�[ ��,���r!l�J�&��V	{��2I�Q��sb޾a3R��əS��t�3L��o�
��)�����ݹX��hP��J��߫G`��,OSX��#@�=� ���\�i�`��`B򓔲ϫmI&�i����u����o&�fa�d�!~(E����@�1�?��3V�����=����TZ���?(�#������=5��{2��G�H ˑ<�ɸW�����ƾ�A.��R �pƩ���nR�kn<a ��iҸ���M�dz6%�i}Y����>��j���հ��D�rP�Dx�@�v4N.�������h�7z{��Y>���-�ބ��=p+���/�5����B�_�ٯ-�j�D��*�B�k&�3��`�cj-x�=BV�;P�~�Z~�b�Ă�3'��$C��pL��6.�-T��j�eu�M���P�U>���μ���bh�w�-㸆?Fp@F��P�N�/�w:<�b�Ϝ;�U���Ϥ�K3�c��(�9������L�� ��ƪ�yCs$�Ԑ�����<`3S���T)�ocz67�T����,�vP.�i���ذـ�!K����-a��#� ����o�ϓ����vϾ5�g�y����=�1�6�+#v6dtcG�z[����(
�L���I���/Hw O7��p��fx��=�
"#^w�F:8w͋�x�(�`�����;k43�J$)����R��&�����E��U�Z4��a|	�u�n�y=��m OV�bOD�.Q���U W���!��",t�aL(�t����6%�x����68�dE$)��6T|���tJa�'��+����=8�
��_��ӷG"D����]��G�`��z&�h0T�@{t��~ײ�ã���h{�"Za������1P5e��7�"� :-������^^��ks��*ڬ#����8]"��������s�a�O��쩸� ��NоJC%\<��*��d�÷U����:D���#�̄�!��2��<���q>E�Fb��R$�Uo�'����$�f�6�f��U|��{W����J/4Ɨ��NE��Нt���'EN)�I>��,��u��E�g�N�}�Y�f%�*�i�Hӓ���[<��%x!�B�p�V��<�F�r�y�;�2���  n�X.�[��ݖ��m^��{��냕 4j�`]&<�!�3�ͳj
�dŊJ��u�~Lap�e�<���k�%уeq�7��#I8�j�]�F
u�牲�%_�M7�bl�c4.6��a�Az%�\n8�KB����m��fY�e���@�p��q�Z�W �m���-
����f��pn_����`��2�Պ�H��0�������2d͙�be��{��⢬�;�X��V�e�+RK�eaˏ�?�/�\�βa�|���T��>q.�����bP���?�����ؓ��s 8vl�<7,G�w7�
S�C�Ie_]/�,OÚ�h �����a�W�֭����;��V���cl�5#*��;�R/�Q��<_��i�t���Zq��Qj>)	���~��P����dBH��c�܂�c�,RK,��l��m����w�]��,As#Mh�J#8"�rO��iDON�����W��v�jQ�ܖ
��l��O�L���	|��C"�7�=M�T�N/�%o����������Z������ɽ�a&�F;���(��5�U�j� <Rr����9� ��T�'U�/ z����\|�O;�nQ��#X����u�x`�	)���,����$^��Z�)����[��H-���]~��Ym�yo.�`�.�aBEcO�&��q�v��z���z