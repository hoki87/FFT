��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ�����������"
"��[Mp� i��tOT���L�5�� ��{q6ab2�Mb��秒5���_�D��>M
3P2�My���[N}�j�����Q�n�g<ߡ?� �]�'�:�#��ܜ�kU�dI��:ZF*Ynd:�-4��s9\�&� ����݄�v������=!��7�0Y�z;LT0PKJt�j��ܓhu�\�0�^J������K��	�&��Žm��>(Rd�_,"������D�X���mK�#~@k$$z;�!S�M�ܑ��WQꥻu�	�,���Z����ߨ�A䷶ 8��a*s���>�<�T�78d���;յ��u�7�	����p?�:E�����i�C`)�M(.�u�T�/D�V�D�7��z�8������Ṷ��Q�!�������՚��#��,:�s�<%d��u�;��:	d���Pw��p�V�q�i%�)���F�@���<`a��ױ��)RO��i�R�;��c����a�:��h�����G�ZPE�w��T�i�m��'��g�M�T�늱_�h�������� 8O	������=�!���܏� �]���鞎���ET�@g�hQ9��M�Q�Q}�k��K�[\z�[�0���H����^���4Obv�0Wf��f �\�-�b��n�E�t�}Vl��ʜ:�ޮ���[���:�ڻ��>.|�����G,Q22)��Q��b�c]���MۡXo���t^č�"��R�؏�)��
p��v\�0RJ�2��|P����!�§�kG��$�;a����[������M(�ί����h�A5sh� g���TR��Ӟ7h@י|�Q(�^�~���o(����,�MƀW��fϴw||O`� ]��\x��/��oB�v�^v�^�W%�� �a[2'A!͘2?`��`-��
���c��(W-��V���b�\�{����a���1��` a�7��ⰽ�]Zd�h�K
��~${�w�+r74@��x��@���7�4��R�x�l;�{�{��bqE>�н�L��Sq,¡5�Ч�Fo�}%,�-�af��0��c�ҵW��F+f���fo#E���G���ߤz�R���k,�������������C���fN��ݻ�u�4?��k�i<쪄�v��+���F�N��¨N�Y��ä�(%�Z�q�[�H��̿8=؋���������Y���[��G����ƊxP+Nc�:�1�#�%f�l��K��H�u�ȇd	�A��N恡�A\�7��G��^�?A4�'$��Òċ*�Qmu���_�K�ƞԒR.�؛|� R1�R�M�I����>�i�wX�-�Q\�A�7���D�g`�`�sJT0}�����SI�%�4"I)���S(>���T��S�_=a9����y�ZGϧ�Ƽ��y��?~%n��T���
H�bn0"�l/���oj�@�_@��M��f�>��d��,���	����]8 I	Ҭ��a���S���/� +(�j=Qv�"�Ÿ���n���2=F�9ch��U��ea�� 1:�ʯ�6Y:ק�ƘB��=�f��������s�N!�V�b����fr�ɳe��Z�璜���S�H���̹�.v�r�����ިLR+��\��P{��B,��E�5�:��ﻖ������g��T ����],�<1��e�h�Z��qR��ⴻO�u�_��q���m��b��DQ�m&������a�z�XW���e�1��47WG5�[��u���V�2k�%8?��i�t�� ����xԯ��&��]��Wݚ��VP2sr+!r
s2����%A� ̋��D������:�������H:����>�y�c�^,�2җl�7
U�W�>C�"��#��zQe���:_d8�'k�ڶ;ޏ��w�䫵���/�!m���F�J�8%WW*e����[ܐ_��!EM��L����S��I�S�o\���lڶ�@�����^#u"<?�qflz��HnX�������$*�D[�k���;��x����^5n��jO���H�{���5���t�ӵT���;�����#����>�)!�Ŀ��� ��J��0[�z+��rǵ�{0���a�<�mO���3����?�oS0]%.vn��[�qMXWL���5�840�؊��8+ƁR�Kf��~��0�=A�����~���mg��G�~��B�
�F�Gg9��e�җ9�@=K/�&<�X��+\/���U��hG�t�8>�	MC>��.ȵ��3�� �F���W�Ӱ�Oږv���������~e�|�������}+i���� ��/�8�㦇�<;�O������6���������lV�@��=�JCHu��dXn�"q�ܩZny��i�Os�T��g�#�D_�^8��b��3~`�N���w�F��@�#��y�s�f�=R\,~r�r���|�g4���4*oāL�ƨ�m�j
����I�,�O������?�]�ZoW����;�����G�kز҈j�S<�J�<�A}�l�S:ƨ�トQ�$Et�ſ���'���I����tDa���x��;K4���Ͳ�����m�4S�E����-��.nC�#�����w^*-���-}�ϙܟ.�ǂ����i��v1lI�8��M��҂�e�jA�4N���s��-��ۉF��]�¤�ZlGr]��MO��C�	
���F�g��E,CE����<P|��d��ՇX8�.S��5*��:��i�:��>m,����]���1�w�)�\]�� ]Z�!���!bw%��{�7o��g�\��o&- $�S�6�1������k��Ս�)<��[�.���$�HJ|�󡥛=HK&&Q~ ���q���J��#�4l�cg�A�=?����UGG���� }l�\����(��yM��u�BM{���.ST�	�D(�H�W����VA�
����
�'v0el;ۺ9SyRs�ιۤSM���'ׇ{�E�`}ӵ�)��%�]���
�v��[�P�_$d�}�Ȍ�U���z�>� �
n�e��� �2���ٝǤ�Ff��V}w�M��RG8��Y�b^f���@�ߧ�Zvb@H�[4d�VD3 sK&���� ǥ�X�-&&�M�ֿh�2��l%N�s"}�P�G�<Y�34,�h5����L���h�lp�]�r�d�C�(��p�J�`߬ќ����`3t���[i�KuPIҀ�1��Qz҂��+;�A.ť ���ݮ�T�۬�{]�`4�S�F��A����#�o���EU_���-��^�:!+��U��0��g�и��p`<��5fc:JD���
�Iݥx�x��@R��#(@/����LY-4��*shq+sy������N1����Fa��e��4i��!3!�����8��o��\m�AcY7pf�s������LS��ʃ??�Л24G�\�H�ﵑ���� p�����;����r��v^[��'����	N�?��L*��7
s�5�3.&��	�J�1,^��عNG��D��Cy�,�&��r��8+�Ў�e� 3Z�p���Bs�Ok	TO�������G�p���Xg�����#�-,�xl�2J�E\�sdh9�6+A��^�IǓf����=��R��o�g�=ڬnO՟v<�BhU��Q���J{!)먃�b�-�2T��^^Rq' !��Vg��߳_#»j��׸�l"zC0e���0�-�r[�I�i�'��`!Z�r�](��S�PV/Â�JM.�	�91���55���h{���F��S]��5�/��3�Y1�+2�(��ye9������1r/��Q2c�j���;ۀ����0�Yg�xB�<���6&R
�pA���?k�T�$�2��`��<��sPyf��% �l�"W�{g�����x�I�>��,��Qn��Ҽ1�#ݜ0��p8&� �^�6���xO�r��ې��m��?��CY��3a.�Q��\d)�h[�QAv�:�Yo��f�6rn�vע��]̕���L��2G��*u�g� O���t��L�s`��f����}\�c߃��$�&�B"�W�m��bw���Y#q~'D�&�$�
�>D�� 6�:~��x�Et'dy�eRrb��N;D�!�OxK���n��l�/��Ȟ`�Vn�z��Q�e��A$7_�*���s͚��|Vd��*p�h�^���K�Yz�:�m9���ݞ���������Ջ"���6%5*E1s�����=߽��'��sn���&�bt�7������C��L�@��F%��Ye/n�`$ ��_��"av���&>Ã��hL6�|�c�7ިn�*�ְ�yX�ܐ�/����1p�I�*�Ȥ��:���?��q4����������O)�q��4ow+?ِa+�4T��s�s�3��!^��TId��;CV8�ȖN��"��U�C_<~LhF��2� �iO�r1����X\���
u�giC:��o.�K�Y@*��O6�!0+n�)ȋ�N{x~iЩ\*B�PΟ�ƾ.k��X�ZL�㘂p�8�ڋ����3x������f�7�] ^fw��='�ƚ���V�>B��^��I��0�ً�7�/���Pݯ!�N���ή��`��0f�����'RQ<^�r+�����m��lO�u]�tph��Ko#�K�d�Ɍ�c�cT&�Hơ`�ѡ�ҋ,�s�_?��k@♘W��f7B���Ъn1���U�P���M�^��{q�v��\x�*1_#�|��g�ӪH&@�&+�ث��'2'O�+�Y���o��W��� Hױ=L	��4-}�d�P�z;���L,Nu��������q�BF���Z83��P�u,�� Q�d�"U�-�ź32l6�:�)�M��ǽ*(V�_G���w��V�`d�J��Xs��R�U�Gp��e�^��]Ȇ.�;$�bG�^�Bn���<���a�q��q����lZ)�#�d�#v���r�����J�(U�k
�J�D:�u��R޻H���"-�*TVH���Q.� ��3��ٖ[Lk[��[��}SMF�yFXIrڗ��P~�H��\y�Kr7�["��t��-O���&���*��Ң��ڝq��w�%g �%C�_�h]ȟ�z�T(����P�F/
0����옢��Q�*�;�~i�z4zAh�ں�<�d�Fom�(�+�C�L��o،2Hu���H�5c���1L�Q���V{Kx�N�f�F n�����ɭv���|��~�I;��z	�C���h�!�9��v�#�P�~?d.A|�IdbW@e齗(�r�[-���:~�F��A���_����o��X�h��[��j6�#`8��fi�el�BD�4Й�T,6+3�9�^8��R�����-�颺�\�f
h�
�݅#+��4�
�O����Q{��7FԳl~(9��ӘR�.�US�eE���7( ۺƲ �S��Q%Q�g�s$^�t�ڳi3�]��~����-ޥ�����A--�����lYw�҉ж%���0�>���.�8��#��87�A\>��f�P��A�ȴ��ǆb�V^ڠw��=Lp|[S���cd$|����5x7�y#U�hL������ ��%�ɒ�	;A�xc��'ϕ�A�F��ܓ6����{�Xo�h����Ȃ��=�i^���N�]��fs�ҕ�>��J[��1����!|G���f�b�L�25���HA��szW��S���XTa�h�<������C�
R�QgAd�k`Q�q�$	�U߷�d֐4�|�󦧲�ADg$�2\_�?k+1�"��)���^U��3��:+��I�O����G����B�W�}qN|G*&"ߏE����r�a?��Jq}c!�KR��9��U.����6(y���i��z~���P$�� V��FBh�� ?�|(KG*g�&>��z�/8*q�\��7�Eej��S�#ҺJ��k�Q��]V*��D�QmӜ*����l����J��)�)Kp������Q�D�_��b�`;�9�)Ô�J뇎���_�밧dj��A�Q�\�(A}o~��s� ƨDR�~�۰G����� +��@9�$�sޝ}���#��+���S�+��+HFm7�K��&�ְ�ҵ�%���l��k�n�v�)-���()�Zf�H�����68�d��_9b�Q��.�x����
�n�A����-�Ҋ�ُ�>ҹ�{�3C�穸`Ѿ�T��RsH�L�	��G�q�@������!�c�`��`�������]W�0�����y�x��GVIgkmg*�偅���ܮ���9-IP|s��5u�V�C���@p��8|�HM��å��C��`�j,��HF���W�_j�:�:����7jwO.�joo	]�Z�4F��8�e��1���`�3�j3c|3��~`^�����o�����[ DB���EM���҄x��d���I��ȬTFق �MO4X
���o�c�����dP�˞2��<X�"��~\i��?R"�����NόZ��1�#(3����6	ۭVD\�C2��핻��ʣ�; i�}�8����,�#�!��V���Ӌ�G��b���Y,x���_�F�ӌ��@̞�S�5��8uG�r�k�/�:���= Z�q�mW��*ۈ�Bq?iK�]R�c��ŋ�c9��E����YC�faw�ӳ�A|�7-��?�15PFfIsHC��.�����x*Qv2�X�7~}#��T��0���6��f���U8kB�$�?�]�L*�nciWwg �Р�i맖��{�����l�fv.�6`�;{:zM~���|n=�Z^���D1��;	�\��dLMl�"5	gf�Sʛ�v��Es��S4l��Bqo�t��y���k��=��@�-@�34M�6�_�+Qdm`���BƮE-	����m ԓ�������my�������IU2km-�-gy��I�ޜ�J����Ox�ˊ��@m�7R!kd�R�wUU{Z��us��>�8����g���v�)7_���r]�l����m���S �'^K����riϧN5XK��w��п��;���ޔ�.�$��v������Sme���.\�	�a�uZ2�<��w�&s6�A�������0Q��ѻ%tzQ�W)��������&���,��z�=67)2bLFQ:w�㯽�^���$��rt�/ғ��l�����tx��mK�Z-��A�j\C��N|}Ӝ��_���O���	����/H��t�P<��#�Xv�JY�$��Vݍ姑 7���L��>�و�e�p�,\� ��Rf3�lI��yihVw��ub�J��IĠ�@�>��|2�i�P���l��a��oEb���a�n���´���s�$NP{3�^�(2OO��nx}�_��W�����|������_�5���˷r�ӊ$��Q���hJ�IE�snG��-5���y)��B����~�6r0�<W��Fq��i��؏�ggk��4�-�~ ��v���O_�=k�C7z�sJp��1_��%5R)[`��0�����r�z|�|��$��*#]X���9�2��^��,!i�}�_8��|Ɠ��!�hCb�:�o�G��~�@1�����@�,������_�Eү�C���'�)���R�pO���ʧ ]4�~�u�،vx��<Gs����;T87�)�2<��+A����!$�i���)H7�q��.��Ro���m߮��bFEn`A����Oy8Y���ǅ��7�:Y��v��G��qnr��X�}���49tv�9�8'g��hڸ���T+�=�w�����(����	�md��U
	��BϬB�{�P)�3�&�ԧYn���5x�0&�OKH	_�ZlvG֩�NB�3a7e���a�\@p�
���Q���:����uj����
��3���إ*\�vf