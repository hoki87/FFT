��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�#&��#�<����軥�JƆ���,����TL�����cߣH�ϫ�о�Vy��/B�h��I��|�I�%=$Q>ߝo�׬9O��7�ٶWf|�$��E7��x�AO�&BGFYHO\oe��V���ન���*����������8��u���e��fATy�Vh����k��B���=��L�U{���M�pϡ�� t��2�ef�M#ߞ�xW�"�H�`�>�;PL{����_-@����(T8�*�ԪA�©~a�q�!
q.�˲Gp*�s�1�Yd&�f��7vl���M�(���$�"Q���XyΓVG�t�D�xU��jH8|�5�<-BoKJ0�	cG~w�������xѩj�B�k��3�~�^F3��:z5l2���k��}�b����ʃNo(��3��:�����~Yz5���m�/���� ��%)Iai�U�SQ#Gq�^�����r��L��-`<���\s��x8�c,�|=�B�ve帰��x�~��#qNP����X���A���&w�� ��D0�k,v�:Le}I}����BP-��_�v���26�;KW��<?1�N�1��e�/_%�X-��/���p�%񆭊�'4+.zm$�)�s�����p��� ܭJb��JQ<o��33n�mAzyb.7z���������̨�f �<��������:��!�LW5�tv��,1�(�m�N�L�;c��)�^��Z��@윓e��:��z�ağ{Q�q 1��F7}Z�i������'+�-։��>	��q�/�3h�m}�C��Z�Y�-��m��Z��!o4�����������N7���4���G�k�l��l�`�a�f{:M��h���ނ:9�P��: ���+�S��W7��w�9|���zC�5>7z�,��\�k1���I��N��9�]{�:cЛã(ߵe��eH\���	|*���!�F1�h	�!�����`g,?��"aZ9��"|E3�Z�r�uf��3�N��MA�G�GL�{�{�D�@N���FP�V
X�$��t�[����rƎ�����h�7⑯(��f�k+�yr��3��p�;?��r��H����\[���r�YH����M%]�a�^U�� Ə�6<S�1�-a� ���:��)��Z��׼L�^Kο�������sI�W���َM�K�������H����B��z#��v+�6���ܭ�g�����0��U\����[�\�`V�Rh��|J�Q��x�œ~}�4�AΝ�>9��n�^�C�Th`����<�\�n	�TCp��w8~?ɫ�����]�0�3 �z�r�y5qb��cٖ�?�&j�Hk2ٻS�]�M+T������e����lѳ�n�Ί�e�:�ccF��k�`�ûMg�T�b ���Y����	y<a}��?|!��B>{������4�|/d��v~�D�z5	l�t�.f;��K�T����^��LD�j�?ut�O@3��뉹�Y�>�xN�,lZ��f�f�)��~��i�U�� �M��C|!3F�@��
h�B>$��AF�9$en�U�8{��<Uh�L}#TD�M6��o*Z?��ȋȕ�WY�ٮ(�֓}õ���*���2Բ�.��RO-��ƾϙ���ʹCRx�2��!v�<yp��w?���A�t�r��"�l� �3�sI\�Z~сƬ�O=��0B��>9r=��Y����7�ݴ�bM��ߛ�<��~q���G4��N�8�whU��|�|U#���D���߭;� �Aksh�uǉ]�Z^O|������C߮d~�2��
���yj���B�������OcEiɣ�A}r%�c �T�� vq^R��T���h�K�}�̆��8{��o&ѵ����k��aw9M���*�8Âr�S/1Ie�~���� �?�J��֘K�,��՘`Y�$�cʟY��Xқ��3������w�
�9ln�6��"�Zu�v�Z�^b�'��Un3֛U';-f!�o�O�8��+�.&c�(\h��p�����rn�!ƖkE��(r�:���Ge���U �#�,��$Ed����$���˯]v^hbC��2����-��[�*�Lq�"��rC�z�"����^C�v{K�<���^X�&�P���$`��]7|�)ts��s�o���լ~��Ǣ�Xa��L۽{�?�O�
���J�k�*��q�W)�����=��0r����up�͊�C/ _�Ӑ듆�"v	b�/v��� ��6������`g���}.�=���H3�����\�y�	)��Yh���0�F<K.���K;�)�si����Z-��ly(��D
�4��g*�WY%ʡ���]7Q�&�em��V�X֖ۅ� �T����CŊ�hTl_H���)D��
���aƶ��V��1�70%�̨�2R����h��>�yp�ӆ����߬

�F|F:HΨ�r��jJ'DC+?��A8F�������A!��o�h̶�?%&u��^!�
[�su�5Z��W�]>���*��sg���oQ��n��߇$ź�:�,	y��h�,n\\w���/Sf��o�N�Z�i��Ro�ꎱ$Ur� W��pB��g�5|i�xC,0�y�8�4�lt5�B!P����9���\-*�k��[->�Y�l:c���x�(^��f��ý�4���8LJ+�=�DDí;��L���*�#���2N�/<�E0���ؓ=�,�{ق������wbB��K)c�U��׆�=P1ŏ��/��?�8Fc�|B����?ׯVP���F$�>Y���צ"�����P���I��8�V{�/U�����)h�2g;�Td��c���U����J��П��d-�m�ó떥�}ʕn��	����^��m^�#�|�\O�M��<��B�	w��B��>z�	CT@��)��88K_G{Ew��A�c@ߞ��1(8l�H�._�]��!�H�J���H�	�)�JA7����*v�{�+s��f��0+���JU�s_4�,�l�������� Hۊ�5g��y�GT�iTE���K!��#�A<o���ȧ0$�p~��g����)�����G8��&|5[Q�_����_�^�^V3`�Zj�,�i�g�2E�3P�x��.fFŇhC��n5��@�I�	c4\���� 3OC�#J :��W����	���˙+z[n	���. g���KZɺ�	L1rߜ�^*�*P��a�挜A_d9WpF)�+��rT�lhϒm�~��d��Q�6��LȘ�<Ǧ��F*�´�7`�Ӻ* }���Te�������p���~�^_����I�jP�L�j�ѢCgx �kW|��t7�ǑA�h�󔳧�r~^a��I�6��2SI��Z���9��ذ,��N	�O�ˇ�,����ֶ��s@�$�8��
���k\_m*�3���'�E�8���'�cg�:t�Ti0�J�Z� ��1=�X0`y����6S��*?*�G��%ͦY�^0�3���7$�~rzq��s�܀��3�?	��'x��������)��O�m���F�"��Q�x/,�^1�V�����$��|�^X0��q��{62�m� _�k[Z�.�F��>g�U-��|�0����2�4��P!a�}~�8 �"ɡ���٧�42]h�~��D�bmQ(O�IfvŅ��xƖ�!*-ݸ13�p�v�[Y����m�ot�@(����sb�G�SB����1䖙Ù@ ����ML4"KaN�
s&{��-���5J�=&U�l����"��sZ���������r\j�{��^V���S����xő��݃Ճ������	�?��]]�y�UB�@*`ܭ�`���f�6#��"'#��ա�=0m�����4��f��P(Q-��y�j:וh��O6��f����P_�v	��"mf���!T�����uL"�lSK��B4
%08��o���S�6���HD�Դ5�����@>B���w��- �c_�-��83Ā�}�g�ѫ%-q�l�]TW��'b�o��9t6�L<Ұ���+�Ux'�Ql.﵈����IV�/�*��`�T�f���{,��`��
c�v𙻮َo}��g
��K�Lw����m1��a�c	��T;.K�U��v�(1/΃�K�b�I��2=1�	�jn�r=�{R{(|w.��+�oS>�S�΂p����s�`|����װ@���+�� >v ��ϣ�ʓR�t`Խ����zQm�(Vҷ�`�I1�(>\[���Z�{�V�,Wq��BzA�wU+T��k��eb��n��y6���~��;�Z	= ���W�$�4��ӟ��nx�u@����l���4�wO�*���nOe��q<����l�C���[3�BVG'��k���k�](i�Y)���cd���te�"`A=1�?5'�$�[Q&�>�����	P�$�b�j�R������@������k#ܠ{PK�X�f^�Y�h��m�i��,�^
*Z��zN?����]J0�)7!�L�\Z�S�7�!��CU�d�1$<��{hL���c��Gʖ���
��.
��-����숈M�fSm���>��׎_7궈'�u��!Ͳ�ʯ��w���fS[�u᭍6�$d$�G��敝�<v��爁�Ql-�@��d��̂һ���^ҙ]�����[#��֭|2)��Y�)9
��"��UL�++V��;�6?����G�B6��ԥ����W-oϿ����qw�:0A/rg�c�Z�ͥнv�����`�o�ç����:z0ѥ�'*f
�WU���Wa.=�[��0z��|���]2�k���F��A��Q(:����B"���<�NE�C�Á����	_3�7 ��5U`�1/�˙��%�Bf�J�}y�̤�G��B���,u�V|@�f�_k�j�g����2 �[�%'f7�#	h� ?��ИmZ��!M���#���y�I
= e�~kv�=+i-���BqH�<!��������T�h`�:xծu��Z�����.ª8!щ��9]ឧG*� 52�vB���=J�������FdZ�+6�Á��w4GH+�8�4��s�-U���G��V���{%�4�*��;k��˝�&w��罟2�~GA�\��a)q��em����:{����t�#��U�0��j�a5���|�)j�z�`��d��҆�h�	V���i��������g����m�]Fn*�?���x�V�L�0"�[6��O�+bK��#t��Ģ��׾s]� 5!W4B+�65�>��o
uu �
�~.�4��`�ceL �D %"2�q깟M0�@V�c�#.�A��� ��3NB{5���d�3��'vY;�	w�w2%S<:rbFj�b�ĒX���['3~w�e��_�-s滐��]`K0�8�ԋLv*�,�H����F����E�?���������o	�
D��(i���WޑO���' Se�g�$g�<X��j�^~N\nȖ?L�Ȇv��Ӓ���O8Sl��ی�Ů��UZ��R?�
g~��ȳ���%8���w��O�G�ﭵ�~377��4U��ZT�Cs��F����z���kcq�蛋�ﰾ�3��({&�gG����3�Bwi�PJ�y�cs��HE�R�|T빠�jέ���������酞��O_�v�#v	�x�M#���|�Ļ�
 �9y��2�o��虴��y�ld�\���FX��s�8��/�V,N��̈́�ȇ�����A3��a�����l��ѲвpLآ9��q{y�X���N��>)����/t؞�,9� �f}���%G0��Y4�*(+g\+	�V��p�z l�*i��������a����[.�J7���R>��a�(5��3&ڱm�����`RjO]��"r����[2 �)�{(�*r�&ʣz�zu�<j-!7����/D�L�&���97>;��c��;������ܨV�Ly�<u��P��m�;h׳1�'����(�vDRF��w� d�"'���_���̓g~��
��{l�Ӷ܌]�/T+Kv��,3�\�4	�5���񙫟�