��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ������������~���aGma�Ko�^LBfD���=�z�]�E���s���j��W 2����ĝ��v�z�9��C�f�Q��e����_��{nl�pU��v�2�]1ko1E��jup�@4�c�{:����-�d�-�#���F+�,�������e$I%o�v.<`����AFO���I���ʺ�)V�v���+#��P�@�(f�w"YM�<d2ޤ���½���FcԾ-��IooOL����-ӯ�-�ߐ���sm�&�a&�ߜ?:�{��Q��P�_��?!��7�B����2I�حY�-b�wp]�{�{�"H���R�5�Ff�}rtˬgb�ͤ>L�,[�M��"L?R��I��)_�9xJ�����ږ!��ףŲ�b�T)���BODV��Lh��Er$�|�ը_�R9<ON���������a��uk�وm�Y���~j	p8�\Ƈ��9P��=��.8k���op�y��{$no�z476�`�1Wdqަm;��vN"�u
����S������ӆұ��kǭ�A��\n|L4�ˢW?�~�F�7�������%ο���_��*N$��tQ�MrR�����$�>
O �[��ɸߑoP?��uK)� 6/�Fr/��������zd��e�,z������
T��`�0<�l�������0�Z����D���B����ya��+s)~2\��e��&>Ul�kPS�<� ���NG��2{"���	`���Q��f�f�Hp�Vk,��$��  &�����.~�<�#���U�r�p�F���
����c��Gó{�X:x�N��p����QS�J��}�>G�~ko�!�9�'~蝖<A����!k�Y��z�3G&�㓁$�K9�l���ҺZ�V�����J����釵1�sW�5�|;�m��Q*`"���F����j~��8m?����[����D�����ᬸ�V��1Gšt:Ţ�҄sBR�J��8�&������K��k-r@~��kp8H�B��2QSCx��[1�T�a����GB��qzR������%*����FF���6��]�D���A�k�e��Pj��Q��n�0wR*�6ԾB�-Ӏrf۝'�ue��(cS��C?x�P�5�eBT�!�[u1R��/���l���~��) T좍 K�z�@�(
�Xyq��*���^@���7�UJ�]l������TT�F$�m�w��\ː�`	_G>.��i��������}���n4�W�8�	��Н#��j+�P$���Z��y�F�}��$_��z����%,i������@޺|�+&�$dM�|�S�$P*x�� ���+� ����pJKtE��X�&��
��_����\C7k���U������-�����9�O�;S�p~�Swb�w����pK7���'	l9Z� ��/y:t4�Ƌ@ۮ�Rz�`ϸ�z���\.3�G	�,I�HǷ�Z�k���RWt�}����Ǩ���t0{�`�\rd�z|�]�S�]�-ᆷ���,��ݕt��O�PZ;*��
Or�0���[~������I���1`Q��Ň�Sφt�
��<c��A\�:�c
��7<gA�˶�?JU�OC[�!�|���.Q�2�=�����c�"�C�Ȝ �+S���:X�M9È
kz�m����M/dV�M�7��>�[bI�S˩�*a��m_x���B��wכ�z���}�	5�d�.�"���2p'��+e�g�}~CD��*&\���M}�S��J�a�j�kGX=ǽM8*.y�K6�G�LD�%x1E��-	�wn��v������H���3��4n�,�/�_e��=�nb�:$ϐ�A���X�$�s�7����8�8�^�0	�+mrݭO����@��P���fnZ�-"�I%��f��o�r=�M���R��d�o��13��O����e��e�[�>�ʖ��~���Z���*M�p#׋��o�Vq�����-��A�����%�A)�#9�ۅ�Z]�}%cj���?E%Z1���b��4��Xk���C�0>9�����Q?�L��EدF�g#�i��$�gp+��C9�Yz���qMy��̭f��m�V��y�y����Y"�3u�0�����!�x
�CW���|0��&������Km�SO�(߀M���#A��_RM�c�s�X�I�}ܮރ�	�ohi�(	�iy�8�����R��R;��}C���d=���+D_��[\��ӸHȇtT@Gu�#���w�4�'��Ry�kT1�o�b�n�4H�����"�@bn�%:	�"?�xE�I�a�#;�P��Q��hgp�Df���s�%�]դ���z�u/{���A�t6�NFR�IV�U�rQ�!�_7��.&ɹ���F��<"�v�Ѓ���g�(�=��B~Lѵ������g�O&�J$������;�O!E�Q���{6?	V�rٔ=�����a�(՜����!��vM�^�������xp�Xtx��Y���vO9{mҷ}�1S���Q��Z��T7l]��T��=9�,3q�N�IJ:�`�ad�ʗ[�je+�[�&���I�`�����5F�>͘	�Ns 6���_L�&�[i�)3K�{~o.���5����eԮ�b>���s�V���j�岧3氩ߒ+;��SE������7�C����Jw��'�ld�2tL��90vu��'�������h�!��5&���/Е�<V�Ri�m.����]I�j��+�d[��c�#İ�!�s�U._����m~!SiVEμAPL17b�,�я
�9�"L���d�3���+c3`��l����Af&�wXغN�;��3��Li�l�Bo8y��	�������8ege����[g�p�k�\��0�w�ʉ���K�";M��I+��2��:����F����!4f�����W�_sa^(+�UKrӋ�h.��8�z�ϖ�@�9o���|b�6R�%����h��D�TɬC�.�M<Z5/��ڲ�n��V�\#^��	F��u �Fwo(6��AR��T��h=�����B�meN�V�M�x�z��.���Oy���`BH�'ʕ�pe�G��D;-sD�&�(�<��Gh�N9k�ռ<��*��+ϚL��RFFqTyY�I��#/�U����b��p��N���H��+��w�x�`[b����ҧ�@%�b>�
�|PA��+?�/LR�L�eD��B>Ř�7�D���W�"t^�J����lm���謼bJ]������h���Y+D��U�HY�'��v
k�%�q[�+b����Ǫ����6W��軜�:>D��S�Qy��O���*8;�:I��ְ&��$+JTh��ל�&���﵎�(�G�ד#�J�Q���K?�ɖJH��yLq���`"�M,�|�J� Ƶ�4�<��	Nɉ�W����aF#��IW�
@ 2rM~o�l��N��,^���YF���]�t�LѵrCR^|�j)��A]T�!��C����Jx����+��}�+:�?��Q#��&�2�i ho���`�7=�8*_��Lp�ڛ5�z�Q#��k�!�o�0i�z�X ���[������;�T��	B�'p0��^���/9�vS��z��-l���g1�~�����<>��C�sF�ezODqG�x����) .?��Ja�E�is['���mȜK&�6��n:6x��ȷ:��c����Y�������<e���V�L���5$WlA;�x3�~KT]�Ô�̪��pue�A��e˚�:u�
�}*]4Z����8��R�eZW���H��+�\?s�T�����
Փw�����T����ا���֎�5����+�
"�Hk��3�{�l�M�O���c�ga޽�1}�C\��"�W�wG����p�Н�%��m��|��-��bs�V����?�gdQOX<�6A�gV5�t����b��K\c�1��M8����l\�`H��b�m{z��s�|�}�K��o0������;Xb8F���&b3�/<���@����yM T.���^+�5�� -\2ЪV�f5�4��c���O�K4O�e���#5�Mz�Q��f�T|L
��!��A[�ʙC�u�����t_.�I+���xU����)��g�$Z�,�n�Onz���]U�K�4p�@�wS�~��%4ڮ^U'�oJ��˼:#�J�+��ٛxْ��g�P�i0kbmZ���Hg�Ċ��|����m���HSxp���~��Ť�һ"�T�����ŗ}�<i6�_��E�m�ʈ�� /�6b�:��V2�V'�U���w�����}>���!����_�.����򺇺�<�fOʤa���T��yi#P�k;�JDi����?@�r*����CU��7 >�|�pIa<��5+�ln���Zی��#�'��Q�}�"�h�:@����Z	D�=�BF<�?��z3gV����;��M��ϳ�!kX�_�j��]���v��52%q��G�I=�1\*�bp�~v��)j�Ե�������aSF���66?�v��!р��qu�A8y��^ԒN!}����ː���N�k �0m���R���Pr� -�ǁ��#J�����8��zݤCw$��NU���(���])�{�S��@H��9h �N�kR�?Mi-�p�8���m���
�?�Gv��,���٦�����ٻ��b�:J����u����5#���c`�C�s��K��vK�B~M�~L�r���܂#I�g͛|�Ki>��u9��lP/&>=��W�󀩉A�t,zh��g��C,�<wF�{�	�4(���A�"9v6rQ�0�6���.dD��$����>]+��3�TF9G���vՅN�{V#l�v��B4kx��P���49�qy�?�(x0���Q�.{�pP��0j�Z����[Dݳ}.�FZV�5���h����_l$r�ef~�L���wy( t�Zu7g�e�WX+�ͬ�Vs���={ ���lƷi�JU	�	���-P
轭����6$l��c����6�LS��������&þ��Hh�Og줁��֛�艬��:X���>���4����P�}�N���y}-�ɾ�W��q��*�<An$��0	��U,���N� �n~S���P����L���F.�!��넄�ӧْ�M�ʴ/8ڹS�{�����.��e'8B*UA?ɻ�e��|���3%��ڻ��,I�Z؊q�%Խ;c���Pe�jU��y
)��DR�z<��\2�H�[�|�t�n���fŧ%�S �!��·ɽ�����M�<�����mv}q$���M��B��W&��CH;nlmѥ�1��].�2wނo�jz_�s���>S.�ᙫ�T���Hq�������ƺ�Rl�=̉���*^�q�~S�AW����wNB+��%�	)���d�7
Ǹ���-�����E2c�<��{�'c���Ges�kw�Cf�+x�EwH��.d�@�^�Y?��°�cf#�:���B#�4W�;h�������%ғ��I��)�&�ڮ�zk���6�b|U�8̾�sɑN��e���G1Eq���`�`>��"�mƿ'��h�1L;c���Ec>�Տ+�>��}�v��*<���|���M�4]���i �F14�S��5�����ϟ�`�i���D��u�	(L��L~��+ŘM��Z�W �}#2�+�v��
��|�UÌ=�9���~��:xHUh��7O�rťp��C��͋���m �ygw�g�J�n��'�Kf	e�mu=��Cw�T��F��}q6�nqD���g�!.�
n��=�wK�H��Ϸ�-�4�JԠm�ܺ�!w{�ذdeS�L�4Iݱ]���BXɘ�x���S\��)��g^��'�υ�XR`�j���x��)O��i`@Ġ�y
7op�/�J�[(�	���k��s1-�8�����8�<�4�Ё�,Ro�6V����/fe�%��dN5�Ȼ���B3X��������`wK��b�©I�iٛ�ē����-��a26��Z]�)����*��T��IQnρ��-��b��r��H���1h�Z�-=nݛID��m��z�E�4�h'��&s��ˊ+��GfK.I�;M��@N��"����3r�F^�M��A��D�d��'��R��e�G���?vܤUWY�Z�{�@�����g��_[���tmę�X��:ڊ�,g��n E��H\B�? �\���}Y�c�UT�a�j��H~im�fn:�0rr���q(���A�Y��syא��Ug�̈�OY�'�UI�J7�@lK���+�i �N]�����{���Q�HI1���g��i�2m�-$#�c�uxKd�8�s��e'�Bp�֗�c5�U��]��?$(yi�Z�mVX�u�Z��g'��N�%������a��^ۂ������施�	��=��t���
�Q�d�3Z�����́�%�#c~�	Ej��z�f��*���Jx�"	�{�JF^������o�D��J��ӆ����	��]٣�Dr�A��ޗ�r�0�uYL]�٠�(=��\=c�ڑļ,��hۡ�7�I�B�/�
FX�����g��-�y����濠)xB�}�m����s�a�Җ�Kn��`�g�̻�҅_	`�!\��5ҕݒ��M�Ђ9_Ɍ�Ӭ��W�_�h
7Xm�Tp���e�{S�+���J.�B1E�q]�\��YOh��^��BF�76�M� E=��O�>�����g��^�X��i:���m�ML����@ğ/��񊡷������|�b�Ol�6�Ev�'��\}����.��H�hK:�������A�u�5qIA ��`,�G�.��|�?R��hUwΣ�n�3J]�砏�V���|	j1KϩO��X�)	J�"�������E�j*��*π5e�lӌ��ϩo$���LN(���4׉¼z�8���w�$�vr�/W�m�݃���h�/�p�2?*v��'B�78Ą@� ��ֈ�'_E�Rf�)&��4H�9�p�c���3��qx첃��2D���T=h�R���P�0�d��+2�l���k�w�Y��mh�L�^\s�/��_��p CWn����c=u�ȓ��)E¡[��&=|ㅤ��{P����f��de㒧��#��ԭ���A����=wKro]�y$������x+�d֊�l
�����"��R@����I?'J��L����tb�"���&�p��l�'�Ö�nTY����%��n��,�w�ǻ^E���%E>����ς(í�j˫0����c��;+��/Y=�؏/�7�b�,g��0-��y7^����U$C�C4J��=d|�0!\2#'��i-kT���X�P���je]U��"11�zKۥC]�a�ㆲe�j�'��S�X �2�5�cc�w�#�x��z��f��v���r����> �u�m��a7X+hظ@�zE��-5��H����ɦ�#�5����8r�m�����n#�E[حk��i�nD���8��Cs���_+=�VJ�Ӡ��8ŭ����aUȉ5D7��E)���H5���`)�>��J"��a�0]
��X�����KoR~ȟVM�y{_A��z&�Y��:��6���s�<*�޲ق�Jq��������/�}�����cm��kF����!Y�-v��ZB��ha(��h���'�$�cK=_<�s2�軁�`�Jn���%�`Bq;��9��{�q���<$+�L�/$9��:=��c��L�� �R�0���
�m=�w!k�rwb-w,�d�wrCV^�'7��Ve����n��S#��e/}Ǻ1v#�/ ��ʬ\f��!��Z��۱��O5w��[���l$w��N���5��]uq	L���:n:6���*��v�a1ub��V�J�J�ʱ�����F��������$J�N��Q�l�M����t��;h�D� 1�[�!L�A�	"?���-��ɇ��&�^�$��:t;�uc:@�+ueȠ@9��t��wa��-�^5�D�pt�m�@���%w,�[�CXMv�@�:\�gtL�LУ;Xs�6K<�AI���x�4�Y��bqT��:���R�P�����m��Q�o#݈�2z�a�5a�1j{t��^���5�g�����N�~"Z�3��>Y
l���,e�FB��,�H�	��;&��x�do2�ƌ�Y���d�㐑���|Y(���#��V�O|Cn�4�����¥��2��2Y�F� &������@|j�� ���@�P�%^��3��F@2
�^T��e��h=4k- ں�`���/,��'N�,�[�R�8�,uG�8uW�)��Y�+��=���6�y�Gu��G�����7S�D��(��]��3�[&Qr��D]��󽸐�T'fV�8?�XK���MՁ�#=S4.�z	�X^V���@�=ކ��hxa�7t&�4�̗_Xh>-k��7Q�Υ[������ގN����	�>���\�8�J�&�ˁ��j�[�k�z��Q��Ȑ�G�)����綑0�q)î�� �N��S�7�����b���� ��ǆ/t��%1��3� >�IHM�Y���"{�lNiT�ZW�"63�/&�g��b}�;�˜�OɆ�WYG5R$�7P%V��;x.ꆓn��S۹���
8���n�3z0��/���E��Wc�C��.�zEf+����V��t$�XBD��3���K�<
�A��:t	��^�X2t�������g��$�W�A@:?��ܖ�{#�j��-��]}�N0�L����<�\/_ꌪ�6�:��O�-���e4O$r��*���٧�pS�:3R�=�O�];䐐�p������Y�V�xp7��U�إv�stvy�R;�*�Dz&f��`�4%a��7�����&���V��Ey�"g��􆬳�+o��m�k$}C�o�>)O$��!(U�Z�>/�]�$�)(�m( +Y��-�ߐTa�L�g��Gz�������z������v*3��:�5D���:�p�( cɿ�V���p�R@���E�f5Ϸ���
��$�_��1��@̴�-u�ϘE��~ �}彗��De�h��39>�Jw�T&_�be�)��R��'���P�0�ȹ��Vɓ)�f�QQ�n� /��K���J]�ɰ�������"x,`�Ճ��=��˭ ��g�
��bv���vMmE~�r�z�/v23���G!����$w:�{�[;�%�`�ͩˑ4������.�;2MM���g_Ym����˙���K�@�{�����=�0.�K:Fb+� �
�LO۟�� J	��-����ɕ|�3�Mc>�IB��I��|���C��/�%��\5cqޝ�l�ٺ�,��6�s��U�S:N(-9��2 ��|Ӈ�����Y�3=�^�KN �g	���Q�k������I��P��@3�-޼��2�Z��X��c\���[�fɳ�Ax�ZAw�y�w���Dn��{o,օ,k;S�kE�<��0MW :�X�L�L����P;X��z�1/���9;�2�>�N:@�(�DW-2Y"a��rG�9��/(!���&O��ǋ���?Dӻ!�q��`��
п�t�;Z�*M�
����V//�mNGS�PsxF��r��n�8dr��uC��>2�KZ����l�v�1���32�����4Xp�ޫk-O���[���@���j�� %�irq{Oa���4�;�Vد�;�-�����x�!��*o�P��J�ҭul�;s>��}���J���c{U���
ۏ0x�3I�I��0�v��+��kS��k<N,.MOi!?l�"p���Xh&��
h��RcV��r�t_hN�p5���%��*2���RP%���[1<-��Y(�h|�%0�����޿�6k�L���M�]]�& �0 �1�������|o��nl7&��c
�Q�R�Uޖ�3ڲ���T���Jd�|�{w��SD]�7B����Ū)&����U�����(�쐥.{-���SL���P[X�Ss�E�J�U�ܱ��:ޙ�:0X4���p�pl��W���ak���`�z���0���whdz|�������h^<*~�46 ��oT�5��HY�3(����v	��%��F@d�n���� �8�������351u�1(2U�Cǀ8��.m-�����F�Q�����s�������	�wT?g����ݷ���A�G	1f��Y�W[PY�+��|��e���)�BÛ��"���� ����P�s���N�dJ�� �'c�_����gq�t�2�<r5="���MBeRW��0	-j�iy���b�c��S��8�n1
#���� m۱�q�P�bA�!\%@�ԯ���+��Xx8��ݿ^� �(�-�7����=^�jtq�f�M��s1O�TW���bYl�a�
���X`C�[��_�[�D�j��mNu�<DN�g�Eҭ	����W��i�^�å_�����񕒽������I!b�=��	���Skqκ����u~��#?�P���������]��fհPI9!�鳝��E�Q��Z�	�
�5̉�YC�����n8�fU�D�V��`6��D5��ǚ;�.d?��p���a&�_�Iɫ�"��>�&N'Kv�C��(�hM�k|;�SQ L,V��1A�:��/c6!T�V��r��S�w��x��|��F1�$��-�І e�$ag�T�4>@&���E���j�n��&��0�b_#�MT9�3�8ɟ�3r�<-P	A�0�����0�W+W����ւ���I�N�d��8�$�/��1 �K"oI��;
^N0""�+�]f�ͱ���q��i�p�S�N���:��n.s�U�_@��JӇ���;�R��)���/�(^