��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ���������>��y|'NԄ&��p�����1Œ�l�~�RF�yX��/�;5ec�A飫���%L4�lޮk�v�r.��B�q�]Q�^d�W�U�o}ܫ�l?.]2��c�c��[)�߻��;7��m�V5ݩ$Yx�S˗�.�~����Z!�2�W���F�j�`N�#����~��I�D�����H/Gk{�����AZ&����3$z�?6��v,Q�<Eo0�L���n���$TarcN�� ����;z�f�v��u4��!�xFw��W���[���z��C�RLP�h���D��S���>#�	t�H�3��尀4��ҽ��2�xO?�˗��4}����
# r�0�ˎ����j���>!��� ��]A ��J����	Pxjg�G�WY���@��T��3�k��=�8�f��� �s�{.\u��� 5��.eS�ѶrF�0o���7�6Ї��ߎrH�o�mJH�ɇc�.6��o�"黚	V��8�f��7f������@#v�W�j��r�"C���	�b[Z����`{`m�:�)h�g��-�/J�\�A�?)�%��)Ǧ�Ar��M�0���m\��tm��l/L -��!����[v`�<��Ӣ��l��η[z3�[*�?�t�UC�� `�W���!a�=�Q#Y��/8�B�0m������ac~�e�>���� �E$��e�ի	��i�h��Zo��7w��Y��_���Nl�UDx�ޖ�%� zf�k�*O3�ψ<	�`(ڏ��S��b'Sv��H9Iq�����[�'_Ts��~ ���5��2�u9OK��U��8�d�����zj��΍�� æ�'��T��`ÙZ�]�������H.�o�����c.M��p"#��(Ħb=&�3�?������J��  D�Q��.����JξC|^�7-��-bW����ջh�����"������tbh�`w4�$�����r n�� �j��I������Jyzi 
���:�A Cz�x��?͇�d�ՙ>&��S�H}=���z$�}���s�3���p&h��-�Ǿi�q�Z9���'����Jk���ud��qf�ϑ�Wb�\�Tx�ҼHFw���:HN���@Lu�BL��}r5�92f�%)�Ă�Ds9�W�_m�J8�Z\>,�'�z��&e�y�E�(����"��w�)����˺�k�r��瑕�+�����,�);����������ÍKC��R�.\+7��s�-joy��a]y�x���>\��z��\ח�4m��^p|��ˡk��x-����΢B�-��e�2:�i�Z��j~���3}�:����O[�+]7ɽ���Fǌ�~�GE��ȣ��E�<�?�T���$l����kŕ�`�4���Z�=]2h�(5H��B�?�B1o��q����z�w~�GV�rO��d-e8R{�_]���'�(E��Żq��ʨ&��'
�1�*�sÀ��g?���0ń�IG5���I�۝��1��@Ᏻ�p-US�S?qexX;(�[�����&����:��bL����o*�ZvG?N8!�{�V�6zm�c��?X���x�or�3[Q	�\s�.�@�Ƿ蓿��G ��X++�'�d�%u�}�,+�:��TL�8)���O�R���dH��<EL�Z:
S�+�����7�������=�([��fQ�~=shd�̐c��@_<�>�<�����!�i�n���_�b�+K��
Oim域0��gzy������)��8�Ei���v�*��Z������GYG��$E�g9�XIA�g �L^R�9>s�����o���8X��*�v��ӄ�|����H/ϠNm��mП�-���}�^��lc��ոa�;`(�BHO��C~���>�B���(�G�#��������f�	���ҤgYh�ٗ���,��V�-�y���GԿ����<�y0��U�
�8�pn@���s�v�� �����d>_���>��:�(s�_��ݲ����
sP,9�H��_`���۠
Tc�a�=�]^.�c?���i�@J�7us�ԩ>���PA�c`�;_L�5�i4
:�%úC^B�����'��D��+�A�/"b�1�YˇAr475�+'�D�7�B�?u9�з7���~��fs��_��hy��em�[���LL$;0���C0,9����5�ػ}tFΥL\S	.�Kh�ʤ���l����?)io�	D�"�qZG��Y�Jmn��K��J$Y�Ѭ�S�GV���5�]��D+�-��x�zL�j�;3
'�[EV�I��?9Ċ�I�����@uP9J=�����@T��lOj�W�9x��j�	�Y�8�gr��$����hO ϛ�MH���X��w�i-��,�X�ٺ�T�h�/��1[پ���2$�|>C~�Q=]#���+JE�u�:	��b�V�嚊ͤ�
o9b�I^�TO�7��*5���X;�zf��7�}G*�P¿�g����0_"J>�4�`Q&��]�i����n�<Lqk|�����u[�h^=l눛Nw
p����9A�%Y�(��`^U�f��[�AJ��N�v,�	���]}����k�Z�eLwNњe�j�%$ȍ� M���JXf���5"sD����rxf#���.4��� �a�Vp���E�ӎ/�tz�8<��U�/���/>��pD�*�s�����:��f#~��"�x4��D��������.����}]���RN$7�dl:��j8��ע�v��Gѣy�u!>�D?JEU�տ���|����fI��Խכ������V��l[�L=F��QN��Oq�`#B�6Eܞ������y��!d*��My ���D9
 �):7IO;L��˗��DI4�0�U��-Z���A(j����w��h�1��ޫy6t���xpT��Z���7X��!Y;�M����B�f�sX�͑[ެ4ֻ�/��z����;�Qn��W�c�`�w�o��4��L�b��cf�5�g@�ٛb�M�]��xs�ۺQθ+k�¡��m��8�ȅ���-%�0�2�2����,Q��șE�S�{c�ֻ<�s�{���f����*6O��.�
��M�*'A��}��kl�ԑ��t�M�JB�0�q��S����Ƴ�|̕�2�+����ݔ�r�-N���.�r���+�4�f��U�l>k�ĵBj��ޮe����]���<��GB�p�ꆃ�v���B�`C�'�&�xE8<�I�����߼�0��e�*^�X���6H3g_T�0��3�s�9]�����R�wt�.�.�Y���Wd��֯�����a�G�Zl��,���R�1r��H��V����?e�%�74�@ ̂�&�.������=��Y�C����Ũ>̽|��݇�k��}��.bv�L�y*cR�K˸!̜�&�){K���o��`m�JDY�"���(�cP�;]ݚ���ى���;�R��V��q�wMV�=b��p�I��R*y�4Q�2�"�������-Լ�������y�,�ӡ����鑆���Q4v�����U��{P��<�,���'H~40_���/���e�Z��\ �&D����1≝�B�M�1Soq����d�/F�2�nk/���͆���2�\�v|�q8&��^s�[YNw����m�c@s.�ARm�o�]��Ri1)���	]���5x�fb.}����3��|���֞w�_�����{�k�`M���T|�����H<+8������h��iTm�c��T����F�km�s�6�dbӲ���!i�zn�'�d����g�4O2�����"~):j���npY���G�����ekW�%�K@�|-)�M��B	�;�^�7ɞl�F6,('#"�������Xj��p�,uڹmF�ܮW��I	Lg0a�Xq���(������T���������s����9�ұ��`���E�P�[o7T�LI�F�FWBw}W����h���5/����\i�B�� �bɩ}�����q�a��38���Q�+��ot��_?����6N��Ea�´�,���/Ȉ����9Չ��\!��'���&�X|�Z@����;�� ���I�9~ �z�c����ś)|���ҽ3�}Xn>�d���?�E������W3DSG=����D.��~'!�Ϝ�r*� R��t}{1�E�4�t�S�c�7�4qe$n�^�("��ҾM���Gm�\)0iD�2�E�"��54IGJ��wM�.EPސH�ұ왔?V�E���θ?5��B�4ToJ�U�q��ӟ=c����������ZX;'^a&\ �5g�U�köxgܮF��BϮVP���1{.0T��DԘk���Qx!>¥3׺�yj�����G��9ń�ki��ls��K; �*-�@���=� ��P?m��3j�Z�D9>�+���}7C�f� ^!�T�|AΔ�RJo�ՙ�;�W��MIٱ(�H���E�5Lu�����Ȳ�(��3:W����8�@Ii5�ϑ s�i,N>)�Se�Ν��`Pi�w.�"�K�|sa��1t�����P��%×��2M�*���
�c?nCFK�Y�SY������Zf���CL{~T�M�>-P�|�4Տ�9⓿�x�W$X�w�{I�Y@B�ob������}��?�)�|AB�x��m�f��%5�|�2Bt���q����u��5����F�-��f�6{�>��z��$�-�F��*5�f����(DK$gh!U
�s����[K�Klh:>�E��?�:�d�i`^�v�e���l+ aX)W���M�jy�i�y��g�6�R�̮�c�JJ�YR�!���H�P�yVQ��i�U��͚X�UX.i;����zށ7�wZS����}�;�ޡ_U�'Wo	B�o��d9�E�������]��z��aUK�l��d@������_07n]��%�~P���IS)Ih��Y���`9�1��p;��W1G��3�~r�e���ԇ�bZ�r%N�8i�S
Y�X�M�>ܐ�f�>ō���.�	t���)FK3�sO�G*e��=�Cԃ٪����'I큱�߬:�j�>��2����"�K����±��͹�u�&���r�n�=��x��]�&�O3��i4f|�yN���F�i�#�0��ci��Ӕ҉T�~*�!RC�8Ѧ���҇O�A���`ܮ�i�)�UC���QЙ����0�>]Mj��Ɩ��b�����R��m�v�m�@1��r龣4�/?_��V���� 9m�)�xS�[qs���\�q^�r�w:>OV�����9s�:w큗�8��\y�1W��6~�_���u��%�Ӑ�|X���L���~�,G���^=�q残�P"��4p܃���P	�la|/<�+ҟ��G*K EA��w
����A))X~ �R$���P��>Dk�W�˟��0�l���{X n)��p�B��*'Y8&����28ƃL듍���l��?[�s�KTg-6�iΟL��]����c`��k~5�'��q2J�W���#5f���f��2�j�+�ư�{2⑁ĉlI�凿҈V�����1.��rᎾ����A�[��%�_���ބ�.nM�f�fq4͢��y��:J����ՍD܋]�H����X�=�qئ=zN<<0#��y��MT]��;𫒣=��m�4�?3ϭ��H�^�vI@肱�p�$�[#64�Ď=E�}�'�&�}���?�}��?0�Q�9���)%(�L]Q�k�O�.�������q�Q��U�C��2/^�90�:��4���RX�@u�hw� ID�n�\NT���FVm.�	b~�w���N՗������^�;t�ax ���h|?pJ<�kIw��+���O��h�f|:�_;\���d��g�,hn�2��9׺��Wt� ڈű�dQ�j����,Ew����ZdOk��a��ܴM8*2��n:��</��W=�\_j��"�x��~�����q�ħ�&+��F$)Q".�S���n���m�Jw�$.�j�i��qk�/k6N�,K���CVdr��1�(���\v��.���A%l�����9���S>6��2��.�����q'2����@�Ny���?L����B�\����57��.��FQ�5� _�,}*zd�(�M�G��"��ﴤ�{�4�RQ���QIZ-@��	}G���t��~�"�Y6���(}�ݤ;��, DA��7y���.>튲�,�_��Me��fc4¥A!2�So/���j��^������Wb�a� U����16�!�� e�&��oη���r�e���#L���9Q�/��q��eo�r�qUB�	���|W��_O4��<��	��I����������$�	��SA:t��:7Sw����ץT���.5ڼ[.��=�D�-#
򀞊�@G�R���R�K>�ж1hA#5[��H>8j�-���B��[S����P<�q-\�t 1�-��6���o��m'/K����5S����s,�6{��.l;?��>A��2�� ����F��!��H���v��/7R�)^x�֗n��X�g$6��n���x<�l��Š��?U�3�� �V
D,�|�򅊢
b����\��&�j��ҝ��f�,qj���&s��d�Y���G+� ���Q5�����[�(�!����Rh-�������y�\N���W�N���X��{|o�C�������{��a�3������<%��XZ8��l!*����<+�-c�_N~��U����]��t}볿ǔ�;������!2t���&`V5��Su�`Kf������B��Ǫ�L�:�����6�M�\���;{�������O�*)���۞�7�h�
	ih��v<k���M�;�^� M�7+:m�L��V:	p������!5���Y��Q6�����wB�۰�y������f'V�]v(�.>����*��TŪsBu����	���C9 ���?Bqw��T��n�@r^�u$��tM�\����R$�q�b ���X������Ko����ҵ�l�4�����@o<��п�L���|D�Ⱦ�m���WۀJ�^����Sv!_���J������R#Wq�~2,����":©��.�ۖ���v3��| �Z:�L�W#����p��&z_��*A�Q6��ĵJiG�?i��r�+�� �t9�DW���2�ְ;�W������x58��*㌍�I�?@^�T�3���0���(���,���@�&��6^T�5�5Vs���F4�=�A��m��jKZ�P��i�ȁ-�Q�`M2D�����6.?vN��鮬��L:�����#�o����&9��x
S7�C9��f"NTR��껠>9wAz��{6N���u��O�mX��Ay�����m�5�@_�?����^���r����ݗ�\���p��d�@Ы ��L��� �S9�C8ځ_�g�w/\�:�`�Am��!ϴП|3����4�Sl�D�p�^2M����&�kD1�oD( �K��������iiYۗ[^�>�A#b!�X�P�uG8�ˊX�6��jth⋳�5�ˬ�����O�x��p�~M?����V/S�{U�5s~%c^F��`�?�R��N��5Z<Y��A�5��n_^�Qv�q_�.�ᮒ�g	��a��z��8��>ge�f����h5���'�k���(WB�Y�Rl�`pq�sp;���6����&?�	0M�

�M�����tb]Tn��ڙ�{���	��Ay1AM��Y�s��=$d��{�k!�F]&%�* ȇu��쨇I����5絍"�t����x�p
���LZ�&�����S�#J= �~>�7�_)��~���E��R�0G~�k��AH��&��Z��c��T��+~�k��7�gA}+�[��.�-����>��Ȇ0z��L���2���]Sb����('>�S�X-C��V��Ytz݉��� �'b����Ӄc�����}��0'�v�O%��	 � S�P����I������ *2;s���ȏ�&V�\���U�f	W��G+�d1B�~����qմ��BZ�X9�X��+�����>�\��r�$n��*W��Jh@���? yV�#�|B�T�H�#��.E��t�N �Î�� v7�����%��7��������Q]�y����;�<���oԙ��S�#��V��B���H�� �g�W<bc�9|�F�`k�:AZM\K�\��gC�������S��Z�{;3��.�F�ϧt�d�E8�n�蹾�Z(*��rc�U���{�s@Ĩ̦���M�ǈ�4;��|��A�*¯?�)b�U�_L�z�L�q|�Oj����,�
Gj�{?i	a7Zl��o��
�Q�F��`��>%s�?7��o�O]��yl7�f��6�X�|_�;R3�0~�+$ǝF�$��ЅK2�pF ��/�*?0:$�H�' laE�4u�5l����7��\�Kf�S?
G�6~���MH�b���X��wE��MG�]�,�h��Z �∆��Aˡ1jvnbm/G���]���r�Ř�%�/�P�0@�WO#F4i�x2���N���~���Ju%M��5��R�E�+)��/��{�����y�Z�%�⢈SI��'����x{���E�iً��=��S�;��5G">�r��E���ɼ�휨����i㪻��w��՘�:D�{4�2�1�P�{n�����/���H���#�5V�qz@G�&�`hⱷ�'��y8�A��o��۵��{�p�$FB�~���@���ڙB�=UlQbW�5c'�c����9o�G�)6@
|W��4��g�SC����)��6��s�ƒ�#�Gc��K�Ø@��{�]�]��k3H����Ⴊ2�Y?�������|͌SxN���0z��.��uP����~*��.�̇�����N`�:-DoIW��� 8}�oAħy	�1�9_pa��MAb��g^u����n��kz�=�~eTt4��	_�uJ�y ,}Ss	�����3�'�{x���|���@�!q�7�;;zX!�4��O쳙v�[�N�ώŐ9l�k�n�̈��Ґ��^�ۭ���C����)�*��X���Z������`Sܼ�%m�*�k2�/�bi�5U�A��qeg������@�ܚ����W��8�#0�kpزRÔ)�5 !�QQ8P��?�z��{� ���ҘXZ�Ey���y�q�~)����U�*�nS5j�=�z4��:11	jy����t���D2��b|���Õ�ܭ%���<�7�'�+rs��� 4��k�&�/�-�T��4��`;lD���+�ux�����0�lDph%����ؑ��Vf%z�~�*��]g�9�.y���е΃8Ln["J�&;���\��֙,x��`dP���@5����K�a�ٽ��m��p��������)E��郸 �R��Y�6��HE����������欹�J���ٸa#�%�������>;0������L�[�3o�B�S��ϝ���78��\
�l������5՚5WS�0����Ô!*k�-J��Ww�t2:o3�a:!�/�J��iGW��2Ba-��W�Z�<ގ�ɖk��.�+?yM��ºա���(.�n0�q�hL�Z5A�3��|AY甕w�o�o60�٘=.�~X�Bu�wx��X�}i�}�׌�	�ͯ�H���ĹFD���]�7�Ư~��q�%ը��=B��~�ڡ�|9 ���e�yOk��Z*? ZJ��_���6\Q� �r�y�$�Ʋ!]�$a��+-��7����R��Q.W��`{��%k0�j�h��J��`�2o{;ǳ�] lb?�%X��'����Є�ձ�
1���}�����jє+^ޕI���\L88�u%85wZ��)�ݯ�j���SY�W��Ѽ�w���ߎ�J;���F~F�_��tQ!�@�%4�'�m���ǆ�31��T��ǒj�y����5���z����E��q�X5�rN�G��g��@��e��?+PYWF�jYd�"�2�zК��y�C�@
�g��
k`T�wtu�U�V\O�M3I5c�@��O�f����;�C��r��������Y�!O�����}P�.�H�8ǣ�q�G��s���?e�t�L�$?�����lĲ��7h������Q�ϖ���QO학�����@����A,�X�p���	�Ou ��o�*ܑ����o�BY�\�L�9C�Oi�����/��#�d�_�;L�}�/�Ъ�}\��-����z)&	D-�_G�o��Gs��u����cT/}���g��o����Wv�Sn�����vd��nZ��a��ƫ�����,u�y�f�x;-J��~~֑����$q��P,��\��K5��&#��-o�gnH�Ņ�	�eӰ��gI��C�X �Χ���m�:\�6�����G�d+�.d�e�}���>�I���g�Vl�Q��k��4^�8M��u]|�B�R�+P
�} ��+SXy����w����~�����I�:4��D�Й�S~��xV%�1,,;�P�],�#���J"��bv#F(��1��������dt/#���!���������4��Rl1�m\O�{GM`�R|Sʟi�-p���{5�O�p��[�!}����2�|�5pև��L6�V�Bi�k�>�R1������\�9��5�x�Ir�MFM���E��g�K�|1��I���h���,��:A�?�u����I#�τ���XZ�Ӻ���2�榿�������ЉRsO*4<��m��LDLd�S��^�o���Z��PR��i�͚����P�7ȧDy/k����,��B��R;�i�w�>��n�Ž�q�V<Ԯ��8)
�n׭���YF�-���n&���'���X�|���4e4�;@a�f��^������ū�����䇖]p����د�32a<�Ҋ�.�1������"�ʨ�����n��1� ��{:�ʙ�s��;���IY��$�?���9�]��/`%��q<��;{�݃�U�_x�+�0d}�ܲ�\v��<��q�2�6?,X��}.��T��߁/�����=^c��lvif��Q�������l5���^{�׌�a1��[f.�Vw�����Ym�s���h-�+�:�P��S��	��	%xha�Z�q"{Z%\��u������ݔ�lq������P���E�0 }��I&e��B7�]�y��Qu|	-C1����I��kso[�cD9�0h_��V�rP�]�#�)'�4�wͶ��լ��K^�p��Ms�^q;n:'w`Z&$�U,x�r���S��A9ST1$r�I^�>��Pr�I	��)I�y��w���_.���dHyAB�W�z�& �,�KΚI��I������#-��;�s`�_�:f7���I�։ȶ,�K�t��,�N�I��װ�X=LEF��yU��=��v��=rR��͞+���#,��B�&�o_񎦫R����S��Y��a M�t[-�(̾N&9�Rv�5�6�L����('F�DC��?|p�T6.#���4��HmB1�� |�,-mS�����O.J��8�vd�{e����򃭨��ƉT�^������4�ʚV��d�dXѦ��5�6&J5w�| 6�TV I�W�l@���ʣָTDxA��UOtr�V���Ȋi-ĥ�LX�ʋ�ٟ\g`�bϦ�V^o�0nq�+ ������&�58
�SL��g�����^�6љ�M�ϱ7�Ψ��i������ow��vu�unrFE"�-����P*s0>�M�������B*ӯo⚃�������=Q.9����8:�G��v� U|�����5�H��j!�������k��Od[;�z-����!�З��<�:�M�p�h?�B\~A�X$�=ڍ<�P���FR}�-��=��7+�)�g�K���O�ء���B*�Ё=�����y�O�g� �H���֛ 	����t5�抳(�˒���08 2u|��G}�*f�Ҡ�(�w��C�O���O��:�������(RU��ȍ$Q\�
A:��P�`�l�����	���{��Y�A =�rPk���������t�t�s|ݼN�B���bkO<CFIm�j��s�3�j\p�w�F���
K��޻	�A$�ܫ���;�R�ɳ��E��dO+��/ť �����Ra����J��ήŹ�U�T惖[�sq3���S��z�VSW'RH�e�=<-��<,��v�(9H �����џ_�3�_������� �7Bk4,�T΃_ �p�;\{��T)�<@F���,�cf����G��a�[e�n�Yt���%�V�3FTlWm
����|�|��+�@�GE�\�-�Y<V�︇�$��1uj=�~�.����3r�x�W�z;�:��/VCn��iA:�W���]�9S�>e^ :�l����^L۲�!��/1lr�k�"'��\Im��x��
$��~����,h@�D�Y�_Zv�P�?���	oX
yܤ�]m>P1/7�7����T��-����q3ƤD�-\<�C����Qsٴ:��*5u��Pݩ[��Q�x{�B���֨����풳��J\�����ϥ�ǯ\@`�}kCߤ��u���g�1/,b |�&��-l/�-��@��X�BNaI�06�K�x�G��h��@�6��n��F�rj}�1�Yl��N$���~�p /3�I�|���K�d�-�o6�X�S7�9�����ˋ�/��6Y�p���{X�)���H��T(��-M�e����͟ݭl2<mk��K1&�q�6ǧ�SO�2��	��a>+l��?�^Sv�o�	��p�?� Y�����B�)T��Ǯy]�\l*T��<�]5(��	�z���M	�P�~�q�õІH����W=��5��r���-�����wP�
PZ]�g�=�KE�ޤQ
sK\���cg:U��"�8�G�`���O�Ԉ����,p�:Y.l��;gж�K'Az�{�1�p ΀�Q�#�9��_�.��h4��}����]��;&����5q�������h����z�3����Ep9-�g`([�Z����E�:KKӴ̑x�e��[���OdE��g>�Q<��-Sm!^>,�Q��=��Jm
�t8߿��<�x3�-D�ĞGS�{��{!�SQ���b�ʤ��i݈.���	h�i<+�o���5�ڻ;?eXE&@�-7]��W�X��ǩ�pp5�&��}moRF�'s��5%exS�l�n��!l�\d�'mL`0�i��X�{u3!���+G~�J�{#�q�-Lv�N��ŵ �xW���s�XT���?-RQ��eP\̖ǂ�7O��[x&=����h��ƌnn�}Q��~2:P��F�E'�Y6����h�w������R�E&��:��!���1��9�V&��:T���H�G&�
Fu+��z�$O٩����ڗL�j�m���+�%���� �����j��2B��f�eR��m��t*1��X�Fz1�ڂE�"�Y��)��aDl�P�T�pJ��̘�C�S���R�m����߂]>)�,ɞ��)|�W�/68�܁	z�Pf�~���z�I�b8��ѷ3��u���ꈽ�% �Ob{Q�`G��l�L�}���ے��1���o��I�Lc�E3���4�����h�� ����JH��t}���ZGP��x�t�yZ1RJఎm���2�	�\F��潰s��R@���y�����Y�d�8ح�I�_����j4*8�b�X�P�RÌ�}b�U�C��r�WԉOd]ji���= ��3���ƺ��1���u�S/öܔ�iU�ֈ�S��B_8C��S�_~�fg�MkFLQ��zr&\8]Y�w8-Yi�;�<��%A+���L����x,1���RA��|y}���8�I�?�K�j]���4�Q�&A'3��������`=aE.�n�g�G�)�jM���4����f2]屫g:�>�܅�Cx�Re�/�����ϓ1OY��Nu)�N�:11q����,ݟ��z&�ue+ͥP�fպ<mb�=}2���c�7W$�iba^���0fO��jc�_�	,��I��hϙ��n<�y��/ﱹuҟi��62^ck�l�r"�T�?/�j�~�ղŌI��=ԕ�ޕv��1z�#��	�c@�7i�S�W��Uvn̎�ăK(e
=J�T�)_��}������?�,#M��#R��� ,Q=���z8��i^O�BD�Mt�OA��$K6fi9Fn��t >SY��K��M#b�OS�HM���a�m������P0Gd������v/�VAI�J�](�����C(��";�p��0��M{���0 &��}��F:�$��wh�#���X����7��
��#QZ����6ƛ��:���ck�����CMq�g���ZX�q�ۤǻ3eN�Q~uC3AwZq���bTJ�^nڙt�֐�����\�c����O�*+����E�(ն��<���V��U$lm�q�w����Bԭ�2�Я>B�CZ�����nN���fc�uDB5��XR��wH��p��ǐ�A/^W|LP~�..��@���`����PO;<C��-^Bs11���%�m2��j�;�B����Jg��J���>gzA0�d��1�ȿ�'k�f��������j4�Z48,�A�Q��܁
7�m��������R��	�k����p�(�KI %�Ӊ��Ԝ��.?�I��"J�0���r�4�b܋�|��I��@/Iu�/�.=Qr�'ɺ�xW�f@-U`�7�N�!|��mpapa�l��&�biR]��UF�����h��8V����/O~���Ҋ�cK��I�4�_�gO!ɾ�Aׅ�
qq��R�R"0�h{�=�S_���=ver.�{5����:��L��g�h�m����i6�Y��gf�1Йf Sl���8UQҔ���$�HA��7��%����_��X�g��.�{����Bl��l�E}E�
����."�,ӊ���h SŜ(^�%�T��ƭ'&��
�r�����:�����!} $#�fH���U�OI��2oߩ�>�����5&i+��4#�ż
/�C�:t�|9~�H����	�Γ�L��*;���a1�w��E/n��z��FxYW����lD&�Ƅ��?�]`�Ɍ��x��C\x
 �6VAR����0c�z����M���f$��}:[�t	Q���Orsl���|�9�uD�כ�3B��+L��,���d����5d%�*��J�b�o����؅�j����rec���C	!zy�ߪ>�������=���Y@:@�q��l#�U��F�0:n���iP����\47QqT7h��|j�6��{��*Œ��}�H�t8<h5�Q2���ەF$��������,����`�G�h�@��$ۚ��@1Q�����vp�z�rt���g�EK&��C�QA�.��xc���g��:��dw��yrA=��n�߫$,o�oKj��g��eig�=�t�?�J�݃J4�2P� ���c���`*Q��^���D�C�u��
 ����5���e���
2A�ٟWd�@�P���̵C�Fd︂iXb�]�� ����'>�G��s��5-gO5f��1�H�z��hQ�
\O*��[�l����(;|�����m�2���U�
\-L����M0]���x�r�+���/4����z4��Ei�	�|�pgzq:ޠ�ͮڝ�򆬺	�L؋�"���'%�1�Qw�pd������۟��u����y~���� ��u��,?��O�
Q�B&��o3�j��{��> �-2�p�t��e�E3�'�F�������wOge)oD�0�N}q�h���ҐN��&:V��rQ��*��p�|F/W���̥�<W�g���b��m����/[H�Fa�)���Ғ������L� ���U��<��m����9��u�ߥ��tB��v�]� �7U���)A&{2`>�Z�郾��B������/z��r.�ЙT�T�xo�4��̌���A8�i�Y���W~t��y�%�0Ӕ�i�K����+oK/5w@!e��.~�k'䰧I���6� �m�����QD�x�
� �Osl?�A��i�|W�L%�7Ɉ�R{������Vn53�>����M��_�_�E{�D��fr2�r{���G�Zs���[%_fˏ���>Q@�0M���M������5kdiS��C���9���h��ǺP`�CL�^'B�]�Z��B(�;���=�ə
�i��b�g�Jx�4�]�"�~}��Ngt�����^�Ӡ��8����c��}H�p�L� @Y�t'��Q��������T�m��}\��9(��<8[��^��w��tiǇ��5�c1��o�;ed\<�
�K"ud5��@�𞛌�$��ؘ)'�~4��
��ra�{��?�_�秋W�����"��h	��t�Y<r!w��v;���o���04)�'N�;Q���d�zj��)rSn��Pg��JJ {���'p m5S�6�3Jjp�ֲ:�Vfw	��6U�-��Jc%�DbV���f��~���m\"��Cd��6hw�����b���e=�O���Є�tƳ*m�~��e��॔hyD�H{���sy\@��]/�[ҤG&�,��!ׇ���P����hf7k�0"��)�q%J�њ��7�\xe�sr�c����J��句�W�� ���lke����<D�����)�x�i!ɳs���9����Yء𿆎2���"��@�s��ћi�
"�_8�� +�rmorI�Ox�\�C��m���' +�^��(���s����@���83��C1���h�]�Yew��Zt����c�4	r>� �������=�ؤ}�|S�BdB�>�f'Sp��E����Z�\��=�e��Z.��Qf>���I�B[E�d�A@k��!~	��F��D�E�i��i�D�����[��:k��r���X3��^����u["��D_d� �f��N�H���*Z�~�!Bk�z:�3+Vu70\MJ`�W;���G���z�r�����6��_0!*bTI����D�+�Z<��h��\���%�/ް=V�H��r�ð�pCA�޳�� ��l��+����!"���X�Ʃ�^*z���}��
Bq�ISՉ�1��-ID�}^gVE�����E�l�g+7�&,u[J�������Z�uɍηwk� �U��8����l���;��N������+#�l�:��]�:`���7e������忧���&u�d7m�d<�>����pSE%�Cz	���Zsf�[�k{vK菥�E�䮃�ҁ�!)�?񖃝�H.�Z}D���1�T���3�Ñ�B&�N#0�Б�o»$�U��3�[�ަ�i
��V9�OFDrp4�@dí�j �'�#��#v �i��Z�h�o����5,���r�h��ͨvkN��k�0��u��0z��(���\� &@�l�F��*0���C�0�ԓ�Ja>7ݝ�3^�L4�J��}�~Δ�$$�dWI1�q�}j�N�C}�"��K�7��P��ޚDAɛ�����'��q��=A&AD:�+E���#�E��?u�#�a\�Ʌ��Y���L������fe���Ob��lN��=>(W�$3}����C�Q#&���/�hS*ϣ���j�M
�b�&����$#ΨҠ4��$�B�~-�����S@���z�#��A"����ܝ�,Z<+r�!Uq
,L�}L���fj���O�?�T|EySf���72�rd���?�$n�"���|���1f�#�P3��r�=s��9�E�$�o�����2Wn+�\�G|�x� ��K1�
d8�9�o���l����g���'}z��,��#)��,���w�c�0tV!n%������+Y�{������9ʡ���{I���|�ȏ]i�N( �w+��a���U��~|�2������wfnL���\���0�N؊ϧ;�Lp�TW8�e�~2��o����)��+?���~���h4��M+wޱ��p@y�p���H7��B���9f�F��'����1��np��j ce.�[	ֺ�O�NF�d���B���g�JG��
\���@�)����2�#���6#G�)�{�}~7c�4ޔ�'s*��M�/���"��-���Sߥ-��SX:�F3���C#󔜂�
��%d?�W�>x�����`,&�W�/�RkD)�}�"�P��k�(��*�qqO���'}Y���(Hr�~��g�>1�P~�R�]��آPD�A�)�kc�,+h9��c��+��d�e��>�.�0��1zO\[�1b|J��]�Y7ڼ��`�G�?�)='�#�=�k�Z4�"Q����'��T��76����/\�ttng�m�Թ \Z� g�>��⠤c�Dv�3%ԘL����e#�fF��L����z����W���Χ!s˄ƥ�Z�PToz�ty3E����o%k&����g�Pl6�a���Oˣ+7�B���-��Q��R$��J[z�W���@Ő�(�C)VY.���w�{�UPWU�;�\[i�W9�E7}p�؟�i8?P��f�j�iAAx;�ݜ�ɧb�ʲ����G���ws8����3y�lf%w�/�o&����w��w��&i}�z�	�v�|5���#|�QB��;���p��a�����W��Y����O��l&=~�l;��|����Z�N�ܖ���4�@��-l���O �����R��V��}�3���T�C��ø>@յ�Ps���*��x.�3U8����m��!J���B,��t�A{�|_���d-��]yN�����c�T܃^1W�}�d<�e�t4�W���Tn�Nl�?3��Q̗���9 �r��|�XŜ��2z�L������b^S����&��l�ܻ3��ϷYFjO�u�)A��?��5�V�1�$'����x���/���emڿ���83���U7Ci>+��!�1���q͚Q�#�1�Ʈ��y�F-��Ո�����^ռ��y �8k��S��4�?k�_�r|����.��T����eW�C2���� ~�� ������4����G���uS�� x���i��1g�V����g�#�ݞ��L>�䌘�3�pK�D��P�Q)�����#D���e�����
�#m(�+'%\�� 1�UEt&�#*�-d}��FR)�)���;����4g���Q��>y�DO5U}p�Ӎ�E�	� �+��'�0�
�~!G���9vڧW�w��tȊ�sv���{�{s�:�K�������WՋd6,�Sŭ/��,�I.����@^�����ņ��Gת�W`&W�D��LK��ˈq�}Yz"sMU���9��77�ޔG�;��=��	u��BT&-E���6��Oc6F��ƕ�n�r��G'*�Ȥ�C�,�d��j%�d�6\�_O$�p)~�����g�O[	�
�eӽlG1�,�qR�Ɖ��{ݑ��D6ʗ��5dKQ:u�(_gs�ػ��,��@�<�V�`#qO�t�|x8ͰgM�����F��.}�v����\�\8V �E�k׍�$ҡ��Ll����Wx{�b���n�>�����R��-`s�ݨ�����:��,�7�y�G`c؇T�ޒ<�⿥��;����N��a��q��1��y7ҕ8�߳t����D���!��JJ�[�yʸ��Q�9���n	�ݣlH��\���	CO��p���ğٕ�� ]�I����@���H*������֔�"i�#�C�1�s@�3��,y�5ڐ���[7�����hҭ���;3_vݺ:3��Z��N�gTt�_	Էt�EZ�]U��L�cK��ʯ�#�%�"*}�~�:��тJ����/���֦�V�@D��,��)���H����Bw���8����a.��P!*޼K;߰������`�ڌҔ=<����N@�>�|�6�D몦s~���ռD�T�c�����y�4D����G;��,T"4�1#�]���3FE���D3�C&2qp&ߏC�QUT�9%f�n�����U���GiF�7�ǅ/^�tiA����3�`��mSE���XAlO����t��uK�ߩc�9�-�zgJe�k^EEm��!�t�=�t�i.ڄi�����+�Lcm�����U)%w�-�.�B�	86�Jw�H�8-� I����9��m�B@.	������4�����9�I���� w�$�S� ���0h9<��N����[;u��(S0��a���c����wq�8����X}&7�"���n4|Yx�bfA����*hN��f;�`��[�`~�:��I�B�f��̹�1,�VByMk�4&�eY��o��s���W��~"��<����)������g��P'��~�{[��&ذ��C&M=Te�� %[1�%ą�?M�3��>ۧ*�t*�p�g��z���$�� 9��|f�>m��L.�B^3��<h[����`�P��������K�EI��+�t���eiRH��=�-J�|FQ�6��A崵�ƻ�$-�{@��5�V6[��l^C�nr���j��Q�ɞɗu��o�\��oa��0��y*	t~� a�&���d�L����"�*���I��&49w~$��~׀jc����!��n��q�*"0�O��X�a�~�/��-�	ʷ�YY��H%��>��nd5^T���ז�9öGY�0N*CM�o�?��E�?�د7�ϴ��֌�-�1�E�

G�EM��x�-��5�� �(�53Ă�B�}��Ă�Ms����y"�*9���Hr�zM(�T����h�KuϋLe���W�������Y�����MJ4�{ZvYT^TB�5Ws��F���s6�Aʌ^����HC6����_3f�z���5�&�/��i���+?�ہ}���aA����WZ�5*�!P���Nb��І�"���fpCu�F�u���Gx�Ŵ:�� e���f��m_V�x��:>dٸY�c��#e2�{���B���#����� +�N��r�C�*�Ba�5�;�W]tʳ��tQ|ޗvCI�(M'��B )J}<*0��(9��6��,�ړ�%�d�9\��+:�u�"9Im	����c�s"����(@�E�#�΋.�.�ĵ��2���-I5 \�⃷>�Z�eɼ�L��Z*�;��y�'��}���vIM�&hdП)���QJA�*4��"ɕ�����*�-D3~	s|L�	�6i]H����k*�{N�c쐇�2�j�xp�F�'$����Xx,�6,3�qI4�� �+Z���|���1�I��1E��$�q�B
L��?o%U�,��r��Đ����-9Ԝ��0YE��k:2������ֿ�y(���"X]Ȇ�
^����JiK�� ������NS���K�w��&���I������I���<V��
��א�m3h*4��O���Ԝ �b��=W�`m+6=zM��+�!�2�>����:C���Y�z^���k�!���f�X�:<��?��/��r�h�l*�(c$�k��!���6��(/`���.��N�28���M!�8�Xg��\u���z.�I�H������5�H��k�.JTì.T�],�o"�N!��a����h.�j5�'cT���O�FS�L������ۮ��P}�4B���fC	~�[0����Ǿ2�D�'�IV���f���~L�|;�$l�cX�:������p�~�^ƕ�%d������pB�t�m'r� �t	A_]�FTU�h�J�3z�92hfہ��C����-��O3�u�X��0��:0���4�\4ۃD�«�_��2��}<L΍�9/�y\*�RA��+0Fz�\�7������7W1�0wy�'�_#Q�	+��Ħ�ݚ�G��\~����v$�QJSV��UOfx�cĊ�;��ܱ�u�
�f������Y�h���T]�&T�����1�"�%F�\tJQ#m�K�>�[�;�(Թ�
�����	]1�$(F���T�p�y�ìj��k��� /V�/��%�-�k�����俽�<ge�a���p�0�䜅�6�T���G��#��綐_CV:FV�S	���%������.�9�»���A7ۖv��x&�X�k#�-����&��t�n��\G򻚱��eW��=�����+�����9�3��En�U���$��U���+�=��PùX/�q$;�����痒k|.!N��̰P���6�o���C��m�������_��`n��;(]>0�`�π���z4�Թw���ݢ�	�|�
���ju�?v�2=�����z.\cXb_�pz�0�}5+.E�~�S�N������o�X�W�g�Q��������A)�;�)[������H�nq� ���)QnbĿ�G�\]����nV=�:k�%�C Z=g�;n]r��_q������O�B��c[y�kw�B>/.��!(M-�<>����跕��}|ě��f%�;L��O�A�QBt�~%,arѐ9�C��a~ի�K_�D�P"M����]�rB��8Ҝ�lL������G����E�5z0��q�$ %),��	aC^�U7͏�� ���ν-L�Iy��?�^�F*RD�`HLs�γ�:�8!���5X2M �����ڈ Ղ�(�#i!�z_����T�;�1G�e.-ω�*�O�#�Ƈ���oIm0`c�B	l -@�U��{��r���&�b����H���^vKyCpp
T��Ai�	�I�v�I�6Q�ε�@�Xl�D$ 6�@ǉg��6A��}�I��<ࣙ�M��������$5K��(!j� �����2��h�Ɯ�ʁ��b����Q��9^pv�!1�����ޝ#{v��"Dc�jQ�N�-s����ٶ=�$��027�q*�4��.P��ֲ����~��\[t�VJ�G����N��U��Bp��(��$����Jz:pP0���3ī'z?�D�%|�I�UPyms ���|{w�� %�<����+�7-X+�ل���`�]��A�����V�l�����4xEq�L����\���-�0]Sѽ��%�C�r,g�N��`i�p�nSMe��1 �~����Z�%M�y����h�~0�T�ua�z�ji��d��!�]��]
�П#��4���LB�S��Q�[�����b��]T��#���ō��v��l���~A�$�؄Sj�:������d�9�S�Cc$�P vCa�b�n�����&�F0\���[q'H'Ӕ�5`q�fC�j��.�X�O�.#�I�;Y���ح�y��,BUߵ���2�,/���<�/V�B����wt�HJ��ӛ䂵�^(�Ts��:�
��.%\k��x˝D�o���#|�'��4Ӻp�/�; �H�l�C?�T����2O�+�$̀"�,*߰�"���-i��kB!��t����sY�̎J,��K:��鄱`�^ ���� 0��HW�<�Y�R�d`��~��`�e�_n/Z�L��2F����ʴ��,"ui�ſ��e�.�c	������p���dd�ke�a��+}W�Z6�f���E��/2!ڔ��3{��\�u��RM\NA���}�R&]tw����N,c5�"�orf�	��l���o�9��H�{q
hg�qT 2�#��i���jE��~)����C�O�"׬����d~��2��^�8(�(I�����Vp��08��f�2��M$�������ŉÖ�2+_�ny�����p�vSľ�O.*����J�gǣ�}��Qm��%����P��U��P�P�����Y܇/
����Tݠb2Nz0�K�p�
E΄�U���%a��[��L����s��C3��P9�lڭ��K-��0q1��y�8tK�~ K����pd7���KP#8'��Pؾ��\��c1�,��3�t
g��Yf_�>F�-��Ճ>�QL�$H8��p̺_�k��y$q�%��	���ܦ�y�t^q��E���g���%��^�,���Jd,��L%f�Q�+6,+@�#3M.D]��ah� �z9-�#���t��4{���H�a�'��lhYՊ��(�]#G��Jn+rњ��Đ)J�P{u��+���AFl�� =�Ea�ߦ�HJ�h����bќU��/�Y����h�(�����J6\�I������no������#e�EV���#��@��ޜ<n�a�;@�F��js�hݤQo���#�������k����<�� z����;PP���WX��i�/��~����iuɦ��6��Ď��������@��j����(�����L��5�5�5��D� 8.;<SD~�[q>�V���4f�n����	�w�I�`L��f��-�)#;�0=��k�/�b�m����LQ���)�v:lG���
j��_�͠U!��{�?��t�?f��>T��fdtD��.��ݞg���~�(������m1�D+@��(��<u/1�W���RE#��S�p���w�_)�`#�0DO�,��l`�/BA�\L��jV�ݧ��?.�)�u+�)�M�?)�e� �U�9G���Uv���kّ���V�ub�q!T�]�V�+Yo/�.�k(�.:V�Y�ˆ̳�n�{c�� ę�g6�e&��:"A�<vx��*P	�� 0~rif��_0�!O�ҷ/V����3�fZb�D?��>$����JE�/^cv�ˤ\��V�=�Ol��`�	��M&&��{���L�i��-�r��uv(�Йu'�/`5�~��b�?S>?��Ӥu!~�l�̳Ȏ9,x�~ϟE�T!ܡ��OY�N�6+2˹��%��>5g�?�
��7���Q��2q��׸�nC�S
���ȟ�֡kw��ț��3�0x�4/2>7���֦�?D�{פ.#�������5jp�T M�������5hN���aW4�J.7<�ƨ�,ۛ�f�0%P7v$�Y_VyV�����v/��e��N2Y�L0���U;��Ub����hSh7���'��ŋ��5@��	���6���>� p��s����J�r\zZ�5�.g�����B���=KK��/uq �Z��*���P�Sj�F�&dk��h�e"�Y̱�)t�L�+}�UI���4M�DjrKvo����L.st��vR�
�4D�.������tu詩2��Qۨ�jd���C�յL�gN�2-W@o�8$�K0wdE�Ee�!'
�\�JP�$�K	��+�Mͼ�b��Hd��f���Hv��U� �+��~+[�0�#�u�m,�BdT��_�mY�0�[���NM�7�
x�[�f�3��Y"���Y�O��C�4�^���J�I�i�҆��؋��Ͼ$4#���Ts�0q1ax}��\�g�Q8U�}O&�n��c8{��k
$��^��R��Fv3���ot�F�h��� 9H?�6B�k��~#ؚ;�)�15��;�T�M���^�D�wx�q8/}���n��"(w�%JS��9����*��<�ELF-�q�
�a\�`'^1��)��O��,D\FO�]I��k�\Y������DQ< �tK5D�D�f��S�1�y� �fʖI1�z�l@k�?V�#b�^8�&���;���ٿ���mN�n�Њ<��C�� Y��Y�-nw��y��Wq�o`����O6����:�(O���c�u�qx�A�:J���7bnN��ה��́/! ҙ:҆Z,WB�Eh��[���W��w���8 6e�0�Q`5oݘ�/���W�[h�ݲݽ+��h��������$�) Bχz����(�F��g�j�S[5�r��\������DO�]���O�X���'nY���ݷ-D�Vz�^OS�8ݞg_O�8��V9�,�U���쑖�@��ֺe�wb?w�f�y���i�I��	����U��BI�{U���X5	uΗ�|)�/��H�S�4�{F�n��H�=�����*u�hO�*3���5��yJ�`QC�
w��T��"yp��\��6�=�\��O�p=��I<~A�����<I;)��Lغ^�����9aO� a�F�	��S:V��K%GW�>XD�i�[�溍-�J;�����1��^�t���"/��fkE�R�V��z�2k����pL�Ca.xvƅa�5��Ź^	fX��&�XFW�H8�.ä��{��X�^�Z-�\WT�Oq�x¶�s����&5�{u@�x�[��y�������<��r!� �@v�9��/���	+L%�~�����й�B�R�/,25���F�%
c�~$�Ǽ[w�/��#���$��	��^_HQύ�b�l�\v�ڜP�_�#x�v��?2zv�u�i%8���؍2C�/ؤ�VQ��آu�|ױV��}e���׀���Wцtz,�W��@i!�M�A�v�F�TT>��'�UN4���A/��R8S/���~9(N�c�&�1�0L�D�1�����ڥJ���3 #c����h���0K����N|^>��� E�[la#�Vx��4�^Q<�����s&�zj(ˊ�^���
G��f���JU�ٝ��Qa2�.�/�����F����j��{M��צ�H-ߓ<A��	��6�a�P	pZZA��1��4�afg�����MoQm�Q	�j@V����#�]�������\B���k7�fp5��$�L�=7X�~
1p"�wE}/�b�P�Fڍ�!�����ԫ�"��p�.���bf���K�T��^��4���������a��%��t|��(����p��o�y��_4K�oo]ʫ�c�*O���s8�����?���l�L7f�[��Z$���ĺ6�"��x!Н���$��Z~W󋐘cߐa'&6"�cC[L�����k�;�d'C�K��E5� E�}a�63C��Dl�<=QR�ǿ��_Ae�]�G�͕RjzrZ�ߠG�K�s�v��ж��F.�Sz6�4^
>[�I��W|;u7��^a�mMG�J/0�J6��z��V��x癵 ��Բb��!b�#s���_'!r`~jX؂Vc6#�i��ddq�v��VדK���*v��	@�_DO���4����M�b�Q�P��vJ������� ��JL�� ,�>�]Ĝ7�k��=��-GԨ�S�c�����=�2���t���Q�F����LͶ㫽s�a.fy�O����1B^�Et�[PW�h<g�:���`6���Ij�d�D���c��ReO�� ��J~C�����8k���j�q�y�{x`���Y���{[�Z�r��*/:�X�H�ZS��%�}�i@ZT���c�l['ZP�~y_%y�
@+m-���f�aC�r���28|ʧ]�g΀�Z����s����g�<��[޴ĀK�_f�?��	��`�樾�&P�'�����
�Y��0o4*�%[�b��}i���}8���u0?����ϊ��+����3��F��.���>�]�ۨ�S�	8�Da��	QEM��ْ=Zh��r��E���|�L*`�;�w"�ipT���(�Ϝ�%���_�lG�p�ð�L����7����;M�T���d�5�1���O�9� ���u��3P��M���q�q(�a)�27w"pY{�Y8�|�N��J��iOs3eV��9P�t�9��M+ʒ��U�0gK,��ؐ�+J1J�Ӱ}�N���Y���Ü��H)������TeT��)G�� ,mE�`�V�T3}dQ�pS/�8�H��� w��^��>�r\u�����P"IE�#H}l3P�E���� ���F���7#q�q8̋��4� ���2�N�X��rm� �xd��Hdwy��R��Vp��C��^_����QaXK(F�oJ���bX���v��+~i���M^�H%�{����)>7�����1��[���yS�=I.#
�1<��h��Ԯa��yw/NZ��q�\��9͂��$�Y����-Z��&e�3~	����(��-V���9��9�Ź�\�l�YI��k�^�p�P�B鏩s���}E�9Z�
���f%���Q����@�~׫A4���1�vy�軓"�*�?��݉Բ)�*���'X��7*^���Sg>Nn��93��dWԪ��(���l���J�2
3�q2:*"pI�|��t���P�rTl�ra�AFW�UYLcm^7h
.��7�ͮ�>בb0,��P�	���ps`*�Eh���>�;Xa����uup$ ݽ��iÒHNvT�$�C��=E�fH��ޙ�k�?=�z���$����w��ư��v8kc����� �@��O�|GI�.��h�;���Զ�U	d�C��ƣ��a��u�ԅ���8�)Du9\�p�l����1$���u(�}����V��"XTt�,2T�]�ǲ��'zѸ�q?��Pc`���;���@K�.{1K�^���z�`Ĥj^�Ν� ����q:51�c�k;^���|�y�՞;Vq��ͥ�s�� �7�&����h�P���	٣>��RDz�6d[V�V�:�O/l��z-%����I �GS�M'�:&f_��s�Y@+;��9jum�<�~��U�e��i�X���5��UC���l,��i70��z�1���hI�L?�5&��)�xO1�Y�+p$�/c$E���k��먭_��i�&z{�2ӣ Gx'�����~,�'�K=H&�kț����Ny0���lj*P��S>C�8g��a�� �>-uj��P&-/�@�Mʽ� =���%Lz=W�{��72�����g��7#^��0N�Ҋ�d~z缐Yd`J�smVk� Z�^ f�Z)TB��^���7���g�4{����;(��$P!�ubΠ˒5������@���׃�������Y��V�PrsG����ҟϷUm#I'g-z� �:�4�5Pٗ4� #E�v $N:
�~�}�e�p���������<�~�O��c\"�O���P�y�7����!�4˙}VC���0d5+ᢘ��3z�=��v�* �Ec�ƧU�C*q�5	啬�����sfh�Bm
}��R�<�r�!�d�`;�!����9�3N�P �m�.^��&P,EC�[��
�-�c|V״w��������2�)H��b�dI"�7俕:��:^�p�N�1<;)�����P��h̎���8�GZ��C�@���.ݐ/iU��Ǌ?�|��4�w�p��ǲ�v �o_K���ӷCl�N��N͢>-T�n��v�8�ѤkԒH��'��O�>�d��)ff��%���Ξ>�~��s�I��6z>@���8>�&��M�R�PAw�?1�z�;N֘���ߵ�{"C�$��U�ʏ�`y�����F7��AňV���{��7�i��~�W�<�ב�+y��އt��F�\��)���'��.ӓ��iT�bh�&��gY݊�g��qw�v��*�4Vfq0�E�D�=�D;)�X���ȯ>�G;ZOQ�N�1=Jn��pd���E{��8{^�ǈ�󎪻̺�,{^��n��޻8��C�C~EF�WO���s���д��ڦ��m�C?��⫶? *��(l�H,C&�d0�2�F[�N�&�_ ��s���ʖ�b9ʓ�AH��>}C��x��'��( ;��H�ysN��
���mg�C�*���ŕn$s���6h����䔰s4����ZV󰅷+V�%h3K',���CRsW�Ұ�nMw��T-e!�F���n����&M��X(���'��Ǽc<Et�ك~fѢ���Uu^r�7�#W�r9���rw�HƾP[�����!�����W�hb���[=�4��A�7<uHV#n��X��O���r��.��wq��&�}��Lb�V=�tay�e����]IXg��׺�������.u駼��W�N�u�(jEs8K!��y�8�GK`�7z��Noe�IB��jD�|/�"��h/�rt;.��RQ9<�YM<e:C�#�D"D���M�+�i�6�C	���R,KbZ\`,�� �Ye!�&X��|�2	�YWB�YR�ko�o���/6 d�J{��t^G&գ�{G�7?����C��kG)�A���4� v�l��
O�4_O��8%���Rz������+5A�EM�
�I���{\�#̜Y/��h;��4pY
��q6������޾��Yڋ�i @�fe�!�X�e�)N��[�ƣ���M�ZLQ�.�n�o1F�Y7�巍?����N����=�}���0 (\��!_E�N���������Y� �*󸏊36ߝ
6��L�/���̷��9#���X^��������]y���~�<�@�s]X/������0�-����h�y�DE&|[���"�w68���g�'_\�z��Z�3U��m*�刾U�{��B�=l����QN��Uץ�����cC�C���2tV@�U���*�?�J�Z[/,��=�Qd�\�9c>�:0�����4֢P5ʋ� ;�+4��(uo��Pe�r2})��c��Ɯ(|ɏ����()B�;���t?��4J���(���1�������ԉ���'T�a�;|�mX�@8��FA*�����r̔/�lF�����f��.:��6�A>�Ӳ>���d~�:윎M���fC8�':�e�x%��0�b�z���ϱo,Y�z�����J��c8 �����gh��=0����b��Jo[�N���꟰2C���������oK��}I�	�-�땸'������� �u\Q%�*;{3�@�)��GT�T���Y:V�����y���ʵG��ߢd�:C�Y%�zӎ^>{\���t�r�t�V��<��?Az���$>	��E|b4�W
$P�V>_�[���J�JqB�E����!R�[�~W��f�CN���|4מС{}���%�;���}!�٪qߕ��.�D�iBD��kX�Y]�x�)�RQ����[U�l���U�3�r#}3���ap�A3�nGנ  ԗ-)r��?GU3�ΡR\,���J�3�-�jR�Ǐ#VDXS����D7�rwe���>1��ׯ�ޠc�q���P���_Bf��n��<�B�Oȣ�{+F��c��B41��ܻ���s���%��{4\ڦ����U�o"��/���/��gAssT�?�72y�EM^uǻ�c���y@�g�_�gC/��0�P��'�B��i��\>m��U�)�&
���.�� �jx &���Q��|�H�o������=��\	͐���R���YM*���/�"���n%�}��Y�B��Ͳ�:�i@��i�]�!v3i�6}ư�<��)#Vf��O�qB�Zk�a�ʅ�=z{���^Q��/T�֪�zc]��2e ~�~.]zq�nn�8t94�3!�`fK�x��!�Ex�꫌�CJ���V�@��<�
1�C3�*�7��l�X�-@I^	Uʭ:/�=�u_BOF̏j�ǳ��2���;� lj�z��m�S�|�����u�M����c��|���]A���D��ܪ.��R|�g�G^ay�ŠI�9IB��{�0��� /�����!��-j��*����W
j�-xް��̊�ۓn�m���7�W�#�� �E��
&S?�&�2��D�i�ժa:[֎QX�h��;�(�����PH��P�^��k�a�6�q�������㔉 :V�ݼkm:T%�9]�WmO�	�)|w6��률�	��r:�vO�c��S'?3,������=�����Iȳ9�J���b�P�J!���kl0���UB����[o�s8c��}��䇃k�}i�R�ф9��+�E��"�ט�=���4��]�`��Hd� �埐I�Y�=�c���ez�9ޙ+Yb��=��~�T=g�X)D�&��@��J*��&�[Jޤ�;�dm�u�Lj��;9*_���C҉�lg+�1�d�&�����N�Y5�E
��v��U!�`�w$��(x�XE�ą~@���XGI�Ԯ��_=��b�}��^R�e�/U!��v6!����fa&��ݡM�2K�ت��!�_>jK�PWI%�Fx���0�w��\Me�͋f@	k����?\��G�����OA��s_�W|x���w?�=.D���oKg�����k�h4����P3���*�����ޣ�q�Fvжg��EP��<�3��z
�=�nL�OWV�[Ɩ���-y��ٔWe��{)1���͗`���'�?i
ڱAw��5�G���z�㔼�1-��'	R���j�]��m�@�L�>��.���?���g�D�YV�7t�*jZFݨ8m�Q����7��$2�_t���r��vC��)����8��\��>N��Y�V�p!�l@�=lF֎�`U���묤���[�-��qƃ�]�y�'F���d���++	���;T"�HQ	xPmݸ�[�d�i44�8;~�������d�%0-T��}b�ĥ.��c�T�:���M�_*r�}��k�
N��*$��2F'������O��ÃJr��OC؍o_f<2�x�����==�����Hs��;�?�o��6��2��ϊ��Zd�Lҩ04�/רj _be�]2�/R�Ȁ�mw���/�+��x�f#��Y�	҆�z�Y2�B�X�DSW'�1¶R,��랃ĳ֝�s<i��%���lOm�������	��FO��12-�6�Q׿(4�Z��:^��N.�I(�y|&0�[9��������#�#��X�*o�m�����Ĕ���h���m�є+�H,�X�_9	*+C�����T�tXfi��1��,B���o���t=�y�����FQ	���ZxH7BGwQ)�m��㹫�d���~����L���2�q/J᳭Sd�C�)f�A�a|�>��@y��9;}�O���f���0l*��/�޵��H��B	Fy{xl�&��x��Q��:��ǐ��Ώ�ax�����Vn,�1�f��+��1u5I��:Q`���k����]B[�q(L�<�����G�rT�(�� Y�����Y��l@�ı6��Z�A�Lޟ˲_�T�zs��v�E5�v��8�"0����u
w厘�귍�`zx���2pC'+ҳv��E3#����$�%�l5RȺ�ӗ��,�'�'��	:�G���#�\MA �iŃ=8���^;u$��D���r4����rɍ�f���o)�W\<o�3�3qgMo�Ɋ���a��I^`�#�Ʋ��o'�#d6�)	s�qS���sf�_��d������ȧ�XD�N���`��i�������!	�]����ݣ�1�9��^I:1[GC'�9UK����W�C��w�����N��5y.^'�L`ɂt�x�y=���2i!��#��h|���|���0�Ng�7��jƸ�����;��.�rbj���w@�V����T�Do~ѹ6z3���Y
_�)k�0����䳋��������#4Jr�K�J֕���#��'�� ��-��<����a:�_��	��t�-�m���ȫ�B95��/-��z�ġ�RIǗ���5Ϥ�e߭#|�C��Ŏ+4��N��P�ĥIy�dc3����=�����9�v���L��Ed�Vo�!�Ѳx���Dc�[NӔ�>�3�/�x�n՟���������T����������v��cB|w�U�#�$Ӷ�0C��/J��ǈ��0���I�R5�i3�ͯJ���T���M�Pb_\���?4���a�^܏Lu~.�Yv��*�^g���rq���t�� �ч��	��P��֒�0�=�͹�^^����]WgS�sv7IJ��ЮE)����|�9��W�<�-�?�Q���J����Z����z��hꭉ]��h��FL�;n�IP�n=��}��7ŕM��ȍDO\���Ⱦ�"+�Id���J�
�S%�O�Lo�!��V�CJ�A~Q������2��)I�\EE��*3��N�C��s���>�O�J���b�%�I��C�8��N��=o¿�����ۡ�	����r�d��3[�BJ���mi��#43Y9$f�kh��)fh�>��O<=JѲ�-b�2*}�e�)@vGٓeT;���������ث��W�����Z{*��]��m��[_�pUUE�q#�F́+���q�U�a����}b I-�˳����ׂo.�s�"�!'�Gg�2(�����q-6��R�R+�8����[?��7��2��MHE��&7@*�"C�4��x��X�x<�:?߻��.�O��W����Y��ϫ+�:�|�8�l��?)�&�Щ O3�0�i����4��$�k}��=�m���_�=�`��L=�B����_���&t���q^��npAY��r�A�����u�k[6��XlmC��:���-�g�#� [���-ݠ��4��T����l���4��L�vX�ǡ�6�
C">
C�k�'�h��,(�%euJj*\qw��g:}]T��SU��d��� ��j���|#�	�9}�����[VY���>_������x���L�D�<ܫ`7���a�x*A�0g,P�e��(��_�F��S�4+&p�{]����#�o��!Z!�H��N9���͏�I���A�CP�g�C{@�D$��E�(=$�5�ވ���m/K�J�l~��dЀ��;A�6�S��H?����(g�~)��-���w�I�FM6-8����];Ű�5�p͔D��oq8``a9�'����:Y�c�������亏Կ"vg.�9� ��5x ���T)7�+���rpzs8d�gY0Y�����u6D��!	����!!��)�lW�"a龼����+�BY�%��D�`��9�66Cj l�O2��V&淭Y�����pc8!G����M�<�]����iX�{�i�Q���k]	8]I���=v���W{�
�,T��B��r�[_�c��jmч�d�kBe�4���^	.W�~w�6g3�a��F�,E	Jw텀0gOnD�I��$0��aK��߇�Bdљ� ��Z唦z�T^ߧ���8h+\s I�vC3�kj!�d���LW������ٹ�������z�����4�)�^'1�z�U0ȓlW�@�jZϻț�gm�QZ{�jhe�0�{�9��c�m;�mn��D�-�)WZY��O�=���w��.(��Y�h�&��w�I�^�r�Z����ϗ��_���n�?�Z	��[f�*y_��o��O�=��ӼыӴ��>6�hf
�5�j)�e���AV��e}�Sv��SX6{t�d������I��m������q;����7��{�ֳC�V�+@�B�>5y���/bƾB�]Q�,P��c���9��oY<k/&ix�g�_�Q�Y����ߚȝ�Sொe#B0l��x�e�X�7j�P����x���N�4O��0p�l�f�/�8%�����J8�� ��!l]���Ț������Nv���+Y����q�����'躝V�gyX+���"V��z��_�+���Z�.\��,1��r��Ul��;d�v�Ԟa�e��M?��&��)�&ASo��YC���h6o}�]�NE��JM�ũ�T�N�i�{k���� ��ޫ�_��;e�[������pؓ�+X���9�e�UKO�2nY�+{�:,f���O8@c�ʛ��Ԣc�k����`u��E��/���%��Nܶ����;Y �1�1�+�&�!In�����(��,w��]�k	����%_��N�۩G穁��抈j�k| .���h"�'gS�mog9Ų;��P�I�Xc����m��Ã���W��#wUe�Q�g���;m]�G-x�Q� No���,R�궢��Q��NY@o��Y�(���"I\Dr��/�u��u	xS�?�+j{���Q�F�,���޼�c�G^�δ=O�_��i�r���BQ��	eB�k=Z��?TZ]1�H�����O����ߣ��z�z�j9�<�����."wd�c����)����M]��  ���B����t�(:t�_ĕ&>������aQ�G[e�"���J׆��v�!�c��kI�(<�M�j�iڳ�1i9`R��i�Dq���<XPq,>ը�>FO��}&!2��p�߁[�A�׆�k��4#�� =g@އ:����L��9k&@�SSl�#�������
Zw����R�ד��8�Y��7� o޴�<d�M�SK�����^i��T����c�5�~��5�DX�P�6��i����1㑧�sV���Yơ1|�ƑI���j�>R�1#���w��n�4*I����?��ʱ}o}��C�Ø^�iΈc��<[�)�u�	Ϋ���zr��"�q����3@�x�$������>� ~4DX�px����%X�+������_a{�ɒ�l!���p�8�\�u���~$�t�me����ͻ?H�+x�l^:4N,gz�K����jF(��R�5��4�.���Q\��<Q����	T�e��� �F�s6`��-�:-�=�Zv7���-�������T���Z5o�!��b[�>��Z:_ST[��t��>����W����[�>4�D���T��g;%���!jZ�;�/q53n\u֞M�������k�K���ʎjU�
N%U����
h�EW�׻.N2��S��ܑ�Zic�m.�}��팳f�����+�h[���A=ɠV����7��qJ���?K�d�Q�׬�j>�m0ft��^��W�Rǉ���ZO���6Rq����`����
�����Vu�gu{ej�C�*�L��:W����Nyc��.�03�]�@���f��:N���Wet,�͝�dc�e{]����	�5AC�҇bă�ճ�,�(b �Yֳ�PWK�جN�NUf�y��@�w�
 �|��^j�����i��~�R�p:[Pu�i�ڿ�JV��@�!��I;���Uf���h>�Vj�=ХN��$>6�g:�W���T9� ��@��V��:(���aT�!������:^>�Y?�{v �L`��R����i�qK�� ?p�$"�1J��7'�t��X.G��m�j��Q�:���fu�7r3Q!�`�5?�Mx�/���K��P����w���
GI_��ɩL�� WJ[b������J��a�fF:_�����B�c��F�[�5� $=_��j�VƤr�/�I�r�;l�j4�Qkc�:�����:L�N�����Z���2J����*��4mា�V�s�X �Ql��N��G`Z�r��0)t*�pB�vc� �Mc�Z�/}�]�<������*(q�_j��E��g ��QT�TT�d!X�3��������2��_c�ζ���ⲁl�Q'�~P��&t��#놀zOշ)�S���Lc?Pz|&��ve	�7?!���;��b�0�ŉ|p�y��M�A�4T��}ɓ�[�;��]��`����½{]�Tgq"�����)~��UX���KJ��5�.��6�e]�L?-k�(�i�&��"��:Z=f����JG�+
����|�֥��*&z	��D�L�'��I?���H�4��ß3�@��*�u�;��Nn�H킡9��Ht��ѓ�E�0������m����������H�T<V��̂$�
�g�?��oY�"�̾��Jet��Xc_L��2��ߵ�n�О�:_�5�a7!�sL�;2vo���7R��6�yt�T�<�����zP�?@*m̶=��J��;��������TC/�ir�G�`�L����'�nfͱQ,H�2��@������Q��N�CU�:���;��~lCQ�T(�{nLЃc�U���1g���1��2���dx�db�M��KH�<��e*�H�c�0�=1E�X.W�M�fA�;Md��d�R0��8��P鵥9$:R��]�?�ǎ����?���f�6;Ʈܪ�z���veMn�~�n7\݁5�C���i����\
��M_� }���KM��{�P��.�(�F���py�����z��?���K<m��/O7��m8R<uר	������*DP�ꖯ�����������2�R��w�SwN��b��s0$F��(��M�5:d�SlQ�*���	����c������{`G����|���2����@�k�G�8_�X�o�A���H��"��E^T��oW�	��g�f���s�_�tN�c͙9�?����N������ը.c��7F뎀����Fmi�[�~������݂:n�j��2��:�����; /�+�0v��O����r`�VK�2�Yl�E]�=��/�ޔ�X��;�[���);���H`p���o˝4�i�Ŭ�c� s���<P�����-�Z�B~tڼ/��O�π��̴��YC����MO�f�=v]��iV�?A:�C�i�Qd���!� gP��7�*�4/��W��rC�iI�ħ�vOސ@���`��+�	l�vƎ�_
�i��X�0��l���qc�Lx%n��i\U.�9}�:�'B��ߕ�(�YVI;f��8���� 9�ٲ�/)�۷՜�0���: �t��);��PV����)EǭC�X��a�i���퉍q�[�r�P����?��0��a"s�Z)$s����~�Uk�������5�I��#aI���l��N�ř�60��H��Gh$�`��nA��Q8���>����e��U˿��VV�Ȓ���9��5R��1�+�J%��E�b��RIn)�x2�I�q�=��[&�ݸd���*����5CN�均�8@�i��83�.��"��-и�k�\[�J�����B�d�?v~�_���k��a�<�R�G�s.c�P �^a�+�e�$f���<�E.���C gǻ�3E��xo[�oc�OX�S�Aȅ^c��ѿ�D���i���'��z��ix#�𥸙OT��a9��_}�jEh�J�xJ��Vw������9[���pP'	�3іCIw��p*�E��D�,O��ф����In�Q�˜�/NCf?�
�5��=چ�;46�����܇�ʱ�	�s��w��!��Z�;z�Y5ڐ�ԟkU�-]~��9�5pr(�\�5��U���v�kZ�+Ff�$k��nBW��t�0nqY:F���t��9@V��ɂ)0&��!�������S�]C�3q3U�/�}TQݟ���Z���w�tϤ0�#��;᫄�����!���>���2k��ߗKT������PSαz�@[��D�L�r���@y���Azk8J3 �^�כ�"]�u�T��	�j>����Av����9���`��~��� ���5��:zH���ee�ċ����i��g��^����QmP�VLi�/�\$nO>(ɰ�12{������)`AVF7]�W�y��~��Н�c���[B�~@����l� <�E}��Q��&���s-�|��W��t��G+����GT�������"�^��Q��<*�a^��{.`��9
����R[��Ņ���?y�Ο�?�T�ባ˿}�}gV�w˳}�I�0�\[�|>���F�6�����V�_�b�m?�m0jkO�1�Q2�E��1��|� N�ѷ7�4���0�t�+L��A)t"��<��:�)�|�!��;�cy"y77Ljk	'� ����?������tRバ5��'����OټR�}�G͊h�M�o�N���=�Yu�����0j.�K]8s\9㊈e��@�l�D��/ro5���t8Fo�a���up.f,�Bh>��z�i�͊���� ^�:QC��Y�''35��q�h�X!�3/2#I����՘�%c�_j3%�<����~wt���J�S ��t�f�f�~v�$S���_�ק�x,���U��\&0�D�'�t��\\���ï�R-_�˝�� �	�RM&@���n�զD�h�p�6��yZ63��LAˇS��]h$�L�:#�К��Z��vߌ�M���k�|�Z/
|�Kȴ;�d n�x��	y�P�3K��xQo߻Ï3���}��)F�D0������������%�pQq|�f��x#�%� ś&: Hw�`�"����L�o����	�mSv�۫�����������֩���x����qs�K9�Ղ2���s���g��A��a�uP�V/�ʵ/Q���#x��'��*����[b<�"��½ȴ����uf;�v]� +�f��[n��%�1�3�tڨ;�zQݺg�m<Ћ(fpc9�]��ѣI��T�����'�˼�i?�e�YOM��oݍ����Up�����4��]�ۣ���*8�DJyh����m��_���Yip�G�9��X(KH��$G`�{��9�2�J�:�Ӽv��:-�0H��7�ɬ"rW��ߑ� Ck�����+��&[��U���2���0:���=����ܑh�~�+ښ���v�1�,�9���Z�"��]�}۟Gư�� E
�ۮɨ��(�I���;�������\�1��"��3�(8��u��+�4��k�@�2#`�|`@3���p�}C4�ϒG1=���Ivu��l_�;�2,��j[�����`��jԧ����{O���侈��������A��Ӛ�2
���E%��|�	�b�f�L��Oʿ������9�xR�n3�s	 �- �+M�!�Z6QjP=P���,lX��I	V�)���t�D�y>�'7�N�m�,�%�������\��A������ mME:�49T[W�b׫��T�ԭ��F띑τ���n�i�ܔ"�+U	ڙ��v:\����M8�Ɵ$>�fFn�ŕ����pSj���w�ǜo����jKw�7"�9ۿ�Z0�p�;�/dz=#L�<n����EXߤu�U� ����P���8F�F����)�q�Uć/>%m����o�b*��o��C�e�Q���)p��v2x/���jA�88��v�L�M\��Mr�(5��V8h{[
Y�By[C��{����R���pkCd�doZ��;�+��F2Q+c��	��g����|�--�����;��݊����A��U^f�6���Ht�Ba�#� 
��P�l�i
�NG���X�
� �,�f�����٭O� 6 �=�6.��M�����������<��8��730�'�;P�fY&$(CP��MߺG�vw���X��[�~�)W���%�
q��;����2���v�k����-�1c��m�������@���T�-*��M��І��{!:�k.7dM��4܀Vy��ﵒ��4=ڕ=�,.��i�ہGʻ�/G���9͹չ�7v.��#�}�����"&�_p�;�|�+P��?�Ƞ�GFc!��F�w-��� �	QTh�_g<)�P�S��S-1���=\:�1FtVn�YHs��J�k�U	�{F��i�-�[��.�TƠ�_c�N`V��v�"��!�N�?֮.���ej�>.iz�:�A�4��˹_tv�V�X�3��21���2���@7=na���;C��,�+}�ݵp�2�<��1L3�X�BF�9q��S�_R��~��3֒���Uxm�U��l'�u9��"�c��m= ��V1�<��]?��H#Q��q�HG��
����*����ίp ��R��f�0�,�)����Nw|����8F��S��dP��Dfr��z�����콓��->q��˩(�ɜ��(B�(J�O���
�Z.���ی�$��@��B���-"�88�{N7)g��q�`ɔ��Z-j�c��fY�ֳ)��8�c�؉���2��~�6�g�G�Ȋm�b��>'��A}w��V8"I *Y��D�-���^s���h�z{ڑ\�{�:���ۼʣ�b���1m <�^	����C��T!v���$�ׂ��4wt�ݗp/�	�\�MWA����XM�o[��H��x�/Q6�-8RO�"��	���XnP2�&W��;�V����������YHH�F�ŵ[�̯�^c�[nYz7��؀A���W!����˴����WS�8�f���0�ó=W�1U9aR�*~����Q�#�q���X����/*��w��B�6[qG,�]���mƱn�o8>�|7D̋�=E³8�Va�A*ف��f)���C氝ݎV�GZC��U2Ms[�/��?ſoh���Y��5�.�.`y�;tۂ�>�a.�\-�-B{�@#$"R̟�(�uJ�G��KMT贻��o&4��pz�
0}�-O��	����<�e�5K Ye��|�"Q1�=D�����n�s��_[7�9���𥗢6 P�& 3b�Wf%!H=T�F.�H��'"yhW�h
�vlC�HeK8A}+�eb%����@�	�-\�3w����j0���}8�O�ǝ�j���媤�=�3���8Q.W�f��b0G1��ů6����_ɞ�M����ķ��'�P��,ɷ�--�	�<�`r���\.��I; �$�C��^=�xJC��t�����#��
v[�<�9˩	* ��x�H ��3�n�@k���hh�	`K�敡�oU�����
�<b=������V���}%?�i�d]��uN��>3�s��v��5ķ�N��-�'Y4TJ���'�q��,��X5�պ����.�pi���������ep�����?�ě{A�,7"��1r�h��5��4�j�;BB{��J��q�x�곒yj<󧕅�Fv�u�xC��x�)BoP�=�;�z;szԮ�N�# ��sR̖�Pk���=��4$>�LxAMI��`���S�bb��E,��Z{�>��l�m�t����I���^p����S�+X00�j3��.�˵��/�D;8V�g��ky�a{$7��E2����pѱ�)��v����8"�R���ZO�#�~	��A(����p��F�.�����n���^�{�&�"����C�d�N� �<�=0B�ˢY(�y&��; �������P`ԒQL�L�V��(�B���E/��N�i� ̂���w����~��uM6ѫ�\�G$��P.@?����G�/��s$��B�ݬ/ց��&�cE�A�>�ޔ�����fh��x����/C�?�g�T#��;���Я;W�(�MP����U@�a\ �E�m?�LP:�L���/�����e���p����>Ֆ[���v�	A'w���&�:<�(�m'e���DJ�f��V�ۮ,�$V���dF0��p��Kӭ����'���a�/��ʥ��L�VY|a�)|`�'T�Q�� o���H�XGUp.��J������L+�%�B7���	���}cv��w�B�c�S�U���￪ `�j�߼��/�}3��qbj�  z@�R�Q����0�i� :Vd�'S����,��4��-}8����2UQ���Y[��A���C��)t �8QnD1���ʣ����,XW�5mr����JD3\j[t� ��E���
JR�4z9�,�N�k�Y�G������ژ$��}/޵6�Y��]�oq�2����x���H��A3E�5��U�:��ǯ��x뾊�غy�9�1���������LhY�y���P���;Z���n�8��Dː{4�����3���.ƣ��3�4G\�wHT����n���.���NH�b�Љ��n�xo���|�B~2㹺��ٰ�LRo���(���"�S��0b�7Z5�F�}���C�����p�?�􆫹�� �2b��bU��NA�<��yh�Ɩ����)j(����Ut�{s�V2TF�P])%	#v�g[����A��E��ѰQ
����!u#��c��I�����V�N{N6���*�Q�eϸ4�C)�>O>�҆�ص�Gn9f3L٧�]�^�������N��U�+̥*Hr���>O�?��E���i��וL���?t*�m��<��>L����U:��&�=�&H�vM�f��%�Z4���+c����f�(ON��h9Yӳ�F�����!�뢔�S�ƹ�k�#�5a`��}xY��Y�+w�y�%��C#R?�!���h��zs�8��~�h ��V~T�	;
��OFgQ�o7��+ji���0�����V���W%���(�K!����q��߷s:ה�l�f>Z�$I��n�*�C~�����T�;7���B�Ԝؾ�����l�ܭ�hZ���z=]�����Wka*@HDQ���.w\����sa����*�̑������[�UP
9��#l��G��}�x�E`�-9�;���RͯTHJ���s͞����j��������rxX�%�l S���*_�*�d�!��i�,O�0*�v/���]��"�mU��AW%�1�HO'��w��F4��gH�7�Ai��n���� /7��^����~E~ҩ<%'3�o p�΅϶..� ��Fv�V7��kѫMc�B}�n9����J����I~��
������_�݈� �W�_cE���Nݜ}�y��l�W������C����H���-��J&���71]����+?�F�9� )I���8����ڌn�ETxh\�΀}Q	]D$���ҡ �k��v9,0�{�c[�9Տ���kV%����;9c�=�Z���@p�ש�u�m���J�)3�J�/�<����Cj��U݈���a�_�&w:��uyA$��{Ӏ4�
��H�58&�+���p�'z��(J�B�Fj"'��Vk���6�/�Yi<L~+͂Yj��HXc����G?;Ҟ��?��#L�,b�'��䛣XD�{`�*:G��D"˚�h�U��`G����r���0�������(�Vɕ�k�A\%{�|Ԏf��tl�ǔ%�I,غ��G%��H2W��Ar�����f[um%cHf�p��Fz۔��5?�̱�gŚ�B���>'-;96k�\�C�B�ll#@z��[����M��p�2C�k�&{ku��V0�� }�#su)��{���B�E��k��q�j��"�{��R�|!�MI�qMg�/�dn�<�VG)P{�R�Y��V�T*1x��Q��@���Ht"���2!�����.C�c�����
k.X"�+�V����΋��,�RFu��u6b_r��B}?.ߐ��'�[�	+��`�=��9�֋�<�Ћ������r�X�K�����4f#߮�{kJ��ÛҜ�i	���YI�
������}��*c�ʿ�O�_{!k5"�\=F��.��=�ſ��$7 J�(��ыȁ�p5+_?����Y�n�JӚy�,��?���̈M��Ɓ�mbJ�:�hB�g��gFV����,�%L�#��c����I*S'�-5Q�8�]0���'䏭B��j^-ߓ�D�C�os���M�ؚ�-��W��%�b	��W9��P�ο^�Y[MbH��'85kb��?�~���|�k�����7}��{�Y��l�� 3�\�ȃ�yy�ڭ�<k���0�=IS�p���m�%��@W��5�a����3cC�Z���(i�Ѳh�Ҿ|���y�����\E��僉�Z��o-E��đ��W�|�rri��i�_1DI���j�m~����僒������ϒ�B+�*���,�t��x�[�Ml#� gD�Yk�U��̬E�H,���"iA5��>�U�%��:Y]����dJb�o4~�&����/J��a!E�+]��%���/<���l]�x�G�&�[��y���k��H�����)F5Rc�)C(�&q��R��WZ��!��f$���!�@I
9c�	bx�y�l��$>�_�1���K�?[�NM~�����fp�1��:? ��OW=������?hQ������C�y����m�{����c� �2 �\����X���JMF�L_T��SeE�I��H7��j��^I��f���V�}��� ���0�TA�'�yVi˷n'R� �Z������.�w�6*m����������M�������+��h`}/z?�`��T2�ޠOF���B�4�yO
aS�>+�9L��k�Dbδ��5�m�����2�U���V��(c���#�z�Cb$o^��^ى�!���GU�������4�붥Ѫܾn9s���\��m���Ų8� �J��|r6��p	��V��3���������Xڪ#��w��ؗ��	=��oW�����B����{p�5im�Nފ+��.UT��}(���ڮ�f��\h2�6Nj�u��-����kA��`eu� >�پ߭�ZQ�$sO��3��m �O�Ю=X�W�O��0�(*�Ž�Qs[�C�<�bh�ǫ�(.c}̟W�}&gA�d;|F�2"ّ�T ��
�rGC���P�Fʝ�ېM(��7�M���q.�.!�a�f����_ɢ�.��񍶮��Ib[��{Ĝ�e��A|���|t:O�
���E�nТ�oqFK��^)9�k����,��a��53�Ǒ�9:c�F �Q�q�
��{}�������Nq�X)n��"�����_��Ѵ��{��2-s(�>�U�s1[R�_�p�]'o�) ��ꢂTK޷�w��(���	(2��Zt\��M���'�Y�a~�D�B�����5�±�o��(�a�R�xI����ٯ�s�Q�4�C3��ܦ!�c���,^T��#]����u�R���tQ�L?�u��i�m��O(K���ԩB9;/��3~`Uo��,e�?��cY�yg͆@��+�N�Ud�&4h�\�Q�������:^��"&�d�ώ��CV�ԟ6pO�.�l�Py�^�d�9���~vfi E��($�~M��q��lN�~nRo�?�"��F�]��3��9�4�>ވü
��Y�Ux�vD&��w��N ����Xs��O��`�p�����:�ylҴM���H.y���t2k���z@ǻ����SӿKeE�Zn�a�(�/p���Ug�-:sIK&#�t�%� -���D��[��LQ?�!V��K玤4��Q��g�����4r��7O���>�6�O���Yno�K޺T{�H��v���}vC?Z���G��t4�UǏ��m3��~)��RW1��&�ZîGr!~S,����^�����F�4-0��͓uǰ��p�1�d(�>ױ�� X:�"��t�Z
��������.�}#$x�J0�������e�c^���ӓb�p����ABV!$-"�{���dz���b�SF)o�eYG�M2[ɣ��~�Q����Gie
�Эb��������TpS'�c��].�
�T2��s�<"`�
R߳���F��� ꚨ/���h��;��N����A:7�n�.�?�ˆ��{�J��$�c cH���CH��B�o_lIg�k
 �-UD��j���K�5;�|��c����ٗ��!`lQ��V�&�;KR�;��e#���OT8�.��R�%�IX{�1V�[>:�R��<�?��(���/�p_.��5�� ����r(�M\0�����!�L(?\�? )Ot�j�ݡ�]@Gy++����o~6��*j�{<�����]D�A�(�nx(��w)Sw@�_.r��O��뤟�'�*��h��C*>���������c�.)�ΩP�i�g�T�.�/o����/Ŭu�N�xH�qp�}e�nZ?$��I:6	x���qa�.�²�}�ը��(�).�!`���&��!O#�b�Q���.hm��$��V��N�κ,�(M���ݡ���@��/��^ͥ�(]-�}`���-�w3�E{+���=�d��嚰wq�_�.��-���o�ǈ1b��G�M�:���"r�C�Uc�0O��?�����Y�-��90�2(�&_w8�'�� |��Du!Ȭ��	�*P�Z����j����uͷ_�۟�г��*P�m��� )��7�UUw�,:�]����kO�����g��֪_$�s�0f�����wCf�)����8�֦;�����(�2�_pQc����!gZ�ʀ���:c�!��Mo�G$�Q�K"O�Jt#�<XI�;�)�>�:�$���+�9;���@��>}36��@��������$ çE^�����}6z�f��Y���O	vAK��j�	�V{��+�=��Js�Eof7��c}���9�!�=��.��GǊ]�nO�|��[�|\�����'�"�����d���G��Ɉ�2M^�G���+��/�-��Љ:�i���EzI}���o�h��������(x7H�뭤ՇI��^�cnuL] [C�ɕ��*rQ��A�|t���$8�\\!��!��2��/Zoo:�}*�M�����9�Y���x���]$�e��b��'�j��1N��÷�C屒E���[4��a����JR�s���f/@��KP�W�;�� ��*Ӎ-�x�@$�y'5�u�Kd���_��&T�
 D���]���w7��=�sX�������{�N(�ϔb���s���S0�Xq�#�YdOH��O2B�##;�3��O��S��	�B���l�R
V :�+�E�|�yY__ܠ�Yi��IQ���7�Zg�>!�Bu5�>跒4 ^Qno��3�d��N��K ��J�����������ɖ0�'����̾��������rD	�O��O�Q��Ȏ.�?�ȓ;	�]�&/W.&Q�-���=y�̗����tp��8�OI�@
�Qg�/[9��\��L% H�]/]���|Y�pA ����9I֍�V�X�����)��ҥE ��x�mU��+r]�1�",�ԓ��E�ͣ�_7��.�}*��&<��7o��8�w\( nl�� �z|�����hh��#�̭ɐ��MZ7��zF�A�֬��@>[㱨e\an��A�z�FX/f�鏖w��&���a���p�qf77�E����9�%�*c3��5�G�|%�tZ� ���ܱ����Qⷚ�#�"GlAd�Y�66�'k3���u���^�Lj�2`ah�
?�S���1A�����C�g(��c�����W���5����/?��{B�:�#]S[+T��bԯٺ9}d�yy�/�U�c�
�=��uM�(����u�e}�=���ڥ�.I�=���>rӤel!�-d�{1Y�N��zǰ#�ۇ�w�]D��./���2ti�Ϥ!Ck]�>wzjZ.�&o�Hm�X�n.�߱�|��)��
n!��!��u� n�*�^D���;-�oV!���_)�*��T�c3��O�ɉ�,��d��?h�6[�.h"�w�V}���*�i��|
ĭ6�;AoFo����.���ni� �ńfu����Â���@& $�%�O7N`��%�/�#@�
�_]��]\�
��0V)����}�i��,��V.l>� 9�~�����W�	*�݋V�L�0��z�0�|D	�hE/z� %��|	^ܸvȡ,��%�.���-��|~��,o�r}����7��zt�[�~����BQy$��Wud]��Q���d��)q�SVt�J��㷙��[�\�B���6ѧoԎ�t���[&[[ � ��=�ï��E巍"2���uE9)��w�� CZ���7uj���<j�JZ>��ă��j�ׅ���tFz~h��aL��˴qn��Z~k&@�bH:D݀x��Q��v7C>���;$���;-{�x�W4c�Xn��;��-������a-~M�I�JS���L�/�.r,��r�I�۠Φ�9�KeWAC�x����vGd>�u��R̙�oՋp�%��� �RX[>�zD�u�V�-�'�������[ Ɔ�]��^#}`0H��.d�}�ߨ��l�mJtz�T�nH�C��}!m`@N��sogs�[�DYe����؜w����r�:�gAp���"�K�o��s��aʝ���{�uu��˵�_�_�M4r���cѠI�5ZA��R3a
1ha�F��k�[�aj���	`I�j>t>ֿK�:�����ֺ�7K��(,��P��8���8Թ�����H�P�"��O�i�ϝ��4o�D7��� _��׶��7o�R;fJ �.�����lrI[>f����$��\� 	"i��K�j�;�P%�����`��g��������%l�>��g�tU4�t̬��J&M�;�w��u�pK(#�.$}<�%`���wԾc�����͗�����.`��;����H4D��boҝ�`��N���ƶ��Frm�,c��&����Ի˼?��F*{���n|M �|�m�(����]�K�l��>��l����ZI���!��zu�%[�������㩁MJ����PZ�z���'�m[��y�3�yY�f��b� ��Êݯ	8Ǫ��%M�����G���UA���&���-���S��qc�l:�1}��r��$�'�u�edsy�;A{��-��-����6�/�a/�\S[:�ˣ�[�ޟ�/���i�k7.O��� �o^�'r�;D�R�	����;�E�ϸ2�op�,��R(���\����	��9���{=��"�`+K#2N�~���;	N̙I���!��,fJ�*=i��ی�i��. ��S��.[���3�~�z�GOQ������4lj�`�?�|ҵ�+XHlv�Y��O�����cT����-����Ɯ�.�t��z^����y�Y�*�W���]�Nƻ"l�A�7C5V�V3���xIJ�ήRJ��_�`���T�/p ��|��jQ�	�����ӅK��Ū،ƆmIyI_Ix5.4�6�]A���8�"~��^y��XÜBd�,�i<�5�M֐$�r��t�S	�3��t�;�:�;�����N�R<*>s�3����h�� ٯ�
Fj��;��6���~�)��9�da�3�m�&��# ��-Qr��-�c�r�J�۸�4Y�5�]�Vo���t/���M�����)@ڻ1N�$}�MG�@a�v*ز���*nb;v���젝�jt"x�"��)��z�ם{
���#̢�U¥"���q��ɏ.���PX/��C{��w��G*b_�ӵ{��@aC�6�a
/w���a+E~�8D�Lv��1v�ԫv�'��R��#'�!%h�el<�Gba%�������\|ۈ\qY;�>�G�N�����6�Q��P}Y�i�������Y$K� d�=�B���K�zǏ�l�H+�'���u�A�6�Gd,}Ad��G9;&@�(��7)4�0��
1��T���S{��M�!�:J�u�ʹ�Ѳeڄ%�S���/\����A��2Íp�e�4Y�	����*h�&����"�|�~��k4@�>�[k�Ŭ}�zֹ����*m�����0�8e4Ӝ
^�K����$5�@�����;���-�}=��{ll����_O}�c^�JB�����b:���+&��̩D�ʧުr���p�a qIQ���Q=�~�ռ���3�����7��K����kX���
��xF��l�;{�_Q��Q���N(R���7�aYG7�o«����@��@#�3�DA��d]����;��
����Cs�ݰ�������������x�7�la���i�ƾ'��hqw$g��MC8��YZ�"��XMj���=��(��{+ �Ϳ�td2e�Ŷ�ߒ��x0�����{ѨUy��!�^�Ac��^v��?>no|���9�X\��-����U���(��:�P�*7���k��-�r��P~�V���b�$�]w���XE]�6�_�v_J>������u�(��P����w\�������J��捶�r��]�]Qp�w���"�;mw}s�E����A�wb`m +��F�t�A���qA��{KuY��v}�r��}D�/��t5F�(̩b��{��o\r�g���6<�ɤ��{8��)1Y�2�@���VԼX��׭�mX��듮��x��`��
g�A��qDJ)DUeY��q���D6@����DP09!�ݘg�Fbj⸹���¡�e��li%��������e��]Oϣ�pY.Ȥ�n涽��sb��뾽T���_讠����1���h�"z0��Z���ｃl�2�ͅ�7�:�E�P��a�h|����'�1R��A���i<���_A�!��J]��5;�r�3��:���0�Պdp�%�Zſ��w׷�ea�yv�_�3��hnIV�݂����[*�P�����M����R<�G����Ի�ߜ�}�r^���Ȧ�\�X\�]?���~�P��g��Vb�qAP<��ru߼~�(?&c�ζ��73�:8.>x� (*���@��&H��0�fn�=T�!
�O��%|~��u���>"�4[�-�}�2{`�|�� �o���m��M&͜+�%�j�  YTFC�J���~��5p9p�2�)콮U��1:_)T�;����N�8^��"Ih�$�|��n��T}�M��	R_��c��qC��h�I��mޙ��/',ܟ��+׫О3�#�S�Q��2�Ţ�+�ݭ�M��s���ߴd�/�=��:QZ�i)|����^����!��"K°��hF���f�A-�U�d�̙{V��P{�܉MJ�A����ެ1L�4	sT<�4賚�K]f����@e�X�h�5ǯ_{�H�x�ND�ʘ�Pi�A0I��!�����T�(��=�ϻ��d�!��*BLAM/m�e����FJ����S�+2��'Űu�L�qS�_4�i��� �4E5i��ʪ��i%9m��~EԈ�1�H:ʉ�-܌ϑ��&�(��QE�Z��unk0Y�W�<Q1���d��I�����$ '�_�wǇ���`�D����!;j�>V(Y��!{��@ĸEEҡ�?�O:x��o$W��@hh#?���
K7E��2[V���B����~� ��v�HB���\h?�Eԝg����S��N a�eY}y������ x�+,��,��M�YV w���T�L��_�Z��)���ؚ��� ����`��\m�,��C�Q� l��Ȣ�9+�~�����(���>ıM��I��"K��پa224������Э��7[ԳT�/�m�v(���r�"Lݓ��O�]�r'/���'M0}a����S� �����x}�?S��Pʕz@AϬ�� MB�&�mJ��+yTWT�$��_����~�4O678i�
���}�_)��uY�b�0o�$���FB���p�/EY/l����ІL�������d�����P�J�;EC�H�T��z �4��s.(W����D���b�O�=�M���<�(k���R�f�Sf��%�7 �ug��y�=Op��zp;�Y:�2�V�j��i��������m�c�x>�\:�C� H����KN_���xA�fr\Q�V�e���X��]���'A\O��n�&V��j\�#
"�����/�yNG��}E�1�ҷ-����Q2S�p�������K<��w:�J�~�r�����X*y�\��.���.v΋}l��iܗR���>
�#W�i�wo�_�mt�#ĵ-�.	���0*�
Mj�u��<G��{B5�����2�����:-sy�4�h�o��[z�ӹ�w"�\I�q49	�- !JBg_v�Z�&L�j�B�@5����N�� �>�r��~�l<����V�3����>X�h� �A�Uⶃ8�`�d��9�=O�x@Y7A�	��,x�X�R���z6ƪhK{��ǿ|�彞�-�-*�c��*�Nur��9��Hh/Oj���i�g�Ȕ99���
�o�!���ڸGbbٿEL�a��A{�����//�6M��q5 �E�s3e!Xzǘi4P`GS���x��ffN�Q���^U:#�.{-8��r��Љ��زu���u�U\&?��8D�3ϲ�S��~w����%ş:�C��Wm�\�8<�Y!��p9pH�����SA����J ��b���h���L��æݠN��N�G���Vf���xq��u73�"�S
���!��:�ʌ#J8��Ե�4ΌF�	?M�KZx�$5���{|Hz����W�W����p�!�E�"���2�YŚ�HSU?��R�/��:�YΗƫ`/�U�2�^�Þtj�^�PU���钦����ύ�U�4���툯��<�p�S� )b��5������jl^.�e�_���[�w�ϓ�HU�6VѾ����];�ᐘ$����(�ryt�o�]�V����X��`�yrr����dK_�ʮxtϖd��|X�W�z�ʏ,|�@�.�W�A�8�	��ut^�r�l<u»���<��r~3êò����$rCb��bݣ�,��SΛ��'H�@��l����������AU؂<{'p�=��[l��Bbm5�˴ǜ�2�Ro$������W�By3<�e炗6 ��l�62��?c��k�z�e����&�����_aQ5?iXW�U�,z��3�#�N
��l������i�su#����ok5;����@����ZV�	����-rI��p����e�a�&���06>W���PJI�\ ��2��R32+�S��{�ɹ�.�*���0��3L�f�%�� ȫ�x��[�չ�Λ�Jat�-���\�Ș%.�q6,��MǚD}��4�_� n�h��]A^.uB%�
�rH�Z�P�6�t$�$�x`:'��rὈ�-b�����W�����2@�9 ��6=@ULxo���5�������ߗ�Lg�ݭOm�bI
'V���)B.=g��+Q:��cK��e�GkL�_��ޕ�t/&k��)M� 5zs�=���R����~���(8���D���Qr�ݧ`�����z`��l�!g�%���:��=c��$E��.�<�C&��˙s�j��[ ��+ܸ����Y�V��nV�����`@E�)g�!Y�Д:�����ƍ�` �y�P2���
n�l�&�*=[�"h�c��K�C�
\����ry:_d#�7��S�3�e/��ɳ�eke�E��I�ۙ1�|��b+��h��*���$s��cW�(:&+�k��+z7q��rs�y=�*��צ������d�ztG�6,�7�.��D��C��"��޾��6/7��80B ����U͖��Ii�o�Mh�7h(�LUMϒ0g���ᅓT�q�)�?R��YPþ&� �9mV�7u���ȋ���kƭI{�*[@��Vi� ��ٶ�$vuv�J���^����T��U=�m`\���_7}�m)-�b�"�&L��;�It�p$���@��u[��Em�8���>I6��<T�AO�D̆�{�����Z�p�30&�G)��B7���k�!���;?�D�ΐ⧶)�N���*x#W�0s�
.�׌w�2�c�_.D�N����Ҷ)�7XEJ'���A����yd/6}�f��T�/�+�������Xx
��!�3��Щ;�t��]�!����!�E=^^��:��f�(��d��ƨ!D��rҾac����gE��A�[f��EF:�Q�1o����(��e�dQՖ�U�M���j����r	7��Q���+G���~Ӭ�^��5�F
�UCOr|��,�)c��~ptՃz��8�G�I�C���̦��ь0VwC_�]/��1{p�:��	#�U���a���A��F�6�;tT}� p�i*�Oe�5KQ�#��o���R�A���҅j�$�?י!gy����_�y�F�ľ{�\w�,zr�%K��ixZ���ABZ~]rjr<意5�XٽY�"�y��X���3K���U���п���5,+t�)��(x��D�|N�/�_� ��*lx���X��)�!oZz,���|��a-��j��7��"N�@"��]:�F��?�&[��9��?��A�>���V_�#c���@�I���W����G���m�������(D7O�*��S���j�+��;I�qֆκ��������[b���Gpg��IJ��8�����ָ�M����08�`��X��g���	W�Ҿ[�������4b�1�[J0�9W��s��\͊��5�HO���pE�Q,�	tZ��_��B}$k�$F�Yǉ�x�>�Yk�
�>W�%J�U\ǈ�K�?i#W�����J�$���-����������}x[�.\5T@�,�XيLY�J��muA��� ��L��M�����G��*������Q��E�FנE���Z`%��F]P��k@�1����;3�ˊ�ad�A.��~��f�s��5m[�uPa����x�,K���%-W�H��W�ƥ����A+hm�Ow�����d_"�1@�[���R���Q�[*:[>h�+4������?�=����h��7���x��� ��@!���o>,g3?���ȳ�M77�U�
&��� ����Ӛ���Ve$�ɿm�qϟ�zL
Z�����^W���'� &�!gFJ�G�=F�~њn���GU L+��ǢO/�ݻ�hA<��������ڬ�L�_Ӭ&� '��r@��s��3�&��1�����$,����RfR">����m��{�H�(��{a@����0L���;u�����q�Ћ̨�?"�7&�c���/���N����+�zLH����#��
��\��W;g�Ѽ鰅6��Ql,���{���D��y�v�-�e}������]���#�.���mJXw#]�5��[��Jo�`NeH(怙����.Zz[7$�Z�
l���+��eM�yt����.8l��Љ��f�1t����6��� w��M�K�
��w~�Ff΢489z5���S2�/�@���r6l�e�Y��ն�� ��t��K��g��:1�LD�O�?-J���p!B�`L�`�RK�;eF�:���d�D�hK����'���T�@$5[Uy=�~��z��=u��JZ���Գn��Ƭ|[������p~>鳗���l��=R��Հ���7�&s��`6�h�oxk������̶␑���B������@uq<���F<7���A�=k����y5V�|�fMi��"��*$r����Pu�}��St�}�`�p���ί�{��K�,����%,�!g���zYu\`�ԋ�Z?ò/֬�t�ѿ��-ʙ7�u��q	��*N"Ol\�N��J*Ȉ����XA��u�V�I+>�C���a�!4�j7�Fy���#}$�}�i�YL]����^}�)0zq��ij�Z��܅��[�s�7���⻼���C���{�C���'@�ȟ��`��rZ<lq�1C�ec�j��1�"�����@V���֥�	ʅB�*�d0�G�v�pg�[g��-'C����B�v[a5d�K�R���{Ίb��_��]"����e�1�����7�N/�7�m/^Gz���^�m�����mhbwU5�AG����-�Ij��I�+��M��T��kV\���0�ά�c6&���I���3[u��KiF���e]򟘭�3�^��=�U��vlli|���|�r�B�ު�ޢ�5���
e�E��s�v�}"�Á���&�d��n
{3a��*������07=�n�srq.Ie���8�=M/��9� �%�
i:�dr��nVOS�� |*&`^�@�ξ�r���g�;S{��ֈw?p��R;�[���n�L�Ğ⬌�V�<cs3�7��[?tE�@M������(\�
ٔ����<�)�B�r��c$�L|H��w���b��O)eh��/������@U[Q.p@���ɺ�e�༖���,����O�XV�A��|�K)� 6=]�Do�ʂb����B00�g�&(W��Π�GE��[�k+���W�����>��\4�h#��v�t.@�.r�h��}��P�l���`ڃ��=�K)������Jʠ�Gs�/�T��]�{`�Ef �ǰ��ρ���4;��+���ʺ��fx/��G�	�7c*�λ�n�eܕK}��(O��Hc���Ԧ��me�����3����\tZ*{�XO�X0���{񈓘��G�i��u�j3C4�p>iz9Xs�e�������Q�XQTê����\�^���쮐�4l��$FCϯG\��ܱ&g�i�#E%�>9��0���;�
8�vR�	x����J���x|����ۮ@�L�����hP8��y1���!92��;#_�2��7���Z��G����@HM������īc$L�3�����+~�^�y�5�HJ(�XAۊ,|��j�"��n��&�"^�kyqX���#�~�۶�aA;-C��:��Y.w�A���!|�~R���s�i&֠�Z#��x�^▖��˻���*8 A**����a9��uıՆ��W�^6|rҽO��wQ�jj�N�+�R:N_>��D�lU'Yzu��Xq������I��e�Kã1�[�o,��4� =7{�~1�M���HnD�A�u�2*ҋFAYt�	b ꟼ�j���(�4!=Ȣ����2c����d?=Y썭��b�l��n?w6"x��0bW�=�"��5調Zx 0��4�#b���k��#c��Ŋ��"��aϜ��a�!2h�w�zC�=k�T֪dy�����^����v3�� {�:+��E��2�;�1^[�����/˅��&�2AS�6��})�)[�X��5���^�ח���j�	%�Sl8�LQ�\�U�pd��-?F��Ur�F?3�D>����
�����;�v١�.��4�3��/!��5���F�2őp��޹���v��WN�1�o��Mps�"���ِ�U}p���}pN6�:�g_�]n�3�eŤ\��O��1�T���J�QK"�
v4�ED�Z�{��$&�ɶ����MҢP��qN���_U��O�cmSJ���?������0I�k}Í�v���A����8H,��>f;Z/���V!M�Vĥ�u �!E�S0Y٩�~�D+�הp� Ɉ�kzam��d�E���|~��������t�l�=4�Iu<�L�� 2|I(�H�8��K�{��~}_FU�Z,	C�\�����apX+`�3�Qy�l2�z��_zGj%��{�n�eטڎ�3%�3_d:b�w��W�s9�V�1ǖ.Yҍ�R�F�(�ٝ�Ƥ'f��>�s�E���7��AH����p�������uO���`0�"3qJ+qC�Ӥ��z>C����,���u]�z!\[�z�SAM�FV���>���˚��O�F����S��R�_lgHkq*��[��./�6-K�(�#��Y�\�T�t��y2ܥ�~���J��J��9v<�>3��T��q�?����4��0y��j����P{���1y���ė
�M(����[��%�I�B �O7<�<���ʝnm8J'�2�:V�=��QE-Ɂ�7�|�}X�t��p��*�B"ƕ��1應?kx��qR ��K�q
�=��5�wj	�W
�F�^�t^��ns��4Y߷H���&4P��� =Z#]��#c�X�?1q`��R��fw�������,/PB�d����Sbj����Y��}ֵDt	�t�C�fOt���'��3�#���̻v�QKb�����RJ#�=��0��J2*(�s2���'"X8���9�����z&��6���t��#`���de�D��Y���e����'�~~�] ���*��x:0
���>5ĲmM��(�>C���*��(4��?z���9P��Yp����������9I<��\I[�r��:I���Y� W�Im�q�P�/�������L��L����?��2����:���i��i�A�ɖuk�%�g���-o��';���ILCs�����$"?8
=��z�b���'W� �!Ksz^�3Y0���¢�&�
e���W�Ƚ��h��~���e�ڽ�Ai�M�5k���pS.%)ִD��΢7��'n��WtD�����#@��	���[�a��f޶�9@v6��.���z��R{�2\��)�-���^u��S�A:�z.�0�El�!>F�K�f��Gu�-;>k�$�]�fOMp����1��3���M���U8�p �<x��d�j懴_��Ƀ��T��/��8�ML�T���V�M����a��k�3���I��Q��7nfr̆�:��>��ţ�?r��$�V��o[���~K��n�&��ެ������S���ƬN$3���]?�V+�e����sJ��}���;U���2f�si˩��sDtapъɚ�����@�kYJv��N��&��Μ�>/����L
q�y�Q�8��y������A]W���	�j=`�F��H�vJaI~i���{0y�r�l�J�y%�����wkQ��^=B���nԫ�o�߂�-3, �O8[����5�ow^a�U8�aw����b���֌L+��sn�p���o�*���9e��j�RL���2���K~JV
P���+�r�)�������	
Z����/��x��RW�(�N�=�w2��
Rxk�Y[�*PK7�)�`E��@�\U���BJ����<qȰ:�$E���N �kHTF:�u	�d��bXʝM0F�1���UOu'�{��W�F^�nEJ�&�P�~�z@����ѓV��%��3�~�u %�eK��(K�W������ 2�.N��s�����
k1(�����5��9ʑ��|�.F��5��6Ѝ�>e'"��?`��i*p�d�2; �ك�oskg�򊓠FB֛AA��(_���UI����Ma�:ob��&��dj�"��lqK�|���������N�w�r9؝j�<�~L�2�g&''�{y�򕞗%�A'�������ꕑ�����:���H�ӫM���;i�&O#t/�T?�(����ujR-�gX��`�"�&PC��`/t������[A�;���h47I�m��'���Ɓ9�:%�S�N���|�zV!���7�E6.odT�P�$��zcgş��Os9d�Mˊ^�o~a�6,�|:��� ���$~�]*�W���:-�r'0G�"e���:
�΃J�����ƱMI��GխO5۹b	�r��i/(H�4�7��s�����ՑI���>���-ߙ�={<5dL�4s����,��W�F2��"=R�̟5��4R��>lxd]���=`-����`���[x����Z�J�x�`g&��z���� �V��h��tג���* =k��Բ^U止��׎9���/��h � g��y�'c�KDJR̓Y�*#��$�0p:��nC���a(�M2�H�)��av��JR�b߁7�x�7D����s*#�OZ4�;��Q�ںX~N�g���Q�з4��4ة���⋞c�4� =̻��z�X́�|��U�.J�D-��mX��+�(=}#R�ti�2�]�O*�z8<��7�:;e��Wݼ��/Ag;�?>
�0�]C��8�㐼h���ng��?�徭�e\��7B����B��Ɇ!�?`ͺ)y��j-�˓���~�[,���q�S��R�{��+!ʁ`�\C�t�_gh�u�ۆn\J�^)�\�������_r��rJg�f�,�Op<�
�?׀��Ei"�����3@�P�Cg��;+dn7k@���m�_�C��q|\zֿ7�e��%��xr���\u5�o���\T[�a�|J�a�!�(=8�|��3��2��Y�N Dr��ϩ�VQ:�s��秕�Kc���k@T�A���E��	=�H�M�2��@C�Ma)��~�*��f���킩�� 9�v�u�Qɡ�&j��͊��+�u�Q��$���R�>yz7t}A��z�)9�梣ԛ�h�
`�l}�^a���VՓ>��"i��z$ Y�,7E�_�W�V*�2�k�q̼ĦHzeY�ï����<� >k*���`4נ�A�^EG0����>����j�%�}Y��V��*M�_���b�K��s��C�-���O��~����g˪f~]����%�'���@`j���ٷ�u,U��4�7��-;.���Vi�ǩ���<�Z$ל�_O����k�ûg�#|�*�c�:0�z�qΒ*ƉS��7�X+K�(�Xro�Y����Këg4���#��WWR�sa�>�g������٠+A_1���.IqS9�E���}e`�xK�x&��2Y�Xbz_g9G�æ푎@h�A7}B���������lɄ�F����%½�����(�s��	C喇�G���&��UNp8X��'I�<�� {,��6`�%�o�B��4�L~�u�)P!��(�%\L����D�D�?>�ߡ!C{>�;��v�C����.I(�ݳ�w�CbT7?��\!�`�`��'S)��v���e�,?�-`������}�nK~�I	Χ�$ͬ��^z�t�V\N�"21c$�	|�2j�qr��2U�Σx�$�K��X!J+S�H>�@^Cc Ā"�jT!-��%�p�� G�@#��d!���1�b�a��[d�������Rǅm�QF���x����?e��G$KC�w�E��������I�E#�_�.�Ozb�){�D�g�+�;#�%�<W��;�Y4�f2�A�#|��wd[h&����zl�.?�����(},��Q��L��㞁����
���`��0f�?j�S|�h�9�5�?� \䢑I2!.�b<�\p�����>�^P�zD:��6tV�q?�,~��GIG��;�g��X��a�G���h;�P��K�}e�b�!��J(
�X1 �\Ty�K��5�7ۖ��2�?޺��U�����F��B�0Ҷz�;�H�~T���.� y�!N�h����4����P�{���J��e+_���`�OսsP�߇�\�Z��kh�E}�0L�uܖ�Y�������km��q�J�����wlX�� &�a0H��������S��S��<�`M~SJr;��.bj���*�÷Ĺ�
!�f��g] gu,�1-U�"���Al��ޝ��D]7���k���V��%c�-UW��_p�J�&w(�V�2��cR�Z8K��_���yX0�D���8�$��U������a�rA��#¹e�s�_�v����Ѐ=�"��_�l�ג�J�ب�E� ��������Ip=�+KЌ�� �^�Sds>�����Hl��pI6y�����O�7�����.+��C���K�ޭ��45Z;��24�a啟�2���_�&�^%�8h�H/7N~	e�F����S��'�
#��!.���XB�{/A/���F�\��V�)����\��[���POϦ� ���T�f�x��wm�x�S*A�te�_.�F>�R��M?2"����F�6ׄ��ɚ�&�N�1��lP����ӻ|+��E,��E�}-f\:���Q��y�!l��t+s����k�f��j�}&�c�q���"�u%���.�&i���dC��[a��]Sj�֠�C3ࢾ�T�~��jP^@�py{���At3�DT��D(��Ln��������~p8�1IPpe�C��C�����;6)�5���\��'!Y.<f�`�A%[�w�U�OdY����S-�b�a(ilD��?�5BŃ�lDw��owG}u�4�f>q��Y�	�&0�~����0�+\T���O�aX����u`G���I�=�C]�^.�Xe�N��v�]����&3CV	����q0�oz�Nz�.玜e�S8'E�`���̻�=Fz%u']<����������h��+�n"������Q�����������U���<.��%*F�\!��~���+��J3�z�lͫ7Q<2z��%G���Z[�w� ��`�w�������˵t��D��d�=�&��67Vˢ)^�y1]���T�?�/o���E[q�J3��Aδٟ8:��z��X�8�?�U@��VC$!�r�k��d��V��ȣ���ѓ�>������9Կ��˗�W��
U�F�M��'ɵ6��/f*�	*�¦C���~�+�>wU�ь���p���`t�����N��I7��|յGB񓺘���{W�WQ��nu�����~W�Ȣ�=�X�Ș�VE�����(� �����!�O����ϏF*2yt�)])3�4���!v�Uh�s�
N���Hֺ���	va"A=���z��0����q��b�o�o?>Z=���wōu�|"��|��];�G�h��2��.��z�5����A�\��}+'z�^�:��|̘��X��N�B�}���5=�fQϋRU&�z��s�h������1#y[-�~��á���i��ۻm����s�ޮR��X􅽐U3"jy�+{�C\�bI��o��K�F�fA~B$��`e�b1N�% ͦUt��'�4��Z_q�a��s~'^����6�
��+�!����E����ULU5�T�hw���ډ
QM�vj��o�|}��Vv% ���Q��_{\/@�M�VQ�=y��2m�9+%�]V��|���T�NЧ��M��	y���08����^�P}�q����e��"�����Ű!��}\��'��*�Y6}��W׷=�\h�9L��b@�H� ��S��ٹ.�憂��8I1[����|	�t���_�37�:����p)�N����ځ�{L���Cdϰn��f�;�t�b�3u.B����N('*?WUF��Ƕ���vqq�8i-��������g�?�j*��x��L�{�r/���ժ���-��7��԰5?�Iؕ�-���Q���h1T��SR�qMf�.;̪U�U�{�V���^���`����������<{�s��Q���L����)=����3�ξw���|��=/�?���T�/�yOLB���2��
�Tz�J�\��ݯ��YmV��o�8��12�\�4"�=:���D��P�X�^E���|�s�T�dPM(�[?YY����)�ȳ�5�DD3�ّ�~��_�����)��T����_���Ź�)f2&Bt�������\OFn%���&!�1;��FK{[Jv.��"l������	��V����_��?X�<��L=��]�=��Z�6��sG�^;8!��.���p�D\��hX�R���XXb�&�|?/��LqT���'ε/�T`��5��ٝ�s�Uާ��ȓ�&�܎#��B����nXB�Z���յ�"G�ߔ튓�� $�i�sK���	����
_,�dq�MT���mᅜ�1O\�qz}��Cg�����ƫS]PQ'"�X��ŀ3�pc��O�:%����A�@pir��	*�mWC#��Z���Jj���v�D2�p��(k�!��ui줓���R�ۂ&+�W>ԟ�R���Q2RQ=3������W�K&O���`��:s��d�^PO��;�V�����	0�{�s-��r��$;g�y�%�k����0;|�2���L���A��\��~ �����bj5f���7�"+Uy.y&� 42�?�����r��_u]<�R�"�n1���%�DK���C4'!M�+�l�^���ĺQ�Kl���m]j��f�P�Pa�,�q@^���tj��89C
���t�&7�o���.�_�Ѫ۫����\��K}���vE�+�_��TMR� e段Î
�h�GK�%ahm׮M]r�kc��%0�d<�H";����٭�&D��Ys:�>��ď����$�ǍՕJ�2 ]FCY��W=꽊����=-޻�P���"{�V^>n6�����|,�� e�Gn��Z &h?��r�G����N
?^$�&)��pRi�\��g����Z�U6E���T���Afn�\ȷS{�`�%q8ܸ,����������� ���-a[N����X�Ѭ�59lY{�{
�����"�"��%#�i )�b;o��ɧꧼ�V��_���
9í3�s��MN\��(; h���s��:,�)���;� R�d�Wy�+{>cR�Q��o�V���kT�Ve�
Eٲ��v��谇v�[��&'q3M9%v0�kp��4�Q���#����|.�k,~(Ec����W��c�O�U�/���7j���h����\^�q�=kI�h��lgbj̳h���&���0��x;j8i��hK`�d"��&�9��x螙�$D�8�SKU�)�Mw9�=�UXF���%sy@[���x��m�a�'e����>8�4mW�ܿ���é�`��:����m�B��j�i�
=.WL�my�˿�0g�s�g�{��^�\G*����R�	�������/���h���.<��-ȵ=#� �-�ٽ����>��xL���QM��}RM���q!^��ʏ���L�@�Є�=x`�9��0x�I �R��=Yߖf3I6a���둍̢�@k���2�07�yrI'�j��S�ڋԵ�.*�D��h�<����l������o��e2�����N6)��h�ya��y�E��c	�?������Xax���-�AD�JD>����:�6J������n�F��q�[��׋�я�����/V�9��e;�lp/��03�$��X�~:Z.*[I�_8�&�}oAL)X� ������?�ઋ^�-��n[�^=R���[ɚP�v�2xH�C��_*��n�_˿�~��^�B��UC7� �X�-�0a`�M/ڟLi�+���Ƭ�����./NqO����L�T7�A������|�%��X�E�q࿥3�]'���(�ˮgD�������~�u��4Z���^�N������֩�B��p^�0�!����߁8�	}��^aye� �Z��d1��r'>$��Ad�ո܌I.��6G�G"�^����S�R�,2w���nL� ���߼]��mS KB^�!����2B�达��I��;@
U�J��|��]|����LGEO����WK���%�XO`m��3'+��Rr<��d!��#]��=����]ɂׂ��#��S+��(���d�wߢb�����>2	����<z22	�_���PH˾}agH@B�xpVH|�!�����Y�{TZ.�;�8Sڦ����f��2��z�7�ͅ��c8���f9X��m8�/�Pt�����f�Sk���)�wQ(.�za�����Y�w?	�0��x��)�Rü�1��W=�E�/)�MsE�L�Q���5�~���[x׫���7:��'h���G�\�O�PYW D��eT	w4�s�kT���@�vV����ߣCd�[��^C�׾3	oW�/�s�