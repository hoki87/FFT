��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n��� �x�vqΕ�8�_��x�0]�
s!N��(��pc�(�},#> E����%�X3C�5_p|���FU�1���o��F2��e�?����`�Q�\� ��Au�U��5N���/��5�q���x���jy�{˽���#������-�r ~HP�u��D(����N �~	�W�����Ԅ��:;��A�HE��/_qq:�bJ]22�������fqh�a��&O�5����B��@m��t�m}�m�#�4,<q5�l�����q�T��q����'0C.}-8=Z[�x�7�S�d�"��H��|7>^����P�u��9.�V�C;cV�:�A�N�
%��Nz�}�)X�:�(��+{2/>�p�7�v���Ə�o��pȠ,�@ف�����B��C�k�b�ߡ�m�Y�Q��7���6�n�쎂�ڽ�!�GAw�[�3)��+�0��Q�f<�uV�t��9L�N�iQ�g�[S^���8��[j90�����F� צ���������./���+����I�E�TF��)Y��/F�k��|��y�����
�`��d���4»%�/9�	B�\�p���du��<��7y@��qVn�һ�������?WJ_�����Jwݍ���L7���B��M�i� � �VT>�<����h�ܦ�4.���V�]�\	���(];��{�l���t�pCŠ�.���y�p��F�=�D��E���;p���g#�T�m��l,2�ό�l��g3w�Ԏ�,z(����A�����ya7�[Di��d�|��[f�-�Ivɺ�X�x����Y�I��.ʖ�R������	�믅u�P����~�� �S�]�u����4��TKl�D�[C����u!���^ao���1��Vyz�%��聣�΍x�+z�G�!CRK�z��LwC�{̈ �T��cl=�~���)hx��3r��r�2~*��� �N뀩��t��ἿQ���ɾb4��x�;���9~sA�ր�u�FΩ�m3	"�*O�ch6����[�V�㋜��!c��K����A�(0�f��A�IΠB�Pؿ�
w���LݭPt!���� ��4����\�U��[u�R@޴�ޤ�i}��4L�$t�Lr���ߞ�!#P<fĴ� �$�#E�R��.z$5��U�^��t�!��3聺RT\��y؋� �7|�9�!u��ֿ����;��!�!]ĝ�}�&RW@9b �`��P�U���`��}�\A�Л��ڗɪO�F�X�%�!h�q�w�_Q�*�:y	FЫ��%T��;*upu�7�5T~�=�i���.�$t7L`J��CLt��^F»�m\�,��C|�PuL�m����]��
�5T�z�>��-�ƣ���wtm�8e��Ԡ��p���s��{IO��[��u�Gd�.q&e��ɠg>�u�RI��4�������
�P`H�,�7�__��²Ѯ$ǍC����Z���ae\�~��gxe��-f�گ�`wy2��c%����da���Z��A�ł�T����t	�H:1$�D��2?��h��*�{\���=)�|$	U s�a�i �~����|>���c�^05��N����G 	�!E{��30	'��
74� [pw���'���U\�ɗ��}2�^X�~����4����&w4!DT6~)t����﬐�C��C�O��ժ��$|'S;vZ�KȘ��ڂ�i���h�&��V���~��u�n3h��wn wb]0AO�Z��::��)��8�!�7�A�=E��*� 	V�3t�m�6{m0�>��TLk���\'����>�H����*/�^�*{D�v� ��^_�W�[(�m"�TWƊ_�.����p3�9zA���ޣ��ރ#�����S_r�BA�vZ2m߲c�!�&�  6|�'ҵ�Kr} X���=�@��S���w��6[�ۯ_���Hf�b���j�����R�/ӽ̔��o$��G��K�7J�T+���8c��D��5���Jx� ��D�5��G�WyT�����Fn���0�W�I�i������b��ILH��#���E,�N�u�-��p$��"�����bmt�:���
ħ������e�4>��H��OE�9m��bp���M�hF�g@�Y�Om�j�I`&�a���b;�+��gdQԾ�WVi_ >ۧߓ<�^.C:1���%5X���N�g�2.D4*侌=l�{&�g�*\7��-�/l�>�po*!�BLz�
�K����ڶ�����̊B��K�FT���Xl�[��7�i��%��Qw��W��$[��*�q�_I=����.W[τ'ɣ
12��ٹ� R�*���1'�$��1��j�}/㬬�Z?V%�5�3�~Bx�r&��t��L6��~5U:�pu8��\J���e�)4K��$���ĵ��	s�x|��QK4�.{s���b̔V����'�s�HLL)5���U�ϑ��1aʰL�.��\q<�]�G�U�����D����TL/δ���(I�"q��<3*���P%�b��^8��N�cQK~N�Ulm� C�G�j(0v!�[��,A(�{�7�f %�QE�YUk�o��-���B٨ܿ+Ƒ^��9��p!KD9����_�&7/�3W�D ��0;���۔���	0#�Z��Q:Z>�0�%��M��t	9��1o92��f�exA)��{�$�Q�Ze��̄�^��[�D���&�Qb#Qe�'"������r�1[S����!��?9� <N���AS��+�����0A�`���ʏ���HΧ#�y���1�o#+�[�D�1��N�,uX�Ӽ[$���K_ބ�^�8����a�+�@�6��4xq-]Ԃr�*���C]LQE����p q�Ą
�F����$C(z^�,m�:#���K��6�ꭦ7���� ��=�(��=v]���S����� ɡ���;�Ej��w�l�5H�K�� 3t��nn"�YF~�YY?`u�$A�
�S ��t~aH��eN`;$֕��`��+�ȼu�<Ґ1j��Ps`��EI� ��?���a�'���1>��*���Y'h}r�vTe?�=�?o��)��ȴ��L] :ϰ>��	}2>Ț�u�q,�蚴�W�Q�|ǣ�jZ�[CW�`��c3o&��# #�6*-��s%�(�vx�=�m,>�Wd6�Dl���̧��5@�+L?Y�:g�^����WEdu�tKj��x���e�|,�L|�����*�h�sJ&�,�n�*�V���B
�	�������G��8��ox���ڿ�w*ǒln���>;�Ȕl�^)}�X&�ݽ�VP��D�k�5It�u	����D���\�G�[�IiW��W� �>��6�;���^�<$���LŢ�U,
�=�p_V"���`���=�Q��hV���(�C|�t��y7|9>%
 �bYL�����KK���䕶��z+��7�*��1�dC0C7��V��o9�&dC����
�m�ô{�R?������o~��w�V����F^���Ա�L���8�0 د]���oA���.�N:檒0�K�rr��"���G\��$UC[����})C^n[E?>L�3��C���q�Z�%2���b�hMkI�"�F��C��j����l3�+�m̛)	tsk/��o�,ta1�k���Jo��}�,�7�1�Ǘ�[Q���DU��f�6׸2���\*]��4�N��yZ��VK�$[�2��7���[êx��S������Rܯ��N�3
������3�k��N�����9X%��g�&��������P�?>h��i��z08Fo��>ϰ�����ӫ���a�vh���ph0`�Y�;���j�{GLŎX	��?�1��<Q'�nJ��@=W���uN�[�C�aJ:��p]�����HI/pjK����2�G`�jw���?˕��6o�Mu��yѼF7��Λ�r��o{+�I�"1��z�VϨ�2�u��~�7�'c(#�o !Z)*/�B��~�!��Cv��FrX��y��� 6��Ra�4�#�ѵ2��0�6)9�Z|8��m�x��v.Y|�2��P/AozfOV^I�3���`����x�9e��<�Pe�gߝ�y� ��<���z���"y�E`�ӽ��L@z}@�?-,��Ar��*�ў!"���T��O�J�[��@�TN�#1�$xJ�x3�~�,�;)�d/v9�#���]�Z3�V����6L�b�ʐd�t�-�
�r�u;f���ق�����g�!U�;�Qġ���A�U;���	D|׋J!�1�=p���X��*���.eR�|�ᜩ��ój�~`q�׌��=��ǷE���
y_��9��מ�}uwST���:��J��B=�)��¿�����ćs��Y�^��{��	ez�h2��A L�Ht���f�S�u�:��b�R��?�a�F�:�3R]J����_Z�C�/�ǇK[Sp8�g+?�v'p~-�{m�06�F~L�:\"�-�
$��e&v[�)��~���BT�)R�v6���FG��k6�,�\���W�A9� ,Y��������ђ�ײ�?�7
���g��~��:
�im -+J�W��4��)=���� UX���lY�pWb��h���[��4�(�,�_����;+�ޯgv<t$ �j=�/}�W+��p�
��`w���6:*����Ys�P��X~]K�5����B���_��x(v��z��E���k�����q-���"� ��^�z}bsB�nؒ��#�vg�?��Ư�~ш��ali:~�52kV[q4�z�\��t��e��,�A��9���M]���I��ɰ���x���^�����+�;fH�L�.}JQpA�m]�V�
�c�+�W�y�a��7���5����oF�����\�K����(O��蜗;��>��V������x��l�r?�l_�i,�ۄ.�Ƅ���U_��M�]�筷!���E Ӥ����m*�V
�����R#D�%^=gN|�*xs39�5�o��;�F�jj�`��ՀV�-ם?����
ڽ[�c����!M	hՅ���<F;��Hy%WGA�	�����6_��[gp��7��fpm�)����v<c�>6^���a�Qf��>�Q~�@���n(~2ʴw;�p#�z�!߭�l�y��(1��E"��w��g��������g� ��?����	V�WJ.�<�8^Ϫ����Q�
[c�2��>3>��g����T�66��-��`�J%�#�&(��ύ�Ƭ�ؠ,#�(���{Q7c��(�����*��R� g-��q�q�\�J�5�� �m�eGn9Y ��t�wj��:��pH��J���f�&��':j�W�;�N|�b����q�y��+�w��W�8���r��MT�%��頹�ێwl�i���J�?O���M���i
j��w���׾p_�-A��]p��Ť�q9�<;�Kk�5�%�b1\�OL���7_D�l˹k��bn��'p��K�|�X+���4�V�v�EO�9���F"��w��u3�ߙ�k�I����B��Tb��;~|��B��̨B¡���#
�|���i�l�����3�i�܎�̄�<R~s	�H�w0��-���0�ƹ�����LV�6Q�;��[����W�o͊/ܾxC��lx����^񭿐ź�K>��%�)���m*XhP���G��Bd�r����V��d��*z�F1֑&d�t�cWa��&�z�b�CH�^۝�+�O�))�ѥ>X���jD��xO��W��!�˽Hm(
4�i�S�]e�N��g��ە	E���}���uM�#�>�!1e>g��;ZY��L2�@�6�u�Ղv7���>��Ɯ�2zy���⛝N��P��Z������q�X/qo����tV�[��o"T�����;x劘��k��Aη�a�1 �G�p�pO��#u��>�ӿU��H�^�r��s{�X�n@�oT��/�)�Ϙ*f���E���e���c��=��Gq���0����3GQ�C�z��vp�sV�6Io�_k�����̆ȤQLSѭ�G�{}؇��T:��.fe �?��׃jyu#=I�f��x����֚@����,;����҈��)���3������`��όG�I睢��W̮�e�}٘�*_���~tԧ6��ޓ�����l�s��xӚ��%�;G����O�n�z��yM��A���%��e��"y^������$`�m|db�'�0c���>`�`����B�	����??��%D��R�4�luȩ� `�CC_�]xy>������;�(/�n�^�`�&%�{I��~�8L��G��o��<P�����/lὸ��6|L �}�ӊ;W���@pI�&x7.���o�����Mɦ���W��f�z]��
dC���7T�AR�D���wcs!�3ʣ��3�V�'�7[��i:�Er`f�3�t����IEN:�2�H;r۞�*�^y*&c7�z;��ߖx
/�����l�w��v�"����-�	��Ć���7YP�����rԢ��ղlx=��1w����q°�eK�D���"9��sB�7C\	}�sia4�����f_��m
�ǡ�J��#m0Y�7�Ƣ,���¹m�%�<N������WC�k;�܄5�<^�"� N`[L%;|�DU!\*Ƭo��p��@8+L1�
�@�m2�S����������s,�#������� ����#,&w�c.��fç�oL\cČ��äP��J`�0)?��ݤ.����>c����Lӣ���mD׼݅�|I�o���o(A :�c�m�g��/_��
�D���ӧ����ϴaȪPUX(/���i�F�v��R����0��J2�۝y��dM旖��0��n�i{�>�4M7�+�#оL)�]��O�,핼�#�٨W(:M�� � �yׯD@���-7�K�ƿ'/�Ge�ɚ_�����v�1_^IU��b��=(��Hh�B�0W�*�.x_���G��tEq��Y�SR��R$��#�?f9^@x@hB�0T,"�M��GH?�n;��� z�x�a>�x�R��I �͑o-~R�v���\���GX𦅮]�ڜ*{�?����n-��[�(�@�ADxE:���S��@F��NI�"TU� O�1K����$��w�����g)�>�M�+ȶ�ϪA�	(�v,xyA����;��N^���o�s�y��b�1_�Y���`p����Q��TG�V���u�,v���v��R���]�����,����}�ƶG��WpfA6iM�T&��=�V59�A�G&����r�~���o��T3���F��pg ��r0?��<z���C��ѷ�� y^��8��:W�� �u����CR�w �u���m�LnR�'���F(��@�|8��;)���3W���t"G��8Z,mcA�v���7�\Y9Ū�\,����jZEKDݣ�6��	����gP�l����~�(����(�i�I	"}DٔąZ���^��wHW�J���W��'cV����ME'��N]W�P�]�֋M�6&��c����P�yx��\dYr��{k��ȃU�"n�@�?Ux ~�e����>���s�.����S�M�[�[ş&4A$7�?��Ċ�0�9��y�%��]���:U���!,eNB�;�%������cȪ$27S#Q�72�О�]3�����I����dCa�r]޳�x�
a4wT4�cІ�{H�����Ǭ��k6�� ����7v�\�ٌ�`�ݘ���a�F�s���b5}P�3L�����2����.� ƌظ���jW-�'�d��ica��`�@7	t�ƨ�`�XqQ��=���,f�GzV���r`��1q��9J��SA����&�G�r?:Ê�����V�u{�1�/.���� E3�M�-#ć��\K�	VnUW��ՙM2�eo#@�������>Ξ��c�Ou{6j:)����-���R����n~ �����ml"���ۇ�?�U�Tڄ3\SW<����A����M�a�J:�@�J��t?�!���	R�fߺ^�,Q-�z�E�s9];�O��5���0PҤ^��?R+��C�*�P���Raׯȴ<�6�{P��-��<��>�5֦;TSy����J}��d�Q�j�I��P&Ω�@�Dyy Ě3�1�/Ű�2�=��'L �CZ:����y��*B��t�9I���T5��UJ@PU#�