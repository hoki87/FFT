��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�#&��#�<�����{�sGq�*MO,.���buD�"���`aő<��<XB�:K�z�9�e~l�9L0n�;��a��$F���8{�u_٬DWdZ�X��2`C��o>r�,��<oU�3Mx���C.X�,o���#2�`Z���}JYf�6�J���_~��J�%��{��!�vr[�=��Fd�k��9s�|�M6�V!`��3�}��6aN�ݤ����sp^�k����|�Bw�^�桕�m��"���$�gܥݼj�a���7J�F to��U/� hKt� _[^�^;P�6�RP�|+�����}���+�WYB�C뫩�o$PW�}Z�l3�ibں���;���4��ݶD���ϐ�[��/��Г,��;����H�8z���;;݉�W����ѯ�I��v��vOB�������$��W�e�0�A�,T�Z�[@�T�ث�������a�� Q#�{�Y����Y�����;���W�����iX�c��ѓ��Hu9R�.��s��G�uQc���z���a��ώ���
lw'<\�>��(�@_W�q�ʉu�&��C�.?}�}�'�4�"E�\�2Ì^h�+�oe��rw�w��S|#N�;,�Nk��Q��Wv�P6 �2 <�`yY��4�ɈV��f�"����x@�z�W>�R;3ԛ25�Rd���da���Y����S�>҇rWd�&��0�e������S��#j��:_�d�tlI�L#{D�"���Sq���d�8u�դ.�[�}fK��F�o*��%��QvR_���<��z�����4mt*��}����< ��������G�w��D5���S���B��׸�gW����̙��N1a�n~Q{���G�
&:�N'�G?���"$���bbo�R�Js�wX+f�c�����i�=!�Y��h�N��JI̸�߲�\��?�B����M���L���)޶��]�_{�K��d��U8Q��\Se�$�) v8-=s���˙B� g��i�x�3)6�n�~�Ԯ%J�^m�#2Ƈ@F�80�L�t��NV1���)�S� Z~����4�u5VZe7�:&s%�	Z��Y�6���{�;6��Y_՞@%������ n�D�SW\dy�c,�>��I�Ju1It��
	�O�,#H0$�8Wl28�'S{b
m#�ڣvm3C��6�u�\#�:��Y��x���`�v��5���� c��#��`.�ZU6�� ��q��89������F_���^�,�Z�j�g��`�/��i���h�a0f6�8���v%z�j^�gI.������N���K�x|7�!��8�O��8"9�!�/�!TG ��k�yÐ�2������6����{��La��y2��ʲPQ�g�_��zci�ϐ�W�R��̂�<i`j��'�DEJ�b�] �S�ujּݦ�u�T<{D��0Z��_L*o;���D~�}�n��~>��n���Rͺl9�a�1��Y/�UpwP�3Z�׊�z�H��
(�H��"&A���A�oKQB<�z�2 �yw�����W���m�W\A�����(%��f�9�F��GV8�(�k{j��TW�АF.��)����)8�;UT8��Lİ��-}�^���jT�n���2�;daG�BD�Z<��L@	���x&oK��6�8�O��a,꥽��F�X?lø�O>��`z�%t��`"�!��(�J�Fn�ܠ�}�W�M5�#F�6��i�	���1ְ)�}w@P�����#���k�e��k]��P�� !^W���[E�9J]����K��ę.�[=[���mu�FU�U�	���Qt5��6���@%��~��D���5},n�o�L_c�������H=�=������s��g?_�7���b� (h\Ks��pt�܋1C��$O�(�3���yԹOm�Ml�p��["�aY8�d�0b��!��+$7�[��QO�Ğd=Gn�[�)��
Rx���-e�Z�Ʒ��ߒ��TɦW��=�e�pJgJ����أMR�QH��Ԡj@��*u�(_#")�Xh�%�h���E��)b�ix��Xe9�����hnEo��񚩋P{��,����#_��A���b�"N����7o�+q֛�88{� W��B�j~E	yq_���=�{u?��a݈Y[W���ߪA��IW��^D�t/��Sat=n�d��WZ�Ϗ<�m���G����#������&h�u�恤���6�s�z������|�T�_|�3�#�W��ܨS�);j��N�(e�IV���3�5ޘ$�D�	���x��[�1���̲a��H%��*3P}U�A�n�����\N�_��������$2#Ȳ�Q�m�����e�$V0�%���E[g�M:L�`,���ڀE��4r��ܗ����-��v~��^H+��[9F��ٹ��h{p�]%LD�Ư֛��5��E(jP�M4����r��~��{R�5x6��&Գ���4,l�2�cn��@$�o��!�ii"��B?n0��GMm7���#8]c��t�d���4\���S�$F�%S5w�8yr�#Ʃ�M�L8	P�{N�p>��zz�QC�����(^T�	 ҬD�a=�]T	9pQH&GOr4	���K� ث�C�?������;V�OD�S��4�=+�\:�{�Y�~X�h�������m.�����>�D���N�(�Uy�eYa�T�>E0����mF]<٘�ϯs��*�o,x�/_hY(AA�0y�-��1VJ�T�|[��!r�ÀY�6����^�m��i�"�	�(��B[8�q�V�g���&�wPfn��H'>(;�,�N���~rT�����#�v��>��p;�o|��5e���s"a�8�T�]����E|�ɼJ �C{�T��T����)��N�<R10*�n�@�#4A`=ʤ��u_�!+��뾜:���4������%gO��I�(��X���kN����Fa���}�S���e����;B<�Bԍ�ծd���_������#�3�e=�59�a�y�ۤ#��B�₺�с��E�����t>���;AЀp�sz�WQ�+�$�������ם�.c��j@�2�[W:u�V�v�>BK�V�
f��n$����A��T��d�Y�݅��6�sJA���s�?�/���qd�E�_,�����+����\�U��m��ޫ7ښQ/cm!$�QB�0�a�\�b�|)Б��b�n�P8"��c�" 2�ҧ~�y9�u:��1�V�xͥ6�m���7:�x��m&
��A��v������C� ����y��*���X��_����j���������	�4}t������<��ruMǞRmj��E@<wX�F=��"���OťZ�w|Z�� ���3iL��0q[1p�q���^���"����Y��mYD��&Jf�r+��E�d��Q�Kv����W�}����o�Y��l6$��M�-��(��������7<6��5��ԛ�e9��1��O�r!� a>D�W������O�ܵ�T�sQ�v��PM�T�.��Gɳm_���N��d��H�t	Ae3I2�v��~�Td,��d���R �����
�g��A7��aޠ��>5uI�o�\�G���ႊ=h�Ɨ���i�ġuO	�dU=�Ic`�T��3
���TM�S,�F�V8-ȋX���,���ɥz7���H湨�k�jS��)G~s-���`Y�쩂j��j����� �f�=Ԡm���$��ۂ���5#  0�Yr���jo���